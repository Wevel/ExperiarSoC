* NGSPICE file created from Video.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt Video sram_addr0[0] sram_addr0[1] sram_addr0[2] sram_addr0[3] sram_addr0[4]
+ sram_addr0[5] sram_addr0[6] sram_addr0[7] sram_addr0[8] sram_addr1[0] sram_addr1[1]
+ sram_addr1[2] sram_addr1[3] sram_addr1[4] sram_addr1[5] sram_addr1[6] sram_addr1[7]
+ sram_addr1[8] sram_clk0 sram_clk1 sram_csb0[0] sram_csb0[1] sram_csb0[2] sram_csb0[3]
+ sram_csb1[0] sram_csb1[1] sram_csb1[2] sram_csb1[3] sram_din0[0] sram_din0[10] sram_din0[11]
+ sram_din0[12] sram_din0[13] sram_din0[14] sram_din0[15] sram_din0[16] sram_din0[17]
+ sram_din0[18] sram_din0[19] sram_din0[1] sram_din0[20] sram_din0[21] sram_din0[22]
+ sram_din0[23] sram_din0[24] sram_din0[25] sram_din0[26] sram_din0[27] sram_din0[28]
+ sram_din0[29] sram_din0[2] sram_din0[30] sram_din0[31] sram_din0[3] sram_din0[4]
+ sram_din0[5] sram_din0[6] sram_din0[7] sram_din0[8] sram_din0[9] sram_dout0[0] sram_dout0[100]
+ sram_dout0[101] sram_dout0[102] sram_dout0[103] sram_dout0[104] sram_dout0[105]
+ sram_dout0[106] sram_dout0[107] sram_dout0[108] sram_dout0[109] sram_dout0[10] sram_dout0[110]
+ sram_dout0[111] sram_dout0[112] sram_dout0[113] sram_dout0[114] sram_dout0[115]
+ sram_dout0[116] sram_dout0[117] sram_dout0[118] sram_dout0[119] sram_dout0[11] sram_dout0[120]
+ sram_dout0[121] sram_dout0[122] sram_dout0[123] sram_dout0[124] sram_dout0[125]
+ sram_dout0[126] sram_dout0[127] sram_dout0[12] sram_dout0[13] sram_dout0[14] sram_dout0[15]
+ sram_dout0[16] sram_dout0[17] sram_dout0[18] sram_dout0[19] sram_dout0[1] sram_dout0[20]
+ sram_dout0[21] sram_dout0[22] sram_dout0[23] sram_dout0[24] sram_dout0[25] sram_dout0[26]
+ sram_dout0[27] sram_dout0[28] sram_dout0[29] sram_dout0[2] sram_dout0[30] sram_dout0[31]
+ sram_dout0[32] sram_dout0[33] sram_dout0[34] sram_dout0[35] sram_dout0[36] sram_dout0[37]
+ sram_dout0[38] sram_dout0[39] sram_dout0[3] sram_dout0[40] sram_dout0[41] sram_dout0[42]
+ sram_dout0[43] sram_dout0[44] sram_dout0[45] sram_dout0[46] sram_dout0[47] sram_dout0[48]
+ sram_dout0[49] sram_dout0[4] sram_dout0[50] sram_dout0[51] sram_dout0[52] sram_dout0[53]
+ sram_dout0[54] sram_dout0[55] sram_dout0[56] sram_dout0[57] sram_dout0[58] sram_dout0[59]
+ sram_dout0[5] sram_dout0[60] sram_dout0[61] sram_dout0[62] sram_dout0[63] sram_dout0[64]
+ sram_dout0[65] sram_dout0[66] sram_dout0[67] sram_dout0[68] sram_dout0[69] sram_dout0[6]
+ sram_dout0[70] sram_dout0[71] sram_dout0[72] sram_dout0[73] sram_dout0[74] sram_dout0[75]
+ sram_dout0[76] sram_dout0[77] sram_dout0[78] sram_dout0[79] sram_dout0[7] sram_dout0[80]
+ sram_dout0[81] sram_dout0[82] sram_dout0[83] sram_dout0[84] sram_dout0[85] sram_dout0[86]
+ sram_dout0[87] sram_dout0[88] sram_dout0[89] sram_dout0[8] sram_dout0[90] sram_dout0[91]
+ sram_dout0[92] sram_dout0[93] sram_dout0[94] sram_dout0[95] sram_dout0[96] sram_dout0[97]
+ sram_dout0[98] sram_dout0[99] sram_dout0[9] sram_dout1[0] sram_dout1[100] sram_dout1[101]
+ sram_dout1[102] sram_dout1[103] sram_dout1[104] sram_dout1[105] sram_dout1[106]
+ sram_dout1[107] sram_dout1[108] sram_dout1[109] sram_dout1[10] sram_dout1[110] sram_dout1[111]
+ sram_dout1[112] sram_dout1[113] sram_dout1[114] sram_dout1[115] sram_dout1[116]
+ sram_dout1[117] sram_dout1[118] sram_dout1[119] sram_dout1[11] sram_dout1[120] sram_dout1[121]
+ sram_dout1[122] sram_dout1[123] sram_dout1[124] sram_dout1[125] sram_dout1[126]
+ sram_dout1[127] sram_dout1[12] sram_dout1[13] sram_dout1[14] sram_dout1[15] sram_dout1[16]
+ sram_dout1[17] sram_dout1[18] sram_dout1[19] sram_dout1[1] sram_dout1[20] sram_dout1[21]
+ sram_dout1[22] sram_dout1[23] sram_dout1[24] sram_dout1[25] sram_dout1[26] sram_dout1[27]
+ sram_dout1[28] sram_dout1[29] sram_dout1[2] sram_dout1[30] sram_dout1[31] sram_dout1[32]
+ sram_dout1[33] sram_dout1[34] sram_dout1[35] sram_dout1[36] sram_dout1[37] sram_dout1[38]
+ sram_dout1[39] sram_dout1[3] sram_dout1[40] sram_dout1[41] sram_dout1[42] sram_dout1[43]
+ sram_dout1[44] sram_dout1[45] sram_dout1[46] sram_dout1[47] sram_dout1[48] sram_dout1[49]
+ sram_dout1[4] sram_dout1[50] sram_dout1[51] sram_dout1[52] sram_dout1[53] sram_dout1[54]
+ sram_dout1[55] sram_dout1[56] sram_dout1[57] sram_dout1[58] sram_dout1[59] sram_dout1[5]
+ sram_dout1[60] sram_dout1[61] sram_dout1[62] sram_dout1[63] sram_dout1[64] sram_dout1[65]
+ sram_dout1[66] sram_dout1[67] sram_dout1[68] sram_dout1[69] sram_dout1[6] sram_dout1[70]
+ sram_dout1[71] sram_dout1[72] sram_dout1[73] sram_dout1[74] sram_dout1[75] sram_dout1[76]
+ sram_dout1[77] sram_dout1[78] sram_dout1[79] sram_dout1[7] sram_dout1[80] sram_dout1[81]
+ sram_dout1[82] sram_dout1[83] sram_dout1[84] sram_dout1[85] sram_dout1[86] sram_dout1[87]
+ sram_dout1[88] sram_dout1[89] sram_dout1[8] sram_dout1[90] sram_dout1[91] sram_dout1[92]
+ sram_dout1[93] sram_dout1[94] sram_dout1[95] sram_dout1[96] sram_dout1[97] sram_dout1[98]
+ sram_dout1[99] sram_dout1[9] sram_web0 sram_wmask0[0] sram_wmask0[1] sram_wmask0[2]
+ sram_wmask0[3] vccd1 vga_b[0] vga_b[1] vga_g[0] vga_g[1] vga_hsync vga_r[0] vga_r[1]
+ vga_vsync vssd1 wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12] wb_adr_i[13]
+ wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19] wb_adr_i[1]
+ wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[2] wb_adr_i[3] wb_adr_i[4]
+ wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_data_i[0]
+ wb_data_i[10] wb_data_i[11] wb_data_i[12] wb_data_i[13] wb_data_i[14] wb_data_i[15]
+ wb_data_i[16] wb_data_i[17] wb_data_i[18] wb_data_i[19] wb_data_i[1] wb_data_i[20]
+ wb_data_i[21] wb_data_i[22] wb_data_i[23] wb_data_i[24] wb_data_i[25] wb_data_i[26]
+ wb_data_i[27] wb_data_i[28] wb_data_i[29] wb_data_i[2] wb_data_i[30] wb_data_i[31]
+ wb_data_i[3] wb_data_i[4] wb_data_i[5] wb_data_i[6] wb_data_i[7] wb_data_i[8] wb_data_i[9]
+ wb_data_o[0] wb_data_o[10] wb_data_o[11] wb_data_o[12] wb_data_o[13] wb_data_o[14]
+ wb_data_o[15] wb_data_o[16] wb_data_o[17] wb_data_o[18] wb_data_o[19] wb_data_o[1]
+ wb_data_o[20] wb_data_o[21] wb_data_o[22] wb_data_o[23] wb_data_o[24] wb_data_o[25]
+ wb_data_o[26] wb_data_o[27] wb_data_o[28] wb_data_o[29] wb_data_o[2] wb_data_o[30]
+ wb_data_o[31] wb_data_o[3] wb_data_o[4] wb_data_o[5] wb_data_o[6] wb_data_o[7] wb_data_o[8]
+ wb_data_o[9] wb_error_o wb_rst_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2] wb_sel_i[3]
+ wb_stall_o wb_stb_i wb_we_i
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2106_ _2046_/A _2105_/B _2105_/Y _2094_/X vssd1 vssd1 vccd1 vccd1 _2406_/D sky130_fd_sc_hd__a211o_1
X_2037_ _2071_/A vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__buf_2
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1270_ _1270_/A1 _1190_/A _1194_/A _1270_/B2 vssd1 vssd1 vccd1 vccd1 _1270_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput401 _1504_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_172_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1606_ _1609_/C _1606_/B vssd1 vssd1 vccd1 vccd1 _2306_/D sky130_fd_sc_hd__nor2_1
Xoutput412 _1424_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1537_ _2283_/Q _1537_/B vssd1 vssd1 vccd1 vccd1 _1538_/A sky130_fd_sc_hd__and2_2
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1468_ input15/X _1443_/X _1447_/X _1467_/X vssd1 vssd1 vccd1 vccd1 _1468_/X sky130_fd_sc_hd__a211o_2
XFILLER_170_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1399_ input1/X _1385_/X _1395_/X _1398_/X vssd1 vssd1 vccd1 vccd1 _1399_/X sky130_fd_sc_hd__o211a_4
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2440_ _2446_/CLK _2440_/D vssd1 vssd1 vccd1 vccd1 _2440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ _2474_/A _2371_/D vssd1 vssd1 vccd1 vccd1 _2371_/Q sky130_fd_sc_hd__dfxtp_1
X_1322_ _1322_/A1 _1187_/A _1224_/X _1322_/B2 vssd1 vssd1 vccd1 vccd1 _1322_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1253_ _1208_/X _1250_/X _1252_/X _1200_/X vssd1 vssd1 vccd1 vccd1 _1259_/A sky130_fd_sc_hd__a22o_1
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1184_ _2294_/Q vssd1 vssd1 vccd1 vccd1 _1327_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_4 _1278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ _2079_/A vssd1 vssd1 vccd1 vccd1 _1940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _2360_/Q _2243_/A _1794_/X _2358_/Q vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2423_ _2435_/CLK _2423_/D vssd1 vssd1 vccd1 vccd1 _2423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2354_ _2459_/CLK _2354_/D vssd1 vssd1 vccd1 vccd1 _2354_/Q sky130_fd_sc_hd__dfxtp_1
X_1305_ _1234_/X _1302_/X _1304_/X _1200_/X vssd1 vssd1 vccd1 vccd1 _1311_/A sky130_fd_sc_hd__a22o_1
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2285_ _2475_/A _2285_/D vssd1 vssd1 vccd1 vccd1 _2285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1236_ _1236_/A1 _1215_/A _1235_/X _1236_/B2 vssd1 vssd1 vccd1 vccd1 _1236_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1167_ _2313_/Q vssd1 vssd1 vccd1 vccd1 _1629_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1098_ _1098_/A vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__buf_4
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ _1102_/X _2054_/A _2069_/X vssd1 vssd1 vccd1 vccd1 _2394_/D sky130_fd_sc_hd__a21o_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1923_ _2346_/Q _1912_/Y _1922_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _2346_/D sky130_fd_sc_hd__a211o_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1854_ _2385_/Q vssd1 vssd1 vccd1 vccd1 _2044_/A sky130_fd_sc_hd__inv_2
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1785_ _1783_/Y _2469_/Q _1808_/A _2363_/Q vssd1 vssd1 vccd1 vccd1 _1789_/C sky130_fd_sc_hd__o22a_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2406_ _2472_/CLK _2406_/D vssd1 vssd1 vccd1 vccd1 _2406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _2337_/CLK _2337_/D vssd1 vssd1 vccd1 vccd1 _2337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2268_ _2272_/B vssd1 vssd1 vccd1 vccd1 _2269_/C sky130_fd_sc_hd__clkinv_2
X_1219_ _2293_/Q vssd1 vssd1 vccd1 vccd1 _1308_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2199_ _2199_/A vssd1 vssd1 vccd1 vccd1 _2443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput301 wb_data_i[7] vssd1 vssd1 vccd1 vccd1 _1118_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1570_ _1577_/D _1570_/B vssd1 vssd1 vccd1 vccd1 _2297_/D sky130_fd_sc_hd__nor2_1
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2122_ _1111_/A _2112_/X _2121_/Y _2116_/X vssd1 vssd1 vccd1 vccd1 _2411_/D sky130_fd_sc_hd__a211o_1
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2053_ _2053_/A vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1906_ _1906_/A vssd1 vssd1 vccd1 vccd1 _2343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1837_ _1681_/X _1836_/C _2336_/Q vssd1 vssd1 vccd1 vccd1 _1838_/C sky130_fd_sc_hd__a21oi_1
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1768_ _2368_/Q vssd1 vssd1 vccd1 vccd1 _1768_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1699_ _2334_/Q vssd1 vssd1 vccd1 vccd1 _1699_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput120 sram_dout0[92] vssd1 vssd1 vccd1 vccd1 _1516_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput142 sram_dout1[111] vssd1 vssd1 vccd1 vccd1 _1293_/C sky130_fd_sc_hd__clkbuf_1
Xinput131 sram_dout1[101] vssd1 vssd1 vccd1 vccd1 _1318_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput153 sram_dout1[121] vssd1 vssd1 vccd1 vccd1 _1256_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput175 sram_dout1[28] vssd1 vssd1 vccd1 vccd1 _1312_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput186 sram_dout1[3] vssd1 vssd1 vccd1 vccd1 _1282_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 sram_dout1[18] vssd1 vssd1 vccd1 vccd1 _1237_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput197 sram_dout1[4] vssd1 vssd1 vccd1 vccd1 _1315_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1622_ _1646_/B vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1553_ _2283_/Q _1553_/A1 _2187_/S vssd1 vssd1 vccd1 vccd1 _1554_/A sky130_fd_sc_hd__mux2_1
X_1484_ _1505_/A vssd1 vssd1 vccd1 vccd1 _1484_/X sky130_fd_sc_hd__buf_2
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2105_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2036_ _1102_/X _2019_/X _2035_/X vssd1 vssd1 vccd1 vccd1 _2383_/D sky130_fd_sc_hd__a21o_1
XFILLER_23_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput402 _1508_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_160_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1605_ _1602_/A _1656_/B _1646_/B vssd1 vssd1 vccd1 vccd1 _1606_/B sky130_fd_sc_hd__o21ai_1
XFILLER_133_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput413 _1428_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_160_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1536_ _1536_/A vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1467_ input71/X _1448_/X _1449_/X _1467_/B2 vssd1 vssd1 vccd1 vccd1 _1467_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1398_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1398_/X sky130_fd_sc_hd__buf_2
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2019_ _2022_/A vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2370_ _2474_/A _2370_/D vssd1 vssd1 vccd1 vccd1 _2370_/Q sky130_fd_sc_hd__dfxtp_1
X_1321_ _1321_/A _1321_/B vssd1 vssd1 vccd1 vccd1 _1321_/X sky130_fd_sc_hd__and2_1
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1252_ _1252_/A1 _1191_/A _1195_/A _1252_/B2 _1251_/X vssd1 vssd1 vccd1 vccd1 _1252_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2413_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1183_ _1183_/A vssd1 vssd1 vccd1 vccd1 _2294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_5 _1315_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1519_ input86/X _1490_/A _1489_/A _1519_/B2 vssd1 vssd1 vccd1 vccd1 _1519_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1870_ _2353_/Q vssd1 vssd1 vccd1 vccd1 _1943_/A sky130_fd_sc_hd__inv_2
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2422_ _2459_/CLK _2422_/D vssd1 vssd1 vccd1 vccd1 _2422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2353_ _2459_/CLK _2353_/D vssd1 vssd1 vccd1 vccd1 _2353_/Q sky130_fd_sc_hd__dfxtp_1
X_1304_ _1304_/A1 _1191_/A _1195_/A _1304_/B2 _1303_/X vssd1 vssd1 vccd1 vccd1 _1304_/X
+ sky130_fd_sc_hd__a221o_1
X_2284_ _2475_/A _2284_/D vssd1 vssd1 vccd1 vccd1 _2284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1235_ _1235_/A vssd1 vssd1 vccd1 vccd1 _1235_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1166_ _1166_/A vssd1 vssd1 vccd1 vccd1 _2287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1097_ _2102_/A vssd1 vssd1 vccd1 vccd1 _1098_/A sky130_fd_sc_hd__inv_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1999_ _2370_/Q _1984_/X _1998_/Y vssd1 vssd1 vccd1 vccd1 _2370_/D sky130_fd_sc_hd__o21a_1
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _1922_/A _1922_/B vssd1 vssd1 vccd1 vccd1 _1922_/X sky130_fd_sc_hd__and2_1
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1853_ _2393_/Q _1805_/A _2267_/A _1851_/Y _1852_/X vssd1 vssd1 vccd1 vccd1 _1853_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1784_ _2366_/Q _2264_/A _2272_/A _1783_/Y vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2405_ _2414_/CLK _2405_/D vssd1 vssd1 vccd1 vccd1 _2405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2336_ _2337_/CLK _2336_/D vssd1 vssd1 vccd1 vccd1 _2336_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2267_ _2267_/A _2267_/B _2267_/C _2267_/D vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__and4_1
X_1218_ _2294_/Q vssd1 vssd1 vccd1 vccd1 _1308_/A sky130_fd_sc_hd__clkbuf_1
X_2198_ _2443_/Q _2198_/A1 _2198_/S vssd1 vssd1 vccd1 vccd1 _2199_/A sky130_fd_sc_hd__mux2_1
X_1149_ _1149_/A vssd1 vssd1 vccd1 vccd1 _1149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput302 wb_data_i[8] vssd1 vssd1 vccd1 vccd1 _1120_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2121_ _2121_/A _2121_/B vssd1 vssd1 vccd1 vccd1 _2121_/Y sky130_fd_sc_hd__nor2_1
X_2052_ _2136_/A _2052_/B _2167_/B vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__nor3_2
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1905_ _2116_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _1906_/A sky130_fd_sc_hd__and2b_1
X_1836_ _1836_/A _2336_/Q _1836_/C vssd1 vssd1 vccd1 vccd1 _1839_/B sky130_fd_sc_hd__and3_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1767_ _2371_/Q _2462_/Q vssd1 vssd1 vccd1 vccd1 _1790_/A sky130_fd_sc_hd__xor2_1
XFILLER_143_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1698_ _1831_/A vssd1 vssd1 vccd1 vccd1 _1698_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2319_/CLK _2319_/D vssd1 vssd1 vccd1 vccd1 _2319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 sram_dout0[83] vssd1 vssd1 vccd1 vccd1 _1481_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput132 sram_dout1[102] vssd1 vssd1 vccd1 vccd1 _1205_/C sky130_fd_sc_hd__clkbuf_1
Xinput143 sram_dout1[112] vssd1 vssd1 vccd1 vccd1 _1306_/C sky130_fd_sc_hd__clkbuf_1
Xinput154 sram_dout1[122] vssd1 vssd1 vccd1 vccd1 _1272_/C sky130_fd_sc_hd__clkbuf_1
Xinput121 sram_dout0[93] vssd1 vssd1 vccd1 vccd1 _1519_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput176 sram_dout1[29] vssd1 vssd1 vccd1 vccd1 _1319_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput165 sram_dout1[19] vssd1 vssd1 vccd1 vccd1 _1261_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput187 sram_dout1[40] vssd1 vssd1 vccd1 vccd1 _1266_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput198 sram_dout1[50] vssd1 vssd1 vccd1 vccd1 _1210_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1621_ _1621_/A _1621_/B _1621_/C vssd1 vssd1 vccd1 vccd1 _1621_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1552_ _1552_/A vssd1 vssd1 vccd1 vccd1 _2282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1483_ input39/X _1463_/X _1477_/X _1482_/X vssd1 vssd1 vccd1 vccd1 _1483_/X sky130_fd_sc_hd__o211a_4
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2104_ _2157_/A _2109_/B _2157_/C vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__nor3_4
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2035_ _2383_/Q _2023_/X _2002_/X vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1819_ _2376_/Q _2468_/Q vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__xor2_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1604_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1646_/B sky130_fd_sc_hd__clkbuf_2
Xoutput414 _1431_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[7] sky130_fd_sc_hd__buf_2
Xoutput403 _1511_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_141_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1535_ _2282_/Q _1537_/B vssd1 vssd1 vccd1 vccd1 _1536_/A sky130_fd_sc_hd__and2_2
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1466_ input35/X _1463_/X _1459_/X _1465_/X vssd1 vssd1 vccd1 vccd1 _1466_/X sky130_fd_sc_hd__o211a_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1397_ _1518_/A vssd1 vssd1 vccd1 vccd1 _1438_/A sky130_fd_sc_hd__buf_2
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _2136_/A _2052_/B _2018_/C vssd1 vssd1 vccd1 vccd1 _2022_/A sky130_fd_sc_hd__nor3_2
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1320_ _1320_/A1 _1200_/X _1208_/X _1320_/B2 _1319_/X vssd1 vssd1 vccd1 vccd1 _1320_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1251_ _1251_/A _1251_/B _1251_/C vssd1 vssd1 vccd1 vccd1 _1251_/X sky130_fd_sc_hd__and3_1
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1182_ _2301_/Q _2319_/Q _1182_/S vssd1 vssd1 vccd1 vccd1 _1183_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_6 _1340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1518_ _1518_/A vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__buf_4
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1449_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1449_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2421_ _2425_/CLK _2421_/D vssd1 vssd1 vccd1 vccd1 _2421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2352_ _2459_/CLK _2352_/D vssd1 vssd1 vccd1 vccd1 _2352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1303_ _1303_/A _1303_/B _1303_/C vssd1 vssd1 vccd1 vccd1 _1303_/X sky130_fd_sc_hd__and3_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2283_ _2446_/CLK _2283_/D vssd1 vssd1 vccd1 vccd1 _2283_/Q sky130_fd_sc_hd__dfxtp_1
X_1234_ _1234_/A vssd1 vssd1 vccd1 vccd1 _1234_/X sky130_fd_sc_hd__buf_2
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1165_ _2305_/Q _2312_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1166_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1096_ _1096_/A _1118_/B vssd1 vssd1 vccd1 vccd1 _2102_/A sky130_fd_sc_hd__nand2_4
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1998_ _1107_/A _1986_/A _1995_/X vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1921_ _2345_/Q _1918_/X _1920_/Y vssd1 vssd1 vccd1 vccd1 _2345_/D sky130_fd_sc_hd__o21a_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1852_ _2388_/Q _1781_/A _1808_/A _2385_/Q vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1783_ _2364_/Q vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2404_ _2414_/CLK _2404_/D vssd1 vssd1 vccd1 vccd1 _2404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2335_ _2434_/CLK _2335_/D vssd1 vssd1 vccd1 vccd1 _2335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2266_ _2261_/A _2267_/B _2267_/D _2267_/C vssd1 vssd1 vccd1 vccd1 _2269_/B sky130_fd_sc_hd__a31o_1
X_1217_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1217_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2197_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1148_ _2444_/Q _1150_/B vssd1 vssd1 vccd1 vccd1 _1149_/A sky130_fd_sc_hd__and2_2
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput303 wb_data_i[9] vssd1 vssd1 vccd1 vccd1 _1122_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2120_ _2410_/Q _2111_/X _2119_/Y vssd1 vssd1 vccd1 vccd1 _2410_/D sky130_fd_sc_hd__o21a_1
XFILLER_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2051_ _2387_/Q _2043_/X _2050_/Y vssd1 vssd1 vccd1 vccd1 _2387_/D sky130_fd_sc_hd__o21a_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1904_ _1121_/Y _2343_/Q _1904_/S vssd1 vssd1 vccd1 vccd1 _1905_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1835_ _1681_/X _1836_/C _1834_/Y vssd1 vssd1 vccd1 vccd1 _2335_/D sky130_fd_sc_hd__a21oi_1
X_1766_ _2372_/Q _2238_/B vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__xor2_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1697_ _2416_/Q vssd1 vssd1 vccd1 vccd1 _2132_/A sky130_fd_sc_hd__inv_2
XFILLER_171_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2319_/CLK _2318_/D vssd1 vssd1 vccd1 vccd1 _2318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2249_ _2262_/A _2249_/B _2249_/C vssd1 vssd1 vccd1 vccd1 _2250_/A sky130_fd_sc_hd__and3_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput111 sram_dout0[84] vssd1 vssd1 vccd1 vccd1 _1487_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput100 sram_dout0[74] vssd1 vssd1 vccd1 vccd1 _1444_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput144 sram_dout1[113] vssd1 vssd1 vccd1 vccd1 _1324_/C sky130_fd_sc_hd__clkbuf_2
Xinput133 sram_dout1[103] vssd1 vssd1 vccd1 vccd1 _1251_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput122 sram_dout0[94] vssd1 vssd1 vccd1 vccd1 _1522_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput177 sram_dout1[2] vssd1 vssd1 vccd1 vccd1 _1279_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput166 sram_dout1[1] vssd1 vssd1 vccd1 vccd1 _1263_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput155 sram_dout1[123] vssd1 vssd1 vccd1 vccd1 _1295_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput199 sram_dout1[51] vssd1 vssd1 vccd1 vccd1 _1250_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput188 sram_dout1[41] vssd1 vssd1 vccd1 vccd1 _1291_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1620_ _1621_/A _1621_/B _1621_/C vssd1 vssd1 vccd1 vccd1 _1620_/X sky130_fd_sc_hd__a21o_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1551_ _2282_/Q _1551_/A1 _2187_/S vssd1 vssd1 vccd1 vccd1 _1552_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1482_ input18/X _1473_/X _1478_/X _1481_/X vssd1 vssd1 vccd1 vccd1 _1482_/X sky130_fd_sc_hd__a211o_2
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2103_ _2405_/Q _2100_/B _2102_/Y _2094_/X vssd1 vssd1 vccd1 vccd1 _2405_/D sky130_fd_sc_hd__a211o_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2034_ _1105_/X _2022_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _2382_/D sky130_fd_sc_hd__a21o_1
XFILLER_35_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1818_ _1806_/X _1818_/B _1818_/C _1818_/D vssd1 vssd1 vccd1 vccd1 _1818_/X sky130_fd_sc_hd__and4b_1
XFILLER_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1749_ _2428_/Q _1749_/B vssd1 vssd1 vccd1 vccd1 _1749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1603_ _1587_/B _1602_/B _1656_/A vssd1 vssd1 vccd1 vccd1 _1648_/A sky130_fd_sc_hd__a21oi_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput415 _1437_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[8] sky130_fd_sc_hd__buf_2
Xoutput404 _1514_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1534_ _2157_/A vssd1 vssd1 vccd1 vccd1 _1534_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1465_ _1465_/A1 _1432_/X _1464_/X _1435_/X vssd1 vssd1 vccd1 vccd1 _1465_/X sky130_fd_sc_hd__a211o_2
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1396_ _2471_/Q _2472_/Q vssd1 vssd1 vccd1 vccd1 _1518_/A sky130_fd_sc_hd__nor2b_4
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2017_ _1121_/Y _2013_/B _2015_/X _2016_/X vssd1 vssd1 vccd1 vccd1 _2376_/D sky130_fd_sc_hd__a211o_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1250_ _1250_/A1 _1201_/X _1202_/X _1250_/B2 _1249_/X vssd1 vssd1 vccd1 vccd1 _1250_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1181_ _1181_/A vssd1 vssd1 vccd1 vccd1 _2293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1517_ input49/X _1505_/X _1501_/X _1516_/X vssd1 vssd1 vccd1 vccd1 _1517_/X sky130_fd_sc_hd__o211a_4
XINSDIODE2_7 _1342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1448_ _1479_/A vssd1 vssd1 vccd1 vccd1 _1448_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1379_ _1379_/A _1379_/B vssd1 vssd1 vccd1 vccd1 _1380_/A sky130_fd_sc_hd__and2_1
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2420_ _2425_/CLK _2420_/D vssd1 vssd1 vccd1 vccd1 _2420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2351_ _2413_/CLK _2351_/D vssd1 vssd1 vccd1 vccd1 _2351_/Q sky130_fd_sc_hd__dfxtp_1
X_1302_ _1302_/A1 _1201_/X _1202_/X _1302_/B2 _1301_/X vssd1 vssd1 vccd1 vccd1 _1302_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2282_ _2446_/CLK _2282_/D vssd1 vssd1 vccd1 vccd1 _2282_/Q sky130_fd_sc_hd__dfxtp_1
X_1233_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1233_/X sky130_fd_sc_hd__buf_2
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1164_ _1164_/A vssd1 vssd1 vccd1 vccd1 _2286_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1095_ _1099_/A vssd1 vssd1 vccd1 vccd1 _1118_/B sky130_fd_sc_hd__buf_6
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1997_ _2369_/Q _1984_/X _1996_/Y vssd1 vssd1 vccd1 vccd1 _2369_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XVideo_418 vssd1 vssd1 vccd1 vccd1 Video_418/HI wb_error_o sky130_fd_sc_hd__conb_1
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ _2089_/A _1918_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1851_ _2389_/Q vssd1 vssd1 vccd1 vccd1 _1851_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1782_ _2469_/Q vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2403_ _2413_/CLK _2403_/D vssd1 vssd1 vccd1 vccd1 _2403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2334_ _2337_/CLK _2334_/D vssd1 vssd1 vccd1 vccd1 _2334_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2265_ _2264_/A _2264_/B _2264_/Y _2239_/A vssd1 vssd1 vccd1 vccd1 _2467_/D sky130_fd_sc_hd__o211a_1
X_1216_ _1287_/A vssd1 vssd1 vccd1 vccd1 _1216_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2196_ _2442_/Q _2196_/A1 _2198_/S vssd1 vssd1 vccd1 vccd1 _2197_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1147_ _1147_/A vssd1 vssd1 vccd1 vccd1 _1147_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput304 wb_rst_i vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__buf_2
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2050_ _2049_/X _2043_/X _2030_/X vssd1 vssd1 vccd1 vccd1 _2050_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ _1952_/A vssd1 vssd1 vccd1 vccd1 _2116_/A sky130_fd_sc_hd__buf_2
X_1834_ _1681_/X _1836_/C _1825_/X vssd1 vssd1 vccd1 vccd1 _1834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1765_ _2461_/Q vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1696_ _1749_/B vssd1 vssd1 vccd1 vccd1 _1696_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2319_/CLK _2317_/D vssd1 vssd1 vccd1 vccd1 _2317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2248_ _2248_/A _2248_/B vssd1 vssd1 vccd1 vccd1 _2249_/C sky130_fd_sc_hd__nand2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2179_ _2434_/Q _2171_/B _1889_/X vssd1 vssd1 vccd1 vccd1 _2179_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput101 sram_dout0[75] vssd1 vssd1 vccd1 vccd1 _1450_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput134 sram_dout1[104] vssd1 vssd1 vccd1 vccd1 _1265_/C sky130_fd_sc_hd__clkbuf_1
Xinput145 sram_dout1[114] vssd1 vssd1 vccd1 vccd1 _1209_/C sky130_fd_sc_hd__clkbuf_1
Xinput123 sram_dout0[95] vssd1 vssd1 vccd1 vccd1 _1526_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput112 sram_dout0[85] vssd1 vssd1 vccd1 vccd1 _1493_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput167 sram_dout1[20] vssd1 vssd1 vccd1 vccd1 _1277_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput156 sram_dout1[124] vssd1 vssd1 vccd1 vccd1 _1308_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput178 sram_dout1[32] vssd1 vssd1 vccd1 vccd1 _1246_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput189 sram_dout1[42] vssd1 vssd1 vccd1 vccd1 _1304_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1550_ _1550_/A vssd1 vssd1 vccd1 vccd1 _2281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2319_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_141_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1481_ input75/X _1479_/X _1480_/X _1481_/B2 vssd1 vssd1 vccd1 vccd1 _1481_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2102_ _2102_/A _2102_/B vssd1 vssd1 vccd1 vccd1 _2102_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2033_ _2382_/Q _2023_/X _2002_/X vssd1 vssd1 vccd1 vccd1 _2033_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1817_ _2384_/Q _2235_/A _2267_/B _2020_/A _1816_/X vssd1 vssd1 vccd1 vccd1 _1818_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1748_ _2429_/Q _2337_/Q vssd1 vssd1 vccd1 vccd1 _1748_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1679_ _2414_/Q vssd1 vssd1 vccd1 vccd1 _1679_/Y sky130_fd_sc_hd__inv_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1602_ _1602_/A _1602_/B vssd1 vssd1 vccd1 vccd1 _1609_/C sky130_fd_sc_hd__and2_1
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput416 _1441_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput405 _1517_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1533_ _2042_/A vssd1 vssd1 vccd1 vccd1 _2157_/A sky130_fd_sc_hd__clkbuf_4
X_1464_ input14/X _1425_/X _1433_/X input70/X vssd1 vssd1 vccd1 vccd1 _1464_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1395_ _1395_/A1 _1443_/A _1492_/A _1394_/X vssd1 vssd1 vccd1 vccd1 _1395_/X sky130_fd_sc_hd__a211o_4
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2016_ _2116_/A vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__buf_4
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1180_ _2300_/Q _2318_/Q _1180_/S vssd1 vssd1 vccd1 vccd1 _1181_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1516_ _1516_/A1 _1489_/X _1515_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__a211o_2
XFILLER_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1447_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_8 _1129_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1378_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1378_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ _2414_/CLK _2350_/D vssd1 vssd1 vccd1 vccd1 _2350_/Q sky130_fd_sc_hd__dfxtp_1
X_1301_ _1301_/A _1301_/B _1301_/C vssd1 vssd1 vccd1 vccd1 _1301_/X sky130_fd_sc_hd__and3_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2281_ _2446_/CLK _2281_/D vssd1 vssd1 vccd1 vccd1 _2281_/Q sky130_fd_sc_hd__dfxtp_1
X_1232_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1314_/A sky130_fd_sc_hd__inv_2
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1163_ _2304_/Q _1621_/C _1168_/S vssd1 vssd1 vccd1 vccd1 _1164_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1094_ _2472_/Q _2471_/Q vssd1 vssd1 vccd1 vccd1 _1099_/A sky130_fd_sc_hd__and2b_1
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1996_ _2093_/A _1986_/A _1995_/X vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2315_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ _2387_/Q _2267_/C vssd1 vssd1 vccd1 vccd1 _1850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1781_ _1781_/A vssd1 vssd1 vccd1 vccd1 _2264_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2402_ _2452_/CLK _2402_/D vssd1 vssd1 vccd1 vccd1 _2402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2333_ _2337_/CLK _2333_/D vssd1 vssd1 vccd1 vccd1 _2333_/Q sky130_fd_sc_hd__dfxtp_1
X_2264_ _2264_/A _2264_/B vssd1 vssd1 vccd1 vccd1 _2264_/Y sky130_fd_sc_hd__nand2_1
X_1215_ _1215_/A vssd1 vssd1 vccd1 vccd1 _1240_/A sky130_fd_sc_hd__buf_2
X_2195_ _2195_/A vssd1 vssd1 vccd1 vccd1 _2441_/D sky130_fd_sc_hd__clkbuf_1
X_1146_ _2443_/Q _1150_/B vssd1 vssd1 vccd1 vccd1 _1147_/A sky130_fd_sc_hd__and2_2
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1979_ _1976_/X _2364_/Q vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__and2b_1
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput305 wb_sel_i[0] vssd1 vssd1 vccd1 vccd1 _1547_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1902_ _1902_/A vssd1 vssd1 vccd1 vccd1 _2342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1833_ _1836_/C _1833_/B vssd1 vssd1 vccd1 vccd1 _2334_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1764_ _1732_/X _1734_/X _1745_/X _1846_/A _1562_/X vssd1 vssd1 vccd1 vccd1 _2329_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1695_ _2424_/Q _1828_/B vssd1 vssd1 vccd1 vccd1 _1695_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_171_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2316_/CLK _2316_/D vssd1 vssd1 vccd1 vccd1 _2316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2255_/C vssd1 vssd1 vccd1 vccd1 _2249_/B sky130_fd_sc_hd__clkinv_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2178_ _2433_/Q _2163_/X _2177_/Y vssd1 vssd1 vccd1 vccd1 _2433_/D sky130_fd_sc_hd__o21a_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1129_ _2040_/A _1909_/A vssd1 vssd1 vccd1 vccd1 _1129_/Y sky130_fd_sc_hd__nor2_2
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 sram_dout0[76] vssd1 vssd1 vccd1 vccd1 _1454_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput135 sram_dout1[105] vssd1 vssd1 vccd1 vccd1 _1290_/C sky130_fd_sc_hd__clkbuf_1
Xinput124 sram_dout0[96] vssd1 vssd1 vccd1 vccd1 _1395_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput113 sram_dout0[86] vssd1 vssd1 vccd1 vccd1 _1496_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput168 sram_dout1[21] vssd1 vssd1 vccd1 vccd1 _1286_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput157 sram_dout1[125] vssd1 vssd1 vccd1 vccd1 _1322_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput146 sram_dout1[115] vssd1 vssd1 vccd1 vccd1 _1249_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput179 sram_dout1[33] vssd1 vssd1 vccd1 vccd1 _1263_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1480_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1480_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2101_ _2404_/Q _2084_/X _2100_/Y _2094_/X vssd1 vssd1 vccd1 vccd1 _2404_/D sky130_fd_sc_hd__a211o_1
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2032_ _2381_/Q _2022_/X _2031_/Y vssd1 vssd1 vccd1 vccd1 _2381_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1816_ _2378_/Q _1777_/Y _1815_/Y _2383_/Q vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1747_ _2429_/Q _2337_/Q vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__or2_1
XFILLER_171_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1678_ _2408_/Q _1749_/B vssd1 vssd1 vccd1 vccd1 _1691_/B sky130_fd_sc_hd__xor2_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1601_ _2305_/Q _1598_/A _1600_/X vssd1 vssd1 vccd1 vccd1 _2305_/D sky130_fd_sc_hd__o21ba_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput417 _2437_/Q vssd1 vssd1 vccd1 vccd1 wb_stall_o sky130_fd_sc_hd__buf_2
Xoutput406 _1521_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[29] sky130_fd_sc_hd__buf_2
X_1532_ _1899_/A vssd1 vssd1 vccd1 vccd1 _2042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1463_ _1505_/A vssd1 vssd1 vccd1 vccd1 _1463_/X sky130_fd_sc_hd__buf_2
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1394_ input54/X _1490_/A _1489_/A input89/X vssd1 vssd1 vccd1 vccd1 _1394_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2015_ _2010_/A _2376_/Q vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__and2b_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1515_ input28/X _1485_/X _1490_/X input85/X vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1446_ input12/X _1442_/X _1438_/X _1445_/X vssd1 vssd1 vccd1 vccd1 _1446_/X sky130_fd_sc_hd__o211a_4
XINSDIODE2_9 _1108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1377_ _1377_/A _1379_/B vssd1 vssd1 vccd1 vccd1 _1378_/A sky130_fd_sc_hd__and2_1
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1300_ _1241_/X _1282_/X _1283_/X _1299_/X vssd1 vssd1 vccd1 vccd1 _1300_/X sky130_fd_sc_hd__a31o_4
XFILLER_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2280_ _2446_/CLK _2280_/D vssd1 vssd1 vccd1 vccd1 _2280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1231_ _1231_/A _1231_/B vssd1 vssd1 vccd1 vccd1 _1231_/X sky130_fd_sc_hd__or2_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1162_ _2311_/Q vssd1 vssd1 vccd1 vccd1 _1621_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1995_ _2079_/A vssd1 vssd1 vccd1 vccd1 _1995_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1429_ input61/X _1409_/X _1410_/X input97/X vssd1 vssd1 vccd1 vccd1 _1429_/X sky130_fd_sc_hd__a22o_1
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1780_ _2467_/Q vssd1 vssd1 vccd1 vccd1 _1781_/A sky130_fd_sc_hd__inv_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2401_ _2413_/CLK _2401_/D vssd1 vssd1 vccd1 vccd1 _2401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2332_ _2414_/CLK _2332_/D vssd1 vssd1 vccd1 vccd1 _2332_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2263_ _2263_/A vssd1 vssd1 vccd1 vccd1 _2466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1214_ _1587_/B vssd1 vssd1 vccd1 vccd1 _1215_/A sky130_fd_sc_hd__clkbuf_2
X_2194_ _2441_/Q _2194_/A1 _2198_/S vssd1 vssd1 vccd1 vccd1 _2195_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1145_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1978_ _2363_/Q _1976_/X _1977_/Y vssd1 vssd1 vccd1 vccd1 _2363_/D sky130_fd_sc_hd__o21a_1
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput306 wb_sel_i[1] vssd1 vssd1 vccd1 vccd1 _1549_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _1889_/X _1901_/B vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__and2b_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ _2334_/Q _1830_/B _1825_/X vssd1 vssd1 vccd1 vccd1 _1833_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1763_ _1763_/A vssd1 vssd1 vccd1 vccd1 _1846_/A sky130_fd_sc_hd__clkbuf_2
X_1694_ _2332_/Q vssd1 vssd1 vccd1 vccd1 _1828_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_171_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2315_/CLK _2315_/D vssd1 vssd1 vccd1 vccd1 _2315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2460_/Q _2461_/Q _2462_/Q _2463_/Q vssd1 vssd1 vccd1 vccd1 _2255_/C sky130_fd_sc_hd__and4_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2177_ _2098_/A _2164_/X _2185_/A vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1128_ _2472_/Q _2471_/Q vssd1 vssd1 vccd1 vccd1 _1909_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput136 sram_dout1[106] vssd1 vssd1 vccd1 vccd1 _1303_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput125 sram_dout0[97] vssd1 vssd1 vccd1 vccd1 _1403_/A1 sky130_fd_sc_hd__buf_2
Xinput114 sram_dout0[87] vssd1 vssd1 vccd1 vccd1 _1498_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput103 sram_dout0[77] vssd1 vssd1 vccd1 vccd1 _1456_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput169 sram_dout1[22] vssd1 vssd1 vccd1 vccd1 _1313_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput158 sram_dout1[12] vssd1 vssd1 vccd1 vccd1 _1236_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput147 sram_dout1[116] vssd1 vssd1 vccd1 vccd1 _1267_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2100_ _2100_/A _2100_/B vssd1 vssd1 vccd1 vccd1 _2100_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2031_ _1107_/A _2022_/A _2030_/X vssd1 vssd1 vccd1 vccd1 _2031_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1815_ _2461_/Q vssd1 vssd1 vccd1 vccd1 _1815_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1746_ _2432_/Q _2334_/Q vssd1 vssd1 vccd1 vccd1 _1761_/A sky130_fd_sc_hd__xor2_1
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1677_ _2338_/Q vssd1 vssd1 vccd1 vccd1 _1749_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2229_ _2457_/Q _2229_/A1 _2231_/S vssd1 vssd1 vccd1 vccd1 _2230_/A sky130_fd_sc_hd__mux2_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1600_ _2305_/Q _1598_/A _1656_/A vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput407 _1413_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_153_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1531_ _2281_/Q _1531_/B vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1462_ input34/X _1442_/X _1459_/X _1461_/X vssd1 vssd1 vccd1 vccd1 _1462_/X sky130_fd_sc_hd__o211a_4
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1393_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2014_ _1124_/X _2013_/B _2013_/Y _1944_/X vssd1 vssd1 vccd1 vccd1 _2375_/D sky130_fd_sc_hd__a211o_1
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1729_ _1749_/B vssd1 vssd1 vccd1 vccd1 _1845_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1514_ input48/X _1505_/X _1501_/X _1513_/X vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__o211a_4
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1445_ input8/X _1443_/X _1408_/X _1444_/X vssd1 vssd1 vccd1 vccd1 _1445_/X sky130_fd_sc_hd__a211o_2
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ _1376_/A vssd1 vssd1 vccd1 vccd1 _1376_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_1230_ _1240_/A _1221_/X _1223_/X _1226_/X _1229_/X vssd1 vssd1 vccd1 vccd1 _1231_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1161_ _1161_/A vssd1 vssd1 vccd1 vccd1 _2285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1994_ _2368_/Q _1984_/X _1993_/Y vssd1 vssd1 vccd1 vccd1 _2368_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1428_ input95/X _1421_/X _1417_/X _1427_/X vssd1 vssd1 vccd1 vccd1 _1428_/X sky130_fd_sc_hd__o211a_4
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1359_ _1359_/A vssd1 vssd1 vccd1 vccd1 _1359_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2400_ _2452_/CLK _2400_/D vssd1 vssd1 vccd1 vccd1 _2400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2331_ _2414_/CLK _2331_/D vssd1 vssd1 vccd1 vccd1 _2331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2262_ _2262_/A _2262_/B _2264_/B vssd1 vssd1 vccd1 vccd1 _2263_/A sky130_fd_sc_hd__and3_1
X_1213_ _2308_/Q _1239_/B vssd1 vssd1 vccd1 vccd1 _1587_/B sky130_fd_sc_hd__and2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2193_ _2193_/A vssd1 vssd1 vccd1 vccd1 _2440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1144_ _2442_/Q _1150_/B vssd1 vssd1 vccd1 vccd1 _1145_/A sky130_fd_sc_hd__and2_2
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1977_ _1126_/A _1976_/X _1940_/X vssd1 vssd1 vccd1 vccd1 _1977_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_162_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput307 wb_sel_i[2] vssd1 vssd1 vccd1 vccd1 _1551_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1900_ _1123_/A _2342_/Q _1904_/S vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__mux2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ _1831_/A _2332_/Q _2333_/Q _2334_/Q vssd1 vssd1 vccd1 vccd1 _1836_/C sky130_fd_sc_hd__and4_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1762_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1763_/A sky130_fd_sc_hd__inv_2
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1693_ _2420_/Q _1692_/Y _1671_/X _2417_/Q vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__o22a_1
XFILLER_171_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2315_/CLK _2314_/D vssd1 vssd1 vccd1 vccd1 _2314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2245_ _2245_/A vssd1 vssd1 vccd1 vccd1 _2462_/D sky130_fd_sc_hd__clkbuf_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2176_ _2432_/Q _2163_/X _2175_/Y vssd1 vssd1 vccd1 vccd1 _2432_/D sky130_fd_sc_hd__o21a_1
X_1127_ _2439_/Q vssd1 vssd1 vccd1 vccd1 _2040_/A sky130_fd_sc_hd__inv_2
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput126 sram_dout0[98] vssd1 vssd1 vccd1 vccd1 _1412_/A1 sky130_fd_sc_hd__buf_2
Xinput115 sram_dout0[88] vssd1 vssd1 vccd1 vccd1 _1503_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput104 sram_dout0[78] vssd1 vssd1 vccd1 vccd1 _1460_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput137 sram_dout1[107] vssd1 vssd1 vccd1 vccd1 _1327_/C sky130_fd_sc_hd__clkbuf_1
Xinput159 sram_dout1[13] vssd1 vssd1 vccd1 vccd1 _1260_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput148 sram_dout1[117] vssd1 vssd1 vccd1 vccd1 _1288_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2030_ _2079_/A vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__buf_2
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1814_ _2377_/Q vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__inv_2
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1745_ _1735_/Y _1681_/X _1738_/X _1741_/X _1744_/X vssd1 vssd1 vccd1 vccd1 _1745_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_171_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1676_ _2413_/Q _1828_/C vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__xor2_1
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _2228_/A vssd1 vssd1 vccd1 vccd1 _2456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2159_ _2046_/A _2158_/B _2158_/Y _2116_/X vssd1 vssd1 vccd1 vccd1 _2426_/D sky130_fd_sc_hd__a211o_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput408 _1524_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1530_ _2162_/A vssd1 vssd1 vccd1 vccd1 _1530_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1461_ input13/X _1443_/X _1447_/X _1460_/X vssd1 vssd1 vccd1 vccd1 _1461_/X sky130_fd_sc_hd__a211o_2
X_1392_ _1386_/B _1392_/B _1392_/C vssd1 vssd1 vccd1 vccd1 _1480_/A sky130_fd_sc_hd__and3b_2
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2013_ _2013_/A _2013_/B vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1728_ _1839_/A vssd1 vssd1 vccd1 vccd1 _1728_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1659_ _1664_/A _1663_/B _1659_/C vssd1 vssd1 vccd1 vccd1 _1660_/A sky130_fd_sc_hd__and3_1
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2316_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1513_ input27/X _1443_/A _1478_/X _1512_/X vssd1 vssd1 vccd1 vccd1 _1513_/X sky130_fd_sc_hd__a211o_2
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1444_ input65/X _1409_/X _1410_/X _1444_/B2 vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1375_ _1375_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1376_/A sky130_fd_sc_hd__and2_1
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1160_ _2303_/Q _1621_/B _1168_/S vssd1 vssd1 vccd1 vccd1 _1161_/A sky130_fd_sc_hd__mux2_2
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1993_ _1958_/X _1986_/X _1940_/X vssd1 vssd1 vccd1 vccd1 _1993_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1427_ input96/X _1400_/X _1426_/X _1404_/X vssd1 vssd1 vccd1 vccd1 _1427_/X sky130_fd_sc_hd__a211o_1
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1358_ _1358_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1359_/A sky130_fd_sc_hd__and2_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1289_ _1289_/A1 _1321_/B _1224_/X _1289_/B2 _1288_/X vssd1 vssd1 vccd1 vccd1 _1289_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2330_ _2474_/A _2330_/D vssd1 vssd1 vccd1 vccd1 _2330_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2261_ _2261_/A _2267_/D vssd1 vssd1 vccd1 vccd1 _2264_/B sky130_fd_sc_hd__nand2_1
X_1212_ _2307_/Q _2306_/Q vssd1 vssd1 vccd1 vccd1 _1239_/B sky130_fd_sc_hd__nor2_1
X_2192_ _2440_/Q _2192_/A1 _2198_/S vssd1 vssd1 vccd1 vccd1 _2193_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1143_ _1537_/B vssd1 vssd1 vccd1 vccd1 _1150_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1976_ _1976_/A vssd1 vssd1 vccd1 vccd1 _1976_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput308 wb_sel_i[3] vssd1 vssd1 vccd1 vccd1 _1553_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2459_ _2459_/CLK _2459_/D vssd1 vssd1 vccd1 vccd1 _2459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _1846_/A _1830_/B _1830_/C vssd1 vssd1 vccd1 vccd1 _2333_/D sky130_fd_sc_hd__nor3_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1761_ _1761_/A _1761_/B _1761_/C _1761_/D vssd1 vssd1 vccd1 vccd1 _1825_/A sky130_fd_sc_hd__or4_1
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1692_ _2336_/Q vssd1 vssd1 vccd1 vccd1 _1692_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2315_/CLK _2313_/D vssd1 vssd1 vccd1 vccd1 _2313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2475_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2244_ _2262_/A _2248_/B _2244_/C vssd1 vssd1 vccd1 vccd1 _2245_/A sky130_fd_sc_hd__and3_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2175_ _1107_/A _2164_/X _2185_/A vssd1 vssd1 vccd1 vccd1 _2175_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1126_ _1126_/A vssd1 vssd1 vccd1 vccd1 _1126_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1959_ _1958_/X _1957_/A _1940_/X vssd1 vssd1 vccd1 vccd1 _1959_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput127 sram_dout0[99] vssd1 vssd1 vccd1 vccd1 _1415_/A1 sky130_fd_sc_hd__buf_2
XFILLER_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput116 sram_dout0[89] vssd1 vssd1 vccd1 vccd1 _1506_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput105 sram_dout0[79] vssd1 vssd1 vccd1 vccd1 _1465_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput138 sram_dout1[108] vssd1 vssd1 vccd1 vccd1 _1226_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput149 sram_dout1[118] vssd1 vssd1 vccd1 vccd1 _1301_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1813_ _2467_/Q vssd1 vssd1 vccd1 vccd1 _2267_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1744_ _2402_/Q _1699_/Y _1671_/X _2397_/Q _1743_/Y vssd1 vssd1 vccd1 vccd1 _1744_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1675_ _2333_/Q vssd1 vssd1 vccd1 vccd1 _1828_/C sky130_fd_sc_hd__buf_2
XFILLER_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2227_ _2456_/Q _2227_/A1 _2231_/S vssd1 vssd1 vccd1 vccd1 _2228_/A sky130_fd_sc_hd__mux2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2158_ _2158_/A _2158_/B vssd1 vssd1 vccd1 vccd1 _2158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1109_ _1109_/A _1118_/B vssd1 vssd1 vccd1 vccd1 _2093_/A sky130_fd_sc_hd__nand2_8
X_2089_ _2089_/A _2100_/B vssd1 vssd1 vccd1 vccd1 _2089_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput409 _1527_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[31] sky130_fd_sc_hd__buf_2
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1460_ input69/X _1448_/X _1449_/X _1460_/B2 vssd1 vssd1 vccd1 vccd1 _1460_/X sky130_fd_sc_hd__a22o_1
X_1391_ _1479_/A vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2012_ _2374_/Q _2013_/B _2011_/Y vssd1 vssd1 vccd1 vccd1 _2374_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1727_ _1727_/A vssd1 vssd1 vccd1 vccd1 _2328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1658_ _1657_/A _2321_/Q _2322_/Q vssd1 vssd1 vccd1 vccd1 _1659_/C sky130_fd_sc_hd__a21o_1
XFILLER_132_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1589_ _1602_/B vssd1 vssd1 vccd1 vccd1 _1656_/B sky130_fd_sc_hd__buf_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1512_ input83/X _1479_/X _1480_/X _1512_/B2 vssd1 vssd1 vccd1 vccd1 _1512_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1443_ _1443_/A vssd1 vssd1 vccd1 vccd1 _1443_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1374_ _1374_/A vssd1 vssd1 vccd1 vccd1 _1374_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1992_ _1117_/X _1984_/X _1991_/X vssd1 vssd1 vccd1 vccd1 _2367_/D sky130_fd_sc_hd__a21o_1
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2475_ _2475_/A vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__buf_2
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1426_ input4/X _1425_/X _1402_/X input60/X vssd1 vssd1 vccd1 vccd1 _1426_/X sky130_fd_sc_hd__a22o_1
X_1357_ _1357_/A vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1288_ _1329_/A _1329_/B _1288_/C vssd1 vssd1 vccd1 vccd1 _1288_/X sky130_fd_sc_hd__and3_1
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2260_ _2261_/A _2267_/D vssd1 vssd1 vccd1 vccd1 _2262_/B sky130_fd_sc_hd__or2_1
X_1211_ _1200_/X _1206_/X _1208_/X _1210_/X vssd1 vssd1 vccd1 vccd1 _1231_/A sky130_fd_sc_hd__a22o_1
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2191_ _2191_/A vssd1 vssd1 vccd1 vccd1 _2439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1142_ _1392_/B vssd1 vssd1 vccd1 vccd1 _1537_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1975_ _2042_/A _2052_/B _2109_/B vssd1 vssd1 vccd1 vccd1 _1976_/A sky130_fd_sc_hd__nor3_1
XFILLER_174_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2458_ _2474_/A _2458_/D vssd1 vssd1 vccd1 vccd1 _2458_/Q sky130_fd_sc_hd__dfxtp_1
Xinput309 wb_stb_i vssd1 vssd1 vccd1 vccd1 _1544_/D sky130_fd_sc_hd__clkbuf_2
X_1409_ _1479_/A vssd1 vssd1 vccd1 vccd1 _1409_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2389_ _2435_/CLK _2389_/D vssd1 vssd1 vccd1 vccd1 _2389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1760_ _2434_/Q _1683_/Y _1672_/Y _2426_/Q _1759_/X vssd1 vssd1 vccd1 vccd1 _1761_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1691_ _1691_/A _1691_/B _1691_/C _1690_/X vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__or4b_1
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2312_ _2315_/CLK _2312_/D vssd1 vssd1 vccd1 vccd1 _2312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2243_ _2243_/A _2243_/B vssd1 vssd1 vccd1 vccd1 _2244_/C sky130_fd_sc_hd__nand2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ _1111_/X _2163_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _2431_/D sky130_fd_sc_hd__a21o_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1125_ _1125_/A _1366_/A vssd1 vssd1 vccd1 vccd1 _1126_/A sky130_fd_sc_hd__nand2_2
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1958_ _2171_/A vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__buf_4
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1889_ _2071_/A vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput117 sram_dout0[8] vssd1 vssd1 vccd1 vccd1 _1437_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput106 sram_dout0[7] vssd1 vssd1 vccd1 vccd1 _1431_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput139 sram_dout1[109] vssd1 vssd1 vccd1 vccd1 _1254_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput128 sram_dout0[9] vssd1 vssd1 vccd1 vccd1 _1441_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1812_ _2275_/A _2374_/Q _2013_/A _2272_/A vssd1 vssd1 vccd1 vccd1 _1818_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1743_ _1730_/Y _1749_/B _1742_/X vssd1 vssd1 vccd1 vccd1 _1743_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1674_ _2407_/Q _1671_/X _1672_/Y _2406_/Q _1673_/X vssd1 vssd1 vccd1 vccd1 _1674_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2226_ _2226_/A vssd1 vssd1 vccd1 vccd1 _2455_/D sky130_fd_sc_hd__clkbuf_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2157_ _2157_/A _2167_/B _2157_/C vssd1 vssd1 vccd1 vccd1 _2158_/B sky130_fd_sc_hd__nor3_4
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1108_ _1926_/A vssd1 vssd1 vccd1 vccd1 _1108_/X sky130_fd_sc_hd__buf_6
X_2088_ _2102_/B vssd1 vssd1 vccd1 vccd1 _2100_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _2448_/Q _2447_/Q _1531_/B vssd1 vssd1 vccd1 vccd1 _1479_/A sky130_fd_sc_hd__and3b_4
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2011_ _1126_/A _2013_/B _1995_/X vssd1 vssd1 vccd1 vccd1 _2011_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1726_ _1726_/A _1726_/B _1726_/C vssd1 vssd1 vccd1 vccd1 _1727_/A sky130_fd_sc_hd__and3_1
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1657_ _1657_/A _2321_/Q _2322_/Q vssd1 vssd1 vccd1 vccd1 _1663_/B sky130_fd_sc_hd__nand3_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1588_ _2341_/Q vssd1 vssd1 vccd1 vccd1 _1613_/A sky130_fd_sc_hd__buf_2
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2209_ _1392_/C _2209_/A1 _2209_/S vssd1 vssd1 vccd1 vccd1 _2210_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1511_ input47/X _1505_/X _1501_/X _1510_/X vssd1 vssd1 vccd1 vccd1 _1511_/X sky130_fd_sc_hd__o211a_4
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1442_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1442_/X sky130_fd_sc_hd__buf_2
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1373_ _1373_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1374_/A sky130_fd_sc_hd__and2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1709_ _2425_/Q _1698_/Y _2336_/Q _1708_/Y vssd1 vssd1 vccd1 vccd1 _1710_/D sky130_fd_sc_hd__o22a_1
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ _2367_/Q _1990_/X _1966_/X vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2474_ _2474_/A vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__buf_2
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1425_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1356_ _1356_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1357_/A sky130_fd_sc_hd__and2_1
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1287_ _1287_/A vssd1 vssd1 vccd1 vccd1 _1321_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1210_ _1210_/A1 _1191_/A _1195_/A _1210_/B2 _1209_/X vssd1 vssd1 vccd1 vccd1 _1210_/X
+ sky130_fd_sc_hd__a221o_1
X_2190_ _2439_/Q _2190_/A1 _2198_/S vssd1 vssd1 vccd1 vccd1 _2191_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1141_ _1531_/B vssd1 vssd1 vccd1 vccd1 _1392_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _2439_/Q _2040_/B _2040_/C vssd1 vssd1 vccd1 vccd1 _2109_/B sky130_fd_sc_hd__or3_4
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2457_ _2474_/A _2457_/D vssd1 vssd1 vccd1 vccd1 _2457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1408_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1408_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2388_ _2435_/CLK _2388_/D vssd1 vssd1 vccd1 vccd1 _2388_/Q sky130_fd_sc_hd__dfxtp_1
X_1339_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1339_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput390 _1462_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1690_ _2121_/A _1836_/A _1671_/X _2407_/Q _1689_/Y vssd1 vssd1 vccd1 vccd1 _1690_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2311_ _2315_/CLK _2311_/D vssd1 vssd1 vccd1 vccd1 _2311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2242_ _2243_/A _2243_/B vssd1 vssd1 vccd1 vccd1 _2248_/B sky130_fd_sc_hd__or2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2173_ _2431_/Q _2171_/B _1889_/X vssd1 vssd1 vccd1 vccd1 _2173_/X sky130_fd_sc_hd__a21o_1
X_1124_ _2046_/A vssd1 vssd1 vccd1 vccd1 _1124_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1888_ _1952_/A vssd1 vssd1 vccd1 vccd1 _2071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput118 sram_dout0[90] vssd1 vssd1 vccd1 vccd1 _1509_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput107 sram_dout0[80] vssd1 vssd1 vccd1 vccd1 _1467_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput129 sram_dout1[0] vssd1 vssd1 vccd1 vccd1 _1246_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1811_ _2375_/Q vssd1 vssd1 vccd1 vccd1 _2013_/A sky130_fd_sc_hd__inv_2
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1742_ _2400_/Q _1692_/Y _1728_/Y _2399_/Q vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__o22a_1
X_1673_ _2410_/Q _2336_/Q vssd1 vssd1 vccd1 vccd1 _1673_/X sky130_fd_sc_hd__xor2_1
XFILLER_144_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2225_ _2455_/Q _2225_/A1 _2231_/S vssd1 vssd1 vccd1 vccd1 _2226_/A sky130_fd_sc_hd__mux2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2156_ _2425_/Q _2137_/X _2155_/Y vssd1 vssd1 vccd1 vccd1 _2425_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1107_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__inv_2
X_2087_ _1730_/Y _2084_/X _2086_/X vssd1 vssd1 vccd1 vccd1 _2398_/D sky130_fd_sc_hd__a21oi_1
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ _2010_/A vssd1 vssd1 vccd1 vccd1 _2013_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1725_ _1725_/A _1725_/B vssd1 vssd1 vccd1 vccd1 _1726_/C sky130_fd_sc_hd__or2_1
XFILLER_172_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1656_ _1656_/A _1656_/B vssd1 vssd1 vccd1 vccd1 _1664_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1587_ _2302_/Q _1587_/B _1602_/B vssd1 vssd1 vccd1 vccd1 _1596_/C sky130_fd_sc_hd__and3_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _2208_/A vssd1 vssd1 vccd1 vccd1 _2447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2139_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1510_ input26/X _1473_/X _1478_/X _1509_/X vssd1 vssd1 vccd1 vccd1 _1510_/X sky130_fd_sc_hd__a211o_2
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1441_ _1441_/A1 _1421_/X _1438_/X _1440_/X vssd1 vssd1 vccd1 vccd1 _1441_/X sky130_fd_sc_hd__o211a_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1372_ _1372_/A vssd1 vssd1 vccd1 vccd1 _1372_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput290 wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1708_ _2420_/Q vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__inv_2
X_1639_ _1639_/A _1641_/C vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__or2_1
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ _2136_/A _2042_/B _2109_/B vssd1 vssd1 vccd1 vccd1 _1990_/X sky130_fd_sc_hd__or3_4
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2468_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1424_ input84/X _1421_/X _1417_/X _1423_/X vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__o211a_4
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1355_ _1379_/B vssd1 vssd1 vccd1 vccd1 _1364_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1286_ _1286_/A1 _1200_/X _1208_/X _1286_/B2 _1285_/X vssd1 vssd1 vccd1 vccd1 _1286_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1140_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1140_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ _2057_/B vssd1 vssd1 vccd1 vccd1 _2052_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_174_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2456_ _2459_/CLK _2456_/D vssd1 vssd1 vccd1 vccd1 _2456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1407_ _1473_/A vssd1 vssd1 vccd1 vccd1 _1407_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2387_ _2435_/CLK _2387_/D vssd1 vssd1 vccd1 vccd1 _2387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1338_ _1338_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _1339_/A sky130_fd_sc_hd__and2_1
X_1269_ _1233_/X _1266_/X _1268_/X _1208_/X vssd1 vssd1 vccd1 vccd1 _1275_/A sky130_fd_sc_hd__a22o_1
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput380 _2330_/Q vssd1 vssd1 vccd1 vccd1 vga_hsync sky130_fd_sc_hd__buf_2
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput391 _1466_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2310_ _2316_/CLK _2310_/D vssd1 vssd1 vccd1 vccd1 _2310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2273_/A vssd1 vssd1 vccd1 vccd1 _2262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2172_ _2430_/Q _2171_/B _2171_/Y _1919_/X vssd1 vssd1 vccd1 vccd1 _2430_/D sky130_fd_sc_hd__a211o_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1123_ _1123_/A vssd1 vssd1 vccd1 vccd1 _2046_/A sky130_fd_sc_hd__buf_4
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1956_ _1869_/Y _1950_/X _1955_/X vssd1 vssd1 vccd1 vccd1 _2356_/D sky130_fd_sc_hd__a21oi_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1887_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1952_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput108 sram_dout0[81] vssd1 vssd1 vccd1 vccd1 _1471_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput119 sram_dout0[91] vssd1 vssd1 vccd1 vccd1 _1512_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2439_ _2446_/CLK _2439_/D vssd1 vssd1 vccd1 vccd1 _2439_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _1807_/Y _2238_/A _2275_/A _2374_/Q _1809_/X vssd1 vssd1 vccd1 vccd1 _1818_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1741_ _2405_/Q _1698_/Y _1739_/Y _2401_/Q _1740_/Y vssd1 vssd1 vccd1 vccd1 _1741_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1672_ _2340_/Q vssd1 vssd1 vccd1 vccd1 _1672_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2224_/A vssd1 vssd1 vccd1 vccd1 _2454_/D sky130_fd_sc_hd__clkbuf_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2155_ _2102_/A _2138_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _2155_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1106_ _1106_/A _1122_/B vssd1 vssd1 vccd1 vccd1 _1107_/A sky130_fd_sc_hd__nand2_8
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2086_ _1985_/A _2085_/Y _1952_/X vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _1952_/A vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput90 sram_dout0[65] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1724_ _1725_/A _1725_/B vssd1 vssd1 vccd1 vccd1 _1726_/B sky130_fd_sc_hd__nand2_1
XFILLER_172_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1655_ _1657_/A _2321_/Q _1654_/Y vssd1 vssd1 vccd1 vccd1 _2321_/D sky130_fd_sc_hd__o21a_1
X_1586_ _1586_/A _1586_/B _1586_/C _1586_/D vssd1 vssd1 vccd1 vccd1 _1602_/B sky130_fd_sc_hd__and4_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _1386_/B _2207_/A1 _2209_/S vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2069_ _2394_/Q _2058_/X _2037_/X vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1440_ input7/X _1407_/X _1408_/X _1439_/X vssd1 vssd1 vccd1 vccd1 _1440_/X sky130_fd_sc_hd__a211o_2
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1371_ _1371_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1372_/A sky130_fd_sc_hd__and2_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput280 wb_data_i[17] vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput291 wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _1371_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1707_ _2417_/Q _1671_/A _1740_/B _2423_/Q vssd1 vssd1 vccd1 vccd1 _1710_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1638_ _1639_/A _1641_/C vssd1 vssd1 vccd1 vccd1 _1638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1569_ _2297_/Q _1567_/A _1562_/X vssd1 vssd1 vccd1 vccd1 _1570_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2472_ _2472_/CLK _2472_/D vssd1 vssd1 vccd1 vccd1 _2472_/Q sky130_fd_sc_hd__dfxtp_1
X_1423_ input94/X _1400_/X _1422_/X _1404_/X vssd1 vssd1 vccd1 vccd1 _1423_/X sky130_fd_sc_hd__a211o_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1354_ _1354_/A vssd1 vssd1 vccd1 vccd1 _1354_/X sky130_fd_sc_hd__clkbuf_1
X_1285_ _1285_/A1 _1284_/X _1223_/X _1285_/B2 vssd1 vssd1 vccd1 vccd1 _1285_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1972_ _1098_/X _1957_/A _1971_/X vssd1 vssd1 vccd1 vccd1 _2362_/D sky130_fd_sc_hd__a21o_1
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2455_ _2459_/CLK _2455_/D vssd1 vssd1 vccd1 vccd1 _2455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1406_ input40/X _1385_/X _1398_/X _1405_/X vssd1 vssd1 vccd1 vccd1 _1406_/X sky130_fd_sc_hd__o211a_4
X_2386_ _2435_/CLK _2386_/D vssd1 vssd1 vccd1 vccd1 _2386_/Q sky130_fd_sc_hd__dfxtp_1
X_1337_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1337_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1268_ _1268_/A1 _1191_/A _1195_/A _1268_/B2 _1267_/X vssd1 vssd1 vccd1 vccd1 _1268_/X
+ sky130_fd_sc_hd__a221o_1
X_1199_ _1609_/A _1609_/B _1602_/A vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__nor3b_2
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput370 _1124_/X vssd1 vssd1 vccd1 vccd1 sram_din0[9] sky130_fd_sc_hd__buf_2
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput392 _1469_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput381 _1247_/X vssd1 vssd1 vccd1 vccd1 vga_r[0] sky130_fd_sc_hd__buf_2
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2240_/A vssd1 vssd1 vccd1 vccd1 _2461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2171_ _2171_/A _2171_/B vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__nor2_1
X_1122_ _1122_/A _1122_/B vssd1 vssd1 vccd1 vccd1 _1123_/A sky130_fd_sc_hd__and2_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1955_ _2089_/A _1957_/A _1952_/X vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1886_ _1656_/A _2239_/A _1873_/X _1885_/X vssd1 vssd1 vccd1 vccd1 _2341_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_174_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput109 sram_dout0[82] vssd1 vssd1 vccd1 vccd1 _1474_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2438_ _2446_/CLK _2438_/D vssd1 vssd1 vccd1 vccd1 _2438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2369_ _2474_/A _2369_/D vssd1 vssd1 vccd1 vccd1 _2369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1740_ _2403_/Q _1740_/B vssd1 vssd1 vccd1 vccd1 _1740_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1671_ _1671_/A vssd1 vssd1 vccd1 vccd1 _1671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2223_ _2454_/Q _2223_/A1 _2231_/S vssd1 vssd1 vccd1 vccd1 _2224_/A sky130_fd_sc_hd__mux2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2154_ _2424_/Q _2137_/X _2153_/Y vssd1 vssd1 vccd1 vccd1 _2424_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1105_ _1105_/A vssd1 vssd1 vccd1 vccd1 _1105_/X sky130_fd_sc_hd__buf_4
X_2085_ _2162_/A _2085_/B _2157_/C vssd1 vssd1 vccd1 vccd1 _2085_/Y sky130_fd_sc_hd__nor3_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1938_ _1938_/A vssd1 vssd1 vccd1 vccd1 _1943_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1869_ _2356_/Q vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput91 sram_dout0[66] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput80 sram_dout0[56] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1723_ _2328_/Q vssd1 vssd1 vccd1 vccd1 _1725_/A sky130_fd_sc_hd__inv_2
XFILLER_8_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1654_ _1657_/A _2321_/Q _1653_/B vssd1 vssd1 vccd1 vccd1 _1654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1585_ _2349_/Q _2322_/Q vssd1 vssd1 vccd1 vccd1 _1586_/D sky130_fd_sc_hd__xnor2_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2137_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ _1105_/X _2054_/X _2067_/X vssd1 vssd1 vccd1 vccd1 _2393_/D sky130_fd_sc_hd__a21o_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_167_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1370_ _1370_/A vssd1 vssd1 vccd1 vccd1 _1370_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput270 wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 _2203_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput281 wb_data_i[18] vssd1 vssd1 vccd1 vccd1 _1351_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput292 wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _1373_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1706_ _2422_/Q _1699_/Y _1672_/Y _2416_/Q _1705_/Y vssd1 vssd1 vccd1 vccd1 _1710_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1637_ _1615_/X _1635_/Y _1636_/X _1622_/X _2315_/Q vssd1 vssd1 vccd1 vccd1 _2315_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1568_ _2297_/Q _2296_/Q _2295_/Q _1568_/D vssd1 vssd1 vccd1 vccd1 _1577_/D sky130_fd_sc_hd__and4_1
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1499_ input22/X _1473_/X _1478_/X _1498_/X vssd1 vssd1 vccd1 vccd1 _1499_/X sky130_fd_sc_hd__a211o_2
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2471_ _2472_/CLK _2471_/D vssd1 vssd1 vccd1 vccd1 _2471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1422_ input3/X _1473_/A _1402_/X input59/X vssd1 vssd1 vccd1 vccd1 _1422_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1353_ _1353_/A _1353_/B vssd1 vssd1 vccd1 vccd1 _1354_/A sky130_fd_sc_hd__and2_1
X_1284_ _1587_/B vssd1 vssd1 vccd1 vccd1 _1284_/X sky130_fd_sc_hd__buf_2
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1971_ _2362_/Q _1950_/A _1966_/X vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2454_ _2459_/CLK _2454_/D vssd1 vssd1 vccd1 vccd1 _2454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1405_ input90/X _1400_/X _1403_/X _1404_/X vssd1 vssd1 vccd1 vccd1 _1405_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2385_ _2435_/CLK _2385_/D vssd1 vssd1 vccd1 vccd1 _2385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1336_ _1336_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _1337_/A sky130_fd_sc_hd__and2_1
Xinput1 sram_dout0[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_1267_ _1303_/A _1303_/B _1267_/C vssd1 vssd1 vccd1 vccd1 _1267_/X sky130_fd_sc_hd__and3_1
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1198_ _2306_/Q vssd1 vssd1 vccd1 vccd1 _1602_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput371 _1140_/Y vssd1 vssd1 vccd1 vccd1 sram_web0 sky130_fd_sc_hd__buf_2
Xoutput360 _1376_/X vssd1 vssd1 vccd1 vccd1 sram_din0[29] sky130_fd_sc_hd__buf_2
XFILLER_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput382 _1264_/X vssd1 vssd1 vccd1 vccd1 vga_r[1] sky130_fd_sc_hd__buf_2
Xoutput393 _1472_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2170_ _1117_/X _2163_/X _2169_/X vssd1 vssd1 vccd1 vccd1 _2429_/D sky130_fd_sc_hd__a21o_1
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1121_ _2049_/A vssd1 vssd1 vccd1 vccd1 _1121_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1954_ _1877_/Y _1950_/X _1953_/X vssd1 vssd1 vccd1 vccd1 _2355_/D sky130_fd_sc_hd__a21oi_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1885_ _1885_/A _1885_/B _1885_/C _1884_/X vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__or4b_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2437_ _2472_/CLK _2437_/D vssd1 vssd1 vccd1 vccd1 _2437_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2368_ _2459_/CLK _2368_/D vssd1 vssd1 vccd1 vccd1 _2368_/Q sky130_fd_sc_hd__dfxtp_1
X_1319_ _1319_/A1 _1284_/X _1235_/X _1319_/B2 vssd1 vssd1 vccd1 vccd1 _1319_/X sky130_fd_sc_hd__a22o_1
X_2299_ _2319_/CLK _2299_/D vssd1 vssd1 vccd1 vccd1 _2299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1670_ _2339_/Q vssd1 vssd1 vccd1 vccd1 _1671_/A sky130_fd_sc_hd__inv_2
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2222_ _2222_/A vssd1 vssd1 vccd1 vccd1 _2231_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2153_ _2100_/A _2138_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _2153_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1104_ _2098_/A vssd1 vssd1 vccd1 vccd1 _1105_/A sky130_fd_sc_hd__inv_2
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2084_ _2102_/B vssd1 vssd1 vccd1 vccd1 _2084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1937_ _2042_/A _2085_/B _2042_/B vssd1 vssd1 vccd1 vccd1 _1938_/A sky130_fd_sc_hd__nor3_1
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1868_ _2273_/A vssd1 vssd1 vccd1 vccd1 _2239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput81 sram_dout0[57] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_1
Xinput70 sram_dout0[47] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
Xinput92 sram_dout0[67] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1799_ _2463_/Q vssd1 vssd1 vccd1 vccd1 _1800_/A sky130_fd_sc_hd__inv_2
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1722_ _1722_/A vssd1 vssd1 vccd1 vccd1 _2327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1653_ _1657_/A _1653_/B vssd1 vssd1 vccd1 vccd1 _2320_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1584_ _2351_/Q _2320_/Q vssd1 vssd1 vccd1 vccd1 _1586_/C sky130_fd_sc_hd__xnor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2446_/Q _2205_/A1 _2209_/S vssd1 vssd1 vccd1 vccd1 _2206_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2136_ _2136_/A _2142_/B _2162_/C vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__nor3_2
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2067_ _2393_/Q _2058_/X _2037_/X vssd1 vssd1 vccd1 vccd1 _2067_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput271 wb_cyc_i vssd1 vssd1 vccd1 vccd1 _1544_/C sky130_fd_sc_hd__buf_2
Xinput260 wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 _2229_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput282 wb_data_i[19] vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput293 wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1705_ _2419_/Q _1839_/A vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1636_ _1629_/A _2314_/Q _1634_/D _2315_/Q vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__a31o_1
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1567_ _1567_/A _1567_/B vssd1 vssd1 vccd1 vccd1 _2296_/D sky130_fd_sc_hd__nor2_1
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1498_ input79/X _1479_/X _1480_/X _1498_/B2 vssd1 vssd1 vccd1 vccd1 _1498_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2119_ _2171_/A _2112_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _2119_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2470_ _2474_/A _2470_/D vssd1 vssd1 vccd1 vccd1 _2470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1421_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1421_/X sky130_fd_sc_hd__buf_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1352_ _1352_/A vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__clkbuf_1
X_1283_ _1283_/A1 _1187_/Y _1191_/Y _1283_/B2 vssd1 vssd1 vccd1 vccd1 _1283_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1619_ _1650_/A _1619_/B vssd1 vssd1 vccd1 vccd1 _2310_/D sky130_fd_sc_hd__nor2_1
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1970_ _1102_/X _1957_/X _1969_/X vssd1 vssd1 vccd1 vccd1 _2361_/D sky130_fd_sc_hd__a21o_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2453_ _2459_/CLK _2453_/D vssd1 vssd1 vccd1 vccd1 _2453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1404_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1404_/X sky130_fd_sc_hd__buf_2
X_2384_ _2474_/A _2384_/D vssd1 vssd1 vccd1 vccd1 _2384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1335_ _1366_/A vssd1 vssd1 vccd1 vccd1 _1342_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput2 sram_dout0[100] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1266_ _1266_/A1 _1201_/X _1202_/X _1266_/B2 _1265_/X vssd1 vssd1 vccd1 vccd1 _1266_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1197_ _2307_/Q vssd1 vssd1 vccd1 vccd1 _1609_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput350 _1102_/X vssd1 vssd1 vccd1 vccd1 sram_din0[1] sky130_fd_sc_hd__buf_2
Xoutput361 _1105_/X vssd1 vssd1 vccd1 vccd1 sram_din0[2] sky130_fd_sc_hd__buf_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput372 _1530_/Y vssd1 vssd1 vccd1 vccd1 sram_wmask0[0] sky130_fd_sc_hd__buf_2
Xoutput394 _1476_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput383 _2324_/Q vssd1 vssd1 vccd1 vccd1 vga_vsync sky130_fd_sc_hd__buf_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2435_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1120_ _1120_/A _1122_/B vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1953_ _1985_/A _1957_/A _1952_/X vssd1 vssd1 vccd1 vccd1 _1953_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1884_ _2359_/Q _2248_/A _1794_/X _2358_/Q _1883_/X vssd1 vssd1 vccd1 vccd1 _1884_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2436_ _2446_/CLK _2436_/D vssd1 vssd1 vccd1 vccd1 _2436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2367_ _2474_/A _2367_/D vssd1 vssd1 vccd1 vccd1 _2367_/Q sky130_fd_sc_hd__dfxtp_1
X_1318_ _1318_/A1 _1187_/Y _1195_/Y _1318_/B2 vssd1 vssd1 vccd1 vccd1 _1318_/X sky130_fd_sc_hd__o22a_1
X_2298_ _2319_/CLK _2298_/D vssd1 vssd1 vccd1 vccd1 _2298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1249_ _1303_/A _1301_/B _1249_/C vssd1 vssd1 vccd1 vccd1 _1249_/X sky130_fd_sc_hd__and3_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2453_/D sky130_fd_sc_hd__clkbuf_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2152_ _1105_/A _2138_/X _2151_/X vssd1 vssd1 vccd1 vccd1 _2423_/D sky130_fd_sc_hd__a21o_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1103_ _1103_/A _1118_/B vssd1 vssd1 vccd1 vccd1 _2098_/A sky130_fd_sc_hd__nand2_4
X_2083_ _2167_/A _2085_/B _2162_/C vssd1 vssd1 vccd1 vccd1 _2102_/B sky130_fd_sc_hd__or3_2
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1936_ _2057_/B vssd1 vssd1 vccd1 vccd1 _2042_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1867_ _1849_/X _1850_/Y _1853_/X _1866_/X vssd1 vssd1 vccd1 vccd1 _2273_/A sky130_fd_sc_hd__a211o_1
XFILLER_174_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput82 sram_dout0[58] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
Xinput71 sram_dout0[48] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput60 sram_dout0[38] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
X_1798_ _1798_/A vssd1 vssd1 vccd1 vccd1 _2257_/A sky130_fd_sc_hd__buf_2
XFILLER_162_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput93 sram_dout0[68] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2419_ _2425_/CLK _2419_/D vssd1 vssd1 vccd1 vccd1 _2419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1721_ _1726_/A _1725_/B _1721_/C vssd1 vssd1 vccd1 vccd1 _1722_/A sky130_fd_sc_hd__and3_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1652_ _1656_/A _1656_/B vssd1 vssd1 vccd1 vccd1 _1653_/B sky130_fd_sc_hd__or2_1
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1583_ _2350_/Q _2321_/Q vssd1 vssd1 vccd1 vccd1 _1586_/B sky130_fd_sc_hd__xnor2_1
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2204_/A vssd1 vssd1 vccd1 vccd1 _2445_/D sky130_fd_sc_hd__clkbuf_1
X_2135_ _2417_/Q _2132_/B _2134_/Y vssd1 vssd1 vccd1 vccd1 _2417_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2066_ _1108_/X _2054_/X _2065_/X vssd1 vssd1 vccd1 vccd1 _2392_/D sky130_fd_sc_hd__a21o_1
XFILLER_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1919_ _2139_/A vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput272 wb_data_i[0] vssd1 vssd1 vccd1 vccd1 _1096_/A sky130_fd_sc_hd__buf_2
Xinput250 wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 _2207_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput261 wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 _2231_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput294 wb_data_i[2] vssd1 vssd1 vccd1 vccd1 _1103_/A sky130_fd_sc_hd__clkbuf_2
Xinput283 wb_data_i[1] vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__buf_2
XFILLER_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1704_ _2423_/Q _1740_/B _1696_/Y _2418_/Q _1703_/X vssd1 vssd1 vccd1 vccd1 _1704_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1635_ _1641_/C vssd1 vssd1 vccd1 vccd1 _1635_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1566_ _2296_/Q _1564_/A _1562_/X vssd1 vssd1 vccd1 vccd1 _1567_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1497_ input43/X _1484_/X _1477_/X _1496_/X vssd1 vssd1 vccd1 vccd1 _1497_/X sky130_fd_sc_hd__o211a_4
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2118_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2049_ _2049_/A vssd1 vssd1 vccd1 vccd1 _2049_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1420_ input73/X _1385_/X _1417_/X _1419_/X vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__o211a_4
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1351_ _1351_/A _1353_/B vssd1 vssd1 vccd1 vccd1 _1352_/A sky130_fd_sc_hd__and2_1
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1282_ _1282_/A1 _1195_/Y _1281_/X _1282_/B2 vssd1 vssd1 vccd1 vccd1 _1282_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1618_ _1621_/B _1618_/B vssd1 vssd1 vccd1 vccd1 _1619_/B sky130_fd_sc_hd__xnor2_1
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1549_ _2281_/Q _1549_/A1 _2187_/S vssd1 vssd1 vccd1 vccd1 _1550_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2452_ _2452_/CLK _2452_/D vssd1 vssd1 vccd1 vccd1 _2452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1403_ _1403_/A1 _1473_/A _1402_/X input55/X vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2383_ _2474_/A _2383_/D vssd1 vssd1 vccd1 vccd1 _2383_/Q sky130_fd_sc_hd__dfxtp_1
X_1334_ _1241_/A _1317_/X _1318_/X _1333_/X vssd1 vssd1 vccd1 vccd1 _1334_/X sky130_fd_sc_hd__a31o_4
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1265_ _1301_/A _1301_/B _1265_/C vssd1 vssd1 vccd1 vccd1 _1265_/X sky130_fd_sc_hd__and3_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 sram_dout0[101] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1196_ _2308_/Q vssd1 vssd1 vccd1 vccd1 _1609_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput340 _1126_/Y vssd1 vssd1 vccd1 vccd1 sram_din0[10] sky130_fd_sc_hd__buf_2
Xoutput351 _1357_/X vssd1 vssd1 vccd1 vccd1 sram_din0[20] sky130_fd_sc_hd__buf_2
Xoutput362 _1378_/X vssd1 vssd1 vccd1 vccd1 sram_din0[30] sky130_fd_sc_hd__buf_2
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput373 _1534_/Y vssd1 vssd1 vccd1 vccd1 sram_wmask0[1] sky130_fd_sc_hd__buf_2
Xoutput395 _1483_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput384 _2436_/Q vssd1 vssd1 vccd1 vccd1 wb_ack_o sky130_fd_sc_hd__buf_2
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _1952_/A vssd1 vssd1 vccd1 vccd1 _1952_/X sky130_fd_sc_hd__buf_2
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1883_ _1874_/Y _2238_/B _2267_/A _1869_/Y vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2435_ _2435_/CLK _2435_/D vssd1 vssd1 vccd1 vccd1 _2435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2366_ _2474_/A _2366_/D vssd1 vssd1 vccd1 vccd1 _2366_/Q sky130_fd_sc_hd__dfxtp_1
X_1317_ _1317_/A1 _1191_/Y _1281_/X _1317_/B2 vssd1 vssd1 vccd1 vccd1 _1317_/X sky130_fd_sc_hd__o22a_1
X_2297_ _2319_/CLK _2297_/D vssd1 vssd1 vccd1 vccd1 _2297_/Q sky130_fd_sc_hd__dfxtp_1
X_1248_ _1327_/B vssd1 vssd1 vccd1 vccd1 _1301_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1179_ _1179_/A vssd1 vssd1 vccd1 vccd1 _2292_/D sky130_fd_sc_hd__clkbuf_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2220_ _2453_/Q _2220_/A1 _2220_/S vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__mux2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2151_ _2423_/Q _2142_/X _2071_/X vssd1 vssd1 vccd1 vccd1 _2151_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1102_ _1930_/A vssd1 vssd1 vccd1 vccd1 _1102_/X sky130_fd_sc_hd__buf_4
X_2082_ _2167_/C vssd1 vssd1 vccd1 vccd1 _2162_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1935_ _1935_/A _1935_/B _2074_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _2057_/B sky130_fd_sc_hd__or4_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1866_ _1866_/A _1866_/B _1862_/X _1865_/X vssd1 vssd1 vccd1 vccd1 _1866_/X sky130_fd_sc_hd__or4bb_1
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput72 sram_dout0[49] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
Xinput61 sram_dout0[39] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
Xinput50 sram_dout0[29] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
X_1797_ _2465_/Q vssd1 vssd1 vccd1 vccd1 _1798_/A sky130_fd_sc_hd__inv_2
Xinput94 sram_dout0[69] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_2
Xinput83 sram_dout0[59] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2418_ _2435_/CLK _2418_/D vssd1 vssd1 vccd1 vccd1 _2418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2349_ _2414_/CLK _2349_/D vssd1 vssd1 vccd1 vccd1 _2349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1720_ _1719_/A _2326_/Q _2327_/Q vssd1 vssd1 vccd1 vccd1 _1721_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1651_ _2320_/Q vssd1 vssd1 vccd1 vccd1 _1657_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1582_ _2348_/Q _2323_/Q vssd1 vssd1 vccd1 vccd1 _1586_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2445_/Q _2203_/A1 _2209_/S vssd1 vssd1 vccd1 vccd1 _2204_/A sky130_fd_sc_hd__mux2_1
X_2134_ _2049_/X _2132_/B _2118_/X vssd1 vssd1 vccd1 vccd1 _2134_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2065_ _2392_/Q _2058_/X _2037_/X vssd1 vssd1 vccd1 vccd1 _2065_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1918_ _1930_/B vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__clkbuf_2
X_1849_ _2387_/Q _2468_/Q vssd1 vssd1 vccd1 vccd1 _1849_/X sky130_fd_sc_hd__or2_1
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput240 sram_dout1[90] vssd1 vssd1 vccd1 vccd1 _1273_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput251 wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 _2209_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput262 wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 _2233_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput295 wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _1377_/A sky130_fd_sc_hd__clkbuf_1
Xinput273 wb_data_i[10] vssd1 vssd1 vccd1 vccd1 _1125_/A sky130_fd_sc_hd__clkbuf_2
Xinput284 wb_data_i[20] vssd1 vssd1 vccd1 vccd1 _1356_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ _2421_/Q _1836_/A vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__xor2_1
XFILLER_172_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1634_ _2313_/Q _2314_/Q _2315_/Q _1634_/D vssd1 vssd1 vccd1 vccd1 _1641_/C sky130_fd_sc_hd__and4_1
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1565_ _2296_/Q _2295_/Q _1568_/D vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__and3_1
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1496_ _1496_/A1 _1489_/X _1495_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1496_/X sky130_fd_sc_hd__a211o_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2117_ _1117_/A _2112_/X _2115_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _2409_/D sky130_fd_sc_hd__a211o_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ _2386_/Q _2043_/X _2047_/Y vssd1 vssd1 vccd1 vccd1 _2386_/D sky130_fd_sc_hd__o21a_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_30 _1191_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1350_ _1350_/A vssd1 vssd1 vccd1 vccd1 _1350_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1281_ _1314_/A vssd1 vssd1 vccd1 vccd1 _1281_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1617_ _1621_/A _1615_/X _1618_/B vssd1 vssd1 vccd1 vccd1 _2309_/D sky130_fd_sc_hd__o21ba_1
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1548_ _1548_/A vssd1 vssd1 vccd1 vccd1 _2280_/D sky130_fd_sc_hd__clkbuf_1
X_1479_ _1479_/A vssd1 vssd1 vccd1 vccd1 _1479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2451_ _2452_/CLK _2451_/D vssd1 vssd1 vccd1 vccd1 _2451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1402_ _1479_/A vssd1 vssd1 vccd1 vccd1 _1402_/X sky130_fd_sc_hd__buf_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2382_ _2474_/A _2382_/D vssd1 vssd1 vccd1 vccd1 _2382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1333_ _1281_/X _1320_/X _1332_/X vssd1 vssd1 vccd1 vccd1 _1333_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1264_ _1259_/X _1262_/X _1263_/X _1241_/X vssd1 vssd1 vccd1 vccd1 _1264_/X sky130_fd_sc_hd__a22o_4
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 sram_dout0[102] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1195_ _1195_/A vssd1 vssd1 vccd1 vccd1 _1195_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput330 _2475_/X vssd1 vssd1 vccd1 vccd1 sram_clk1 sky130_fd_sc_hd__clkbuf_1
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput341 _1337_/X vssd1 vssd1 vccd1 vccd1 sram_din0[11] sky130_fd_sc_hd__buf_2
Xoutput352 _1359_/X vssd1 vssd1 vccd1 vccd1 sram_din0[21] sky130_fd_sc_hd__buf_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput374 _1536_/X vssd1 vssd1 vccd1 vccd1 sram_wmask0[2] sky130_fd_sc_hd__buf_2
Xoutput396 _1406_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput385 _1399_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[0] sky130_fd_sc_hd__buf_2
Xoutput363 _1380_/X vssd1 vssd1 vccd1 vccd1 sram_din0[31] sky130_fd_sc_hd__buf_2
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ _2162_/A _2085_/B _2042_/B vssd1 vssd1 vccd1 vccd1 _1957_/A sky130_fd_sc_hd__nor3_2
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1882_ _2359_/Q _2248_/A _2470_/Q _1880_/Y _1881_/X vssd1 vssd1 vccd1 vccd1 _1885_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2434_ _2434_/CLK _2434_/D vssd1 vssd1 vccd1 vccd1 _2434_/Q sky130_fd_sc_hd__dfxtp_1
X_2365_ _2459_/CLK _2365_/D vssd1 vssd1 vccd1 vccd1 _2365_/Q sky130_fd_sc_hd__dfxtp_1
X_1316_ _1311_/X _1314_/X _1315_/X _1241_/X vssd1 vssd1 vccd1 vccd1 _1316_/X sky130_fd_sc_hd__a22o_4
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2296_ _2319_/CLK _2296_/D vssd1 vssd1 vccd1 vccd1 _2296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1247_ _1231_/X _1238_/X _1241_/X _1246_/X vssd1 vssd1 vccd1 vccd1 _1247_/X sky130_fd_sc_hd__a22o_4
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1178_ _2299_/Q _2317_/Q _1180_/S vssd1 vssd1 vccd1 vccd1 _1179_/A sky130_fd_sc_hd__mux2_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _1108_/X _2138_/X _2149_/X vssd1 vssd1 vccd1 vccd1 _2422_/D sky130_fd_sc_hd__a21o_1
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2081_ _2397_/Q _2076_/Y _2080_/Y vssd1 vssd1 vccd1 vccd1 _2397_/D sky130_fd_sc_hd__o21a_1
X_1101_ _2100_/A vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__clkinv_2
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _1949_/B vssd1 vssd1 vccd1 vccd1 _2085_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1865_ _2391_/Q _1794_/A _2465_/Q _1863_/Y _1864_/X vssd1 vssd1 vccd1 vccd1 _1865_/X
+ sky130_fd_sc_hd__o221a_1
Xinput40 sram_dout0[1] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
X_1796_ _2373_/Q _2235_/A _2261_/A _1793_/Y _1795_/X vssd1 vssd1 vccd1 vccd1 _1796_/X
+ sky130_fd_sc_hd__a221o_1
Xinput51 sram_dout0[2] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 sram_dout0[3] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xinput73 sram_dout0[4] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput95 sram_dout0[6] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
Xinput84 sram_dout0[5] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2417_ _2452_/CLK _2417_/D vssd1 vssd1 vccd1 vccd1 _2417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2348_ _2414_/CLK _2348_/D vssd1 vssd1 vccd1 vccd1 _2348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2279_ _2279_/A1 _1898_/A _2277_/X vssd1 vssd1 vccd1 vccd1 _2472_/D sky130_fd_sc_hd__a21oi_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1650_ _1650_/A _1650_/B vssd1 vssd1 vccd1 vccd1 _2319_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1581_ _2301_/Q _1579_/A _1580_/Y vssd1 vssd1 vccd1 vccd1 _2301_/D sky130_fd_sc_hd__o21a_1
XFILLER_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2133_ _2046_/A _2132_/B _2132_/Y _2116_/X vssd1 vssd1 vccd1 vccd1 _2416_/D sky130_fd_sc_hd__a211o_1
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2064_ _1111_/X _2054_/X _2063_/X vssd1 vssd1 vccd1 vccd1 _2391_/D sky130_fd_sc_hd__a21o_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1917_ _2344_/Q _1912_/Y _1914_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _2344_/D sky130_fd_sc_hd__a211o_1
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1848_ _1847_/A _1847_/B _1847_/Y _1763_/A vssd1 vssd1 vccd1 vccd1 _2340_/D sky130_fd_sc_hd__a211oi_1
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1779_ _1772_/Y _2238_/A _1808_/A _2363_/Q _1778_/X vssd1 vssd1 vccd1 vccd1 _1779_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput230 sram_dout1[81] vssd1 vssd1 vccd1 vccd1 _1325_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput241 sram_dout1[91] vssd1 vssd1 vccd1 vccd1 _1296_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput252 wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 _2212_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput263 wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 _2187_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput274 wb_data_i[11] vssd1 vssd1 vccd1 vccd1 _1336_/A sky130_fd_sc_hd__clkbuf_4
Xinput285 wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _1358_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput296 wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _1379_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1702_ _1828_/C vssd1 vssd1 vccd1 vccd1 _1740_/B sky130_fd_sc_hd__inv_2
X_1633_ _2314_/Q _1631_/Y _1632_/Y vssd1 vssd1 vccd1 vccd1 _2314_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1564_ _1564_/A _1564_/B vssd1 vssd1 vccd1 vccd1 _2295_/D sky130_fd_sc_hd__nor2_1
X_1495_ input21/X _1485_/X _1490_/X input78/X vssd1 vssd1 vccd1 vccd1 _1495_/X sky130_fd_sc_hd__a22o_1
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2116_ _2116_/A vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__buf_2
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2047_ _2046_/Y _2043_/X _2030_/X vssd1 vssd1 vccd1 vccd1 _2047_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_31 _1187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_20 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1280_ _1275_/X _1278_/X _1279_/X _1241_/X vssd1 vssd1 vccd1 vccd1 _1280_/X sky130_fd_sc_hd__a22o_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1616_ _1648_/A _2309_/Q vssd1 vssd1 vccd1 vccd1 _1618_/B sky130_fd_sc_hd__and2b_1
XFILLER_160_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1547_ _2280_/Q _1547_/A1 _2187_/S vssd1 vssd1 vccd1 vccd1 _1548_/A sky130_fd_sc_hd__mux2_1
X_1478_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1478_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2450_ _2472_/CLK _2450_/D vssd1 vssd1 vccd1 vccd1 _2450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1401_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1473_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2381_ _2474_/A _2381_/D vssd1 vssd1 vccd1 vccd1 _2381_/Q sky130_fd_sc_hd__dfxtp_1
X_1332_ _1332_/A _1332_/B _1332_/C vssd1 vssd1 vccd1 vccd1 _1332_/X sky130_fd_sc_hd__or3_1
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1263_ _1263_/A0 _1263_/A1 _1263_/A2 _1263_/A3 _1251_/B _1251_/A vssd1 vssd1 vccd1
+ vccd1 _1263_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 sram_dout0[103] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1194_ _1194_/A vssd1 vssd1 vccd1 vccd1 _1195_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput320 _2284_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[0] sky130_fd_sc_hd__buf_2
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput331 _1539_/Y vssd1 vssd1 vccd1 vccd1 sram_csb0[0] sky130_fd_sc_hd__buf_2
Xoutput342 _1339_/X vssd1 vssd1 vccd1 vccd1 sram_din0[12] sky130_fd_sc_hd__buf_2
Xoutput353 _1361_/X vssd1 vssd1 vccd1 vccd1 sram_din0[22] sky130_fd_sc_hd__buf_2
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput375 _1538_/X vssd1 vssd1 vccd1 vccd1 sram_wmask0[3] sky130_fd_sc_hd__buf_2
Xoutput386 _1446_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput364 _1108_/X vssd1 vssd1 vccd1 vccd1 sram_din0[3] sky130_fd_sc_hd__buf_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput397 _1488_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _1950_/A vssd1 vssd1 vccd1 vccd1 _1950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1881_ _2357_/Q _2257_/A _2264_/A _2355_/Q vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2433_ _2435_/CLK _2433_/D vssd1 vssd1 vccd1 vccd1 _2433_/Q sky130_fd_sc_hd__dfxtp_1
X_2364_ _2459_/CLK _2364_/D vssd1 vssd1 vccd1 vccd1 _2364_/Q sky130_fd_sc_hd__dfxtp_1
X_1315_ _1315_/A0 _1315_/A1 _1315_/A2 _1315_/A3 _1251_/B _1251_/A vssd1 vssd1 vccd1
+ vccd1 _1315_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2295_ _2319_/CLK _2295_/D vssd1 vssd1 vccd1 vccd1 _2295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1246_ _1246_/A0 _1246_/A1 _1246_/A2 _1246_/A3 _1251_/B _1251_/A vssd1 vssd1 vccd1
+ vccd1 _1246_/X sky130_fd_sc_hd__mux4_1
X_1177_ _1177_/A vssd1 vssd1 vccd1 vccd1 _2291_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1100_ _1100_/A _1122_/B vssd1 vssd1 vccd1 vccd1 _2100_/A sky130_fd_sc_hd__nand2_4
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2080_ _2049_/X _2076_/Y _2079_/X vssd1 vssd1 vccd1 vccd1 _2080_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ _2351_/Q _1918_/X _1932_/Y vssd1 vssd1 vccd1 vccd1 _2351_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 sram_dout0[126] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
X_1864_ _1801_/Y _2386_/Q _1851_/Y _2466_/Q vssd1 vssd1 vccd1 vccd1 _1864_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput63 sram_dout0[40] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
Xinput52 sram_dout0[30] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput41 sram_dout0[20] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
X_1795_ _2366_/Q _2264_/A _1794_/X _2369_/Q vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput96 sram_dout0[70] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
Xinput85 sram_dout0[60] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 sram_dout0[50] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2474_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2416_ _2425_/CLK _2416_/D vssd1 vssd1 vccd1 vccd1 _2416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2347_ _2413_/CLK _2347_/D vssd1 vssd1 vccd1 vccd1 _2347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2278_ _2279_/A1 _1150_/B _2277_/X vssd1 vssd1 vccd1 vccd1 _2471_/D sky130_fd_sc_hd__o21ba_1
X_1229_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1580_ _2301_/Q _1579_/A _1714_/B vssd1 vssd1 vccd1 vccd1 _1580_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2444_/Q _2201_/A1 _2209_/S vssd1 vssd1 vccd1 vccd1 _2202_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2132_ _2132_/A _2132_/B vssd1 vssd1 vccd1 vccd1 _2132_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2063_ _2391_/Q _2058_/X _2037_/X vssd1 vssd1 vccd1 vccd1 _2063_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1916_ _2139_/A vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__buf_4
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1847_ _1847_/A _1847_/B vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1778_ _1775_/Y _2463_/Q _1777_/Y _2367_/Q vssd1 vssd1 vccd1 vccd1 _1778_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput220 sram_dout1[72] vssd1 vssd1 vccd1 vccd1 _1266_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput231 sram_dout1[82] vssd1 vssd1 vccd1 vccd1 _1210_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput242 sram_dout1[92] vssd1 vssd1 vccd1 vccd1 _1309_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput253 wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 _2214_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput286 wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__clkbuf_1
Xinput297 wb_data_i[3] vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__buf_2
Xinput264 wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 _2190_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput275 wb_data_i[12] vssd1 vssd1 vccd1 vccd1 _1338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1701_ _2418_/Q _1696_/Y _1847_/A _2132_/A _1700_/Y vssd1 vssd1 vccd1 vccd1 _1701_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1632_ _2314_/Q _1631_/Y _1650_/A vssd1 vssd1 vccd1 vccd1 _1632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1563_ _2295_/Q _1568_/D _1562_/X vssd1 vssd1 vccd1 vccd1 _1564_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1494_ input42/X _1484_/X _1477_/X _1493_/X vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__o211a_4
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2115_ _2112_/A _2409_/Q vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__and2b_1
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2046_ _2046_/A vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_10 _1111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_32 _1316_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1615_ _1615_/A vssd1 vssd1 vccd1 vccd1 _1615_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1546_ _2233_/S vssd1 vssd1 vccd1 vccd1 _2187_/S sky130_fd_sc_hd__buf_2
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1477_ _1518_/A vssd1 vssd1 vccd1 vccd1 _1477_/X sky130_fd_sc_hd__buf_2
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2029_ _2380_/Q _2022_/X _2028_/Y vssd1 vssd1 vccd1 vccd1 _2380_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1400_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1400_/X sky130_fd_sc_hd__buf_2
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2380_ _2474_/A _2380_/D vssd1 vssd1 vccd1 vccd1 _2380_/Q sky130_fd_sc_hd__dfxtp_1
X_1331_ _1233_/A _1328_/X _1330_/X _1234_/A vssd1 vssd1 vccd1 vccd1 _1332_/C sky130_fd_sc_hd__a22o_1
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1262_ _1314_/A _1262_/B vssd1 vssd1 vccd1 vccd1 _1262_/X sky130_fd_sc_hd__or2_1
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput6 sram_dout0[104] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1193_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput321 _2285_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[1] sky130_fd_sc_hd__buf_2
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput332 _1540_/Y vssd1 vssd1 vccd1 vccd1 sram_csb0[1] sky130_fd_sc_hd__buf_2
Xoutput343 _1341_/X vssd1 vssd1 vccd1 vccd1 sram_din0[13] sky130_fd_sc_hd__buf_2
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput387 _1452_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput376 _1316_/X vssd1 vssd1 vccd1 vccd1 vga_b[0] sky130_fd_sc_hd__buf_2
Xoutput365 _1111_/X vssd1 vssd1 vccd1 vccd1 sram_din0[4] sky130_fd_sc_hd__buf_2
Xoutput354 _1363_/X vssd1 vssd1 vccd1 vccd1 sram_din0[23] sky130_fd_sc_hd__buf_2
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput398 _1494_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[21] sky130_fd_sc_hd__buf_2
X_1529_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2162_/A sky130_fd_sc_hd__buf_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1880_ _2352_/Q vssd1 vssd1 vccd1 vccd1 _1880_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2432_ _2435_/CLK _2432_/D vssd1 vssd1 vccd1 vccd1 _2432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2363_ _2459_/CLK _2363_/D vssd1 vssd1 vccd1 vccd1 _2363_/Q sky130_fd_sc_hd__dfxtp_1
X_1314_ _1314_/A _1314_/B vssd1 vssd1 vccd1 vccd1 _1314_/X sky130_fd_sc_hd__or2_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2294_ _2316_/CLK _2294_/D vssd1 vssd1 vccd1 vccd1 _2294_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1245_ _1329_/A vssd1 vssd1 vccd1 vccd1 _1251_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1176_ _2298_/Q _1639_/A _1180_/S vssd1 vssd1 vccd1 vccd1 _1177_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ _2102_/A _1922_/B _1919_/X vssd1 vssd1 vccd1 vccd1 _1932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1863_ _2390_/Q vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__inv_2
Xinput31 sram_dout0[127] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
Xinput20 sram_dout0[117] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput64 sram_dout0[41] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
Xinput53 sram_dout0[31] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput42 sram_dout0[21] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
X_1794_ _1794_/A vssd1 vssd1 vccd1 vccd1 _1794_/X sky130_fd_sc_hd__clkbuf_2
Xinput97 sram_dout0[71] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput86 sram_dout0[61] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
Xinput75 sram_dout0[51] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2415_ _2446_/CLK _2415_/D vssd1 vssd1 vccd1 vccd1 _2415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2346_ _2414_/CLK _2346_/D vssd1 vssd1 vccd1 vccd1 _2346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2277_ _2472_/Q _2471_/Q _2079_/A _2185_/B vssd1 vssd1 vccd1 vccd1 _2277_/X sky130_fd_sc_hd__a211o_1
X_1228_ _1301_/A _1303_/B vssd1 vssd1 vccd1 vccd1 _1232_/A sky130_fd_sc_hd__nor2_2
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1159_ _2310_/Q vssd1 vssd1 vccd1 vccd1 _1621_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2233_/S vssd1 vssd1 vccd1 vccd1 _2209_/S sky130_fd_sc_hd__buf_2
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2131_ _2157_/A _2142_/B _2157_/C vssd1 vssd1 vccd1 vccd1 _2132_/B sky130_fd_sc_hd__nor3_2
XFILLER_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2062_ _2390_/Q _2054_/X _2061_/Y vssd1 vssd1 vccd1 vccd1 _2390_/D sky130_fd_sc_hd__o21a_1
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1915_ _1952_/A vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1846_ _1846_/A _1846_/B _1847_/B vssd1 vssd1 vccd1 vccd1 _2339_/D sky130_fd_sc_hd__nor3_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1777_ _2267_/A vssd1 vssd1 vccd1 vccd1 _1777_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2329_ _2434_/CLK _2329_/D vssd1 vssd1 vccd1 vccd1 _2329_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput210 sram_dout1[61] vssd1 vssd1 vccd1 vccd1 _1322_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput232 sram_dout1[83] vssd1 vssd1 vccd1 vccd1 _1250_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput243 sram_dout1[93] vssd1 vssd1 vccd1 vccd1 _1321_/A sky130_fd_sc_hd__clkbuf_1
Xinput221 sram_dout1[73] vssd1 vssd1 vccd1 vccd1 _1291_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput254 wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 _2216_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput265 wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 _2192_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput276 wb_data_i[13] vssd1 vssd1 vccd1 vccd1 _1340_/A sky130_fd_sc_hd__buf_2
Xinput287 wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _1362_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput298 wb_data_i[4] vssd1 vssd1 vccd1 vccd1 _1109_/A sky130_fd_sc_hd__buf_2
XFILLER_29_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1700_ _2425_/Q _1698_/Y _1699_/Y _2422_/Q vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_172_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ _1646_/B _1631_/B vssd1 vssd1 vccd1 vccd1 _1631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1562_ _1714_/B vssd1 vssd1 vccd1 vccd1 _1562_/X sky130_fd_sc_hd__buf_4
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1493_ _1493_/A1 _1489_/X _1491_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1493_/X sky130_fd_sc_hd__a211o_2
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2114_ _2408_/Q _2111_/X _2113_/Y vssd1 vssd1 vccd1 vccd1 _2408_/D sky130_fd_sc_hd__o21a_1
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2045_ _1126_/Y _2043_/X _2044_/Y _2016_/X vssd1 vssd1 vccd1 vccd1 _2385_/D sky130_fd_sc_hd__a211o_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1829_ _1824_/A _1828_/B _1828_/C vssd1 vssd1 vccd1 vccd1 _1830_/C sky130_fd_sc_hd__a21oi_1
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_33 _1334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_22 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_11 _1121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1614_ _1648_/A _1650_/A vssd1 vssd1 vccd1 vccd1 _1615_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1545_ _2222_/A vssd1 vssd1 vccd1 vccd1 _2233_/S sky130_fd_sc_hd__buf_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1476_ input38/X _1463_/X _1459_/X _1475_/X vssd1 vssd1 vccd1 vccd1 _1476_/X sky130_fd_sc_hd__o211a_4
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ _2093_/A _2019_/X _1995_/X vssd1 vssd1 vccd1 vccd1 _2028_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1330_ _1330_/A1 _1190_/A _1194_/A _1330_/B2 _1329_/X vssd1 vssd1 vccd1 vccd1 _1330_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1261_ _1261_/A1 _1233_/X _1234_/X _1261_/B2 _1260_/X vssd1 vssd1 vccd1 vccd1 _1262_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1192_ _2294_/Q _2293_/Q vssd1 vssd1 vccd1 vccd1 _1224_/A sky130_fd_sc_hd__and2b_1
Xinput7 sram_dout0[105] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput322 _2286_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[2] sky130_fd_sc_hd__buf_2
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput311 _1135_/Y vssd1 vssd1 vccd1 vccd1 sram_addr0[0] sky130_fd_sc_hd__buf_2
Xoutput333 _1541_/Y vssd1 vssd1 vccd1 vccd1 sram_csb0[2] sky130_fd_sc_hd__buf_2
Xoutput344 _1343_/X vssd1 vssd1 vccd1 vccd1 sram_din0[14] sky130_fd_sc_hd__buf_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput377 _1334_/X vssd1 vssd1 vccd1 vccd1 vga_b[1] sky130_fd_sc_hd__buf_2
Xoutput366 _1922_/A vssd1 vssd1 vccd1 vccd1 sram_din0[5] sky130_fd_sc_hd__buf_2
Xoutput355 _1365_/X vssd1 vssd1 vccd1 vccd1 sram_din0[24] sky130_fd_sc_hd__buf_2
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput388 _1455_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput399 _1497_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[22] sky130_fd_sc_hd__buf_2
X_1528_ _2280_/Q _1531_/B vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__nand2_2
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1459_ _1518_/A vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__buf_2
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2431_ _2434_/CLK _2431_/D vssd1 vssd1 vccd1 vccd1 _2431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2362_ _2425_/CLK _2362_/D vssd1 vssd1 vccd1 vccd1 _2362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1313_ _1313_/A1 _1233_/X _1234_/X _1313_/B2 _1312_/X vssd1 vssd1 vccd1 vccd1 _1314_/B
+ sky130_fd_sc_hd__a221o_1
X_2293_ _2316_/CLK _2293_/D vssd1 vssd1 vccd1 vccd1 _2293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1244_ _2294_/Q vssd1 vssd1 vccd1 vccd1 _1329_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1175_ _2316_/Q vssd1 vssd1 vccd1 vccd1 _1639_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1931_ _2350_/Q _1912_/Y _1930_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _2350_/D sky130_fd_sc_hd__a211o_1
XFILLER_147_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1862_ _2392_/Q _1800_/A _1801_/Y _2386_/Q _1861_/X vssd1 vssd1 vccd1 vccd1 _1862_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput21 sram_dout0[118] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 sram_dout0[108] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput54 sram_dout0[32] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 sram_dout0[22] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput32 sram_dout0[12] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
X_1793_ _2367_/Q vssd1 vssd1 vccd1 vccd1 _1793_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput98 sram_dout0[72] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
Xinput87 sram_dout0[62] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput76 sram_dout0[52] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_1
Xinput65 sram_dout0[42] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2414_ _2414_/CLK _2414_/D vssd1 vssd1 vccd1 vccd1 _2414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2345_ _2414_/CLK _2345_/D vssd1 vssd1 vccd1 vccd1 _2345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2276_ _2275_/A _2275_/B _2275_/Y _2239_/A vssd1 vssd1 vccd1 vccd1 _2470_/D sky130_fd_sc_hd__o211a_1
X_1227_ _1327_/A vssd1 vssd1 vccd1 vccd1 _1301_/A sky130_fd_sc_hd__clkbuf_1
X_1158_ _1158_/A vssd1 vssd1 vccd1 vccd1 _2284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _2415_/Q _2111_/X _2129_/Y vssd1 vssd1 vccd1 vccd1 _2415_/D sky130_fd_sc_hd__o21a_1
X_2061_ _1958_/X _2054_/A _2030_/X vssd1 vssd1 vccd1 vccd1 _2061_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1914_ _1914_/A _1922_/B vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__and2_1
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1845_ _1845_/A _2339_/Q _1845_/C vssd1 vssd1 vccd1 vccd1 _1847_/B sky130_fd_sc_hd__and3_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1776_ _2466_/Q vssd1 vssd1 vccd1 vccd1 _2267_/A sky130_fd_sc_hd__buf_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2337_/CLK _2328_/D vssd1 vssd1 vccd1 vccd1 _2328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2259_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput211 sram_dout1[64] vssd1 vssd1 vccd1 vccd1 _1246_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput200 sram_dout1[52] vssd1 vssd1 vccd1 vccd1 _1268_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput244 sram_dout1[96] vssd1 vssd1 vccd1 vccd1 _1246_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput233 sram_dout1[84] vssd1 vssd1 vccd1 vccd1 _1268_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput222 sram_dout1[74] vssd1 vssd1 vccd1 vccd1 _1304_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput266 wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 _2194_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput277 wb_data_i[14] vssd1 vssd1 vccd1 vccd1 _1342_/A sky130_fd_sc_hd__buf_2
Xinput255 wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 _2218_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput288 wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _1364_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput299 wb_data_i[5] vssd1 vssd1 vccd1 vccd1 _1112_/A sky130_fd_sc_hd__buf_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1630_ _1615_/X _1628_/X _1631_/B _1622_/X _1629_/A vssd1 vssd1 vccd1 vccd1 _2313_/D
+ sky130_fd_sc_hd__a32o_1
X_1561_ _2329_/Q vssd1 vssd1 vccd1 vccd1 _1714_/B sky130_fd_sc_hd__buf_2
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1492_ _1492_/A vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2113_ _1985_/X _2112_/X _2079_/X vssd1 vssd1 vccd1 vccd1 _2113_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2044_ _2044_/A _2044_/B vssd1 vssd1 vccd1 vccd1 _2044_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1828_ _1831_/A _1828_/B _1828_/C vssd1 vssd1 vccd1 vccd1 _1830_/B sky130_fd_sc_hd__and3_1
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1759_ _2433_/Q _1828_/C vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__xor2_1
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_12 _1530_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _1280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1613_ _1613_/A _2329_/Q vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__nor2_4
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1544_ _1887_/A _1898_/A _1544_/C _1544_/D vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__and4b_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1475_ input17/X _1473_/X _1447_/X _1474_/X vssd1 vssd1 vccd1 vccd1 _1475_/X sky130_fd_sc_hd__a211o_2
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2027_ _2379_/Q _2022_/X _2026_/Y vssd1 vssd1 vccd1 vccd1 _2379_/D sky130_fd_sc_hd__o21a_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ _1260_/A1 _1215_/A _1235_/X _1260_/B2 vssd1 vssd1 vccd1 vccd1 _1260_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1191_ _1191_/A vssd1 vssd1 vccd1 vccd1 _1191_/Y sky130_fd_sc_hd__inv_2
Xinput8 sram_dout0[106] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput323 _2287_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[3] sky130_fd_sc_hd__buf_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput312 _1129_/Y vssd1 vssd1 vccd1 vccd1 sram_addr0[1] sky130_fd_sc_hd__buf_2
Xoutput334 _1542_/Y vssd1 vssd1 vccd1 vccd1 sram_csb0[3] sky130_fd_sc_hd__buf_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput378 _1280_/X vssd1 vssd1 vccd1 vccd1 vga_g[0] sky130_fd_sc_hd__buf_2
Xoutput367 _1117_/X vssd1 vssd1 vccd1 vccd1 sram_din0[6] sky130_fd_sc_hd__buf_2
Xoutput345 _1346_/X vssd1 vssd1 vccd1 vccd1 sram_din0[15] sky130_fd_sc_hd__buf_2
Xoutput356 _1368_/X vssd1 vssd1 vccd1 vccd1 sram_din0[25] sky130_fd_sc_hd__buf_2
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1527_ input53/X _1442_/A _1518_/X _1526_/X vssd1 vssd1 vccd1 vccd1 _1527_/X sky130_fd_sc_hd__o211a_4
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput389 _1458_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1458_ input33/X _1442_/X _1438_/X _1457_/X vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__o211a_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1389_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1492_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2430_ _2435_/CLK _2430_/D vssd1 vssd1 vccd1 vccd1 _2430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2361_ _2425_/CLK _2361_/D vssd1 vssd1 vccd1 vccd1 _2361_/Q sky130_fd_sc_hd__dfxtp_1
X_1312_ _1312_/A1 _1215_/A _1235_/A _1312_/B2 vssd1 vssd1 vccd1 vccd1 _1312_/X sky130_fd_sc_hd__a22o_1
X_2292_ _2475_/A _2292_/D vssd1 vssd1 vccd1 vccd1 _2292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1243_ _1329_/B vssd1 vssd1 vccd1 vccd1 _1251_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1174_ _1174_/A vssd1 vssd1 vccd1 vccd1 _2290_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _1930_/A _1930_/B vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__and2_1
XFILLER_174_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1861_ _2393_/Q _1805_/A _1798_/A _2390_/Q vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput22 sram_dout0[119] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
Xinput11 sram_dout0[109] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput55 sram_dout0[33] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
Xinput44 sram_dout0[23] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
Xinput33 sram_dout0[13] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
X_1792_ _2267_/A vssd1 vssd1 vccd1 vccd1 _2261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput88 sram_dout0[63] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput77 sram_dout0[53] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput66 sram_dout0[43] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
Xinput99 sram_dout0[73] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2413_ _2413_/CLK _2413_/D vssd1 vssd1 vccd1 vccd1 _2413_/Q sky130_fd_sc_hd__dfxtp_1
X_2344_ _2414_/CLK _2344_/D vssd1 vssd1 vccd1 vccd1 _2344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2275_ _2275_/A _2275_/B vssd1 vssd1 vccd1 vccd1 _2275_/Y sky130_fd_sc_hd__nand2_1
X_1226_ _1226_/A1 _1187_/A _1225_/X vssd1 vssd1 vccd1 vccd1 _1226_/X sky130_fd_sc_hd__a21o_1
X_1157_ _2302_/Q _1621_/A _1168_/S vssd1 vssd1 vccd1 vccd1 _1158_/A sky130_fd_sc_hd__mux2_2
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2060_ _1851_/Y _2058_/X _2059_/X vssd1 vssd1 vccd1 vccd1 _2389_/D sky130_fd_sc_hd__a21oi_1
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ _1930_/B vssd1 vssd1 vccd1 vccd1 _1922_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1844_ _1845_/A _1845_/C _2339_/Q vssd1 vssd1 vccd1 vccd1 _1846_/B sky130_fd_sc_hd__a21oi_1
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1775_ _2370_/Q vssd1 vssd1 vccd1 vccd1 _1775_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2327_ _2337_/CLK _2327_/D vssd1 vssd1 vccd1 vccd1 _2327_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2258_ _2262_/A _2258_/B _2258_/C vssd1 vssd1 vccd1 vccd1 _2259_/A sky130_fd_sc_hd__and3_1
X_1209_ _1303_/A _1303_/B _1209_/C vssd1 vssd1 vccd1 vccd1 _1209_/X sky130_fd_sc_hd__and3_1
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2189_ _2233_/S vssd1 vssd1 vccd1 vccd1 _2198_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput201 sram_dout1[53] vssd1 vssd1 vccd1 vccd1 _1289_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput223 sram_dout1[75] vssd1 vssd1 vccd1 vccd1 _1328_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput212 sram_dout1[65] vssd1 vssd1 vccd1 vccd1 _1263_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput245 sram_dout1[97] vssd1 vssd1 vccd1 vccd1 _1263_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput234 sram_dout1[85] vssd1 vssd1 vccd1 vccd1 _1289_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput267 wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 _2196_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput278 wb_data_i[15] vssd1 vssd1 vccd1 vccd1 _1345_/A sky130_fd_sc_hd__clkbuf_2
Xinput256 wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 _2220_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput289 wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2459_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ _2295_/Q _1568_/D vssd1 vssd1 vccd1 vccd1 _1564_/A sky130_fd_sc_hd__and2_1
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1491_ input20/X _1485_/X _1490_/X input77/X vssd1 vssd1 vccd1 vccd1 _1491_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2112_ _2112_/A vssd1 vssd1 vccd1 vccd1 _2112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2043_ _2044_/B vssd1 vssd1 vccd1 vccd1 _2043_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1827_ _1824_/A _1828_/B _1826_/Y vssd1 vssd1 vccd1 vccd1 _2332_/D sky130_fd_sc_hd__a21oi_1
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1758_ _1758_/A _1758_/B _1757_/X vssd1 vssd1 vccd1 vccd1 _1761_/C sky130_fd_sc_hd__or3b_1
XFILLER_171_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1689_ _2409_/Q _1839_/A vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_13 _1534_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_24 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_35 _1264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1612_ _1612_/A vssd1 vssd1 vccd1 vccd1 _2308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1543_ _1909_/A vssd1 vssd1 vccd1 vccd1 _1898_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1474_ input74/X _1448_/X _1449_/X _1474_/B2 vssd1 vssd1 vccd1 vccd1 _1474_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2026_ _1958_/X _2019_/X _1995_/X vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1190_ _1190_/A vssd1 vssd1 vccd1 vccd1 _1191_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 sram_dout0[107] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput324 _2288_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[4] sky130_fd_sc_hd__buf_2
Xoutput335 _1281_/X vssd1 vssd1 vccd1 vccd1 sram_csb1[0] sky130_fd_sc_hd__buf_2
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput313 _1935_/B vssd1 vssd1 vccd1 vccd1 sram_addr0[2] sky130_fd_sc_hd__buf_2
X_1526_ _1526_/A1 _1489_/X _1525_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1526_/X sky130_fd_sc_hd__a211o_2
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput368 _1914_/A vssd1 vssd1 vccd1 vccd1 sram_din0[7] sky130_fd_sc_hd__buf_2
Xoutput346 _1348_/X vssd1 vssd1 vccd1 vccd1 sram_din0[16] sky130_fd_sc_hd__buf_2
Xoutput357 _1370_/X vssd1 vssd1 vccd1 vccd1 sram_din0[26] sky130_fd_sc_hd__buf_2
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput379 _1300_/X vssd1 vssd1 vccd1 vccd1 vga_g[1] sky130_fd_sc_hd__buf_2
X_1457_ input11/X _1443_/X _1447_/X _1456_/X vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__a211o_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1388_ _1392_/C _1386_/B _1392_/B vssd1 vssd1 vccd1 vccd1 _1478_/A sky130_fd_sc_hd__o21ai_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2009_ _2042_/A _2042_/B _2142_/B vssd1 vssd1 vccd1 vccd1 _2010_/A sky130_fd_sc_hd__nor3_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2360_ _2459_/CLK _2360_/D vssd1 vssd1 vccd1 vccd1 _2360_/Q sky130_fd_sc_hd__dfxtp_1
X_2291_ _2475_/A _2291_/D vssd1 vssd1 vccd1 vccd1 _2291_/Q sky130_fd_sc_hd__dfxtp_1
X_1311_ _1311_/A _1311_/B vssd1 vssd1 vccd1 vccd1 _1311_/X sky130_fd_sc_hd__or2_1
XFILLER_173_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1242_ _2293_/Q vssd1 vssd1 vccd1 vccd1 _1329_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1173_ _2297_/Q _2315_/Q _1180_/S vssd1 vssd1 vccd1 vccd1 _1174_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1509_ input82/X _1479_/X _1480_/X _1509_/B2 vssd1 vssd1 vccd1 vccd1 _1509_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _1857_/Y _2460_/Q _2461_/Q _1858_/Y _1859_/X vssd1 vssd1 vccd1 vccd1 _1866_/B
+ sky130_fd_sc_hd__a221o_1
Xinput12 sram_dout0[10] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1791_ _2460_/Q vssd1 vssd1 vccd1 vccd1 _2235_/A sky130_fd_sc_hd__clkinv_2
Xinput45 sram_dout0[24] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
Xinput34 sram_dout0[14] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput23 sram_dout0[11] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput89 sram_dout0[64] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
Xinput78 sram_dout0[54] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 sram_dout0[44] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
Xinput56 sram_dout0[34] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2412_ _2452_/CLK _2412_/D vssd1 vssd1 vccd1 vccd1 _2412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2343_ _2472_/CLK _2343_/D vssd1 vssd1 vccd1 vccd1 _2343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2274_ _2274_/A vssd1 vssd1 vccd1 vccd1 _2469_/D sky130_fd_sc_hd__clkbuf_1
X_1225_ _1225_/A1 _1190_/A _1224_/X _1225_/B2 vssd1 vssd1 vccd1 vccd1 _1225_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1156_ _1182_/S vssd1 vssd1 vccd1 vccd1 _1168_/S sky130_fd_sc_hd__buf_2
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2136_/A sky130_fd_sc_hd__buf_2
XFILLER_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1912_ _1930_/B vssd1 vssd1 vccd1 vccd1 _1912_/Y sky130_fd_sc_hd__inv_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1843_ _1845_/A _1845_/C _1842_/Y vssd1 vssd1 vccd1 vccd1 _2338_/D sky130_fd_sc_hd__a21oi_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1774_ _2470_/Q vssd1 vssd1 vccd1 vccd1 _1808_/A sky130_fd_sc_hd__inv_2
XFILLER_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2326_ _2337_/CLK _2326_/D vssd1 vssd1 vccd1 vccd1 _2326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ _2257_/A _2257_/B vssd1 vssd1 vccd1 vccd1 _2258_/C sky130_fd_sc_hd__nand2_1
X_1208_ _1234_/A vssd1 vssd1 vccd1 vccd1 _1208_/X sky130_fd_sc_hd__buf_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2188_ _2188_/A vssd1 vssd1 vccd1 vccd1 _2438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1139_ _1379_/B vssd1 vssd1 vccd1 vccd1 _1140_/A sky130_fd_sc_hd__buf_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput202 sram_dout1[54] vssd1 vssd1 vccd1 vccd1 _1302_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput235 sram_dout1[86] vssd1 vssd1 vccd1 vccd1 _1302_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput224 sram_dout1[76] vssd1 vssd1 vccd1 vccd1 _1225_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput213 sram_dout1[66] vssd1 vssd1 vccd1 vccd1 _1279_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput246 sram_dout1[98] vssd1 vssd1 vccd1 vccd1 _1279_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput268 wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 _2198_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput279 wb_data_i[16] vssd1 vssd1 vccd1 vccd1 _1347_/A sky130_fd_sc_hd__clkbuf_2
Xinput257 wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 _2223_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1490_ _1490_/A vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2111_ _2121_/B vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2042_ _2042_/A _2042_/B _2167_/B vssd1 vssd1 vccd1 vccd1 _2044_/B sky130_fd_sc_hd__nor3_2
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1826_ _1824_/A _1828_/B _1825_/X vssd1 vssd1 vccd1 vccd1 _1826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1757_ _2434_/Q _1683_/Y _1692_/Y _2430_/Q _1756_/Y vssd1 vssd1 vccd1 vccd1 _1757_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1688_ _2337_/Q vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_14 _1300_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2309_ _2316_/CLK _2309_/D vssd1 vssd1 vccd1 vccd1 _2309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_25 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_36 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1611_ _1609_/X _1646_/B _1611_/C vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__and3b_1
XFILLER_157_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1542_ _1342_/B _1438_/A _1407_/X vssd1 vssd1 vccd1 vccd1 _1542_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1473_ _1473_/A vssd1 vssd1 vccd1 vccd1 _1473_/X sky130_fd_sc_hd__buf_2
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2025_ _1117_/X _2022_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _2378_/D sky130_fd_sc_hd__a21o_1
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1809_ _2382_/Q _1805_/A _1777_/Y _2378_/Q vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput325 _2289_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[5] sky130_fd_sc_hd__buf_2
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput314 _1935_/A vssd1 vssd1 vccd1 vccd1 sram_addr0[3] sky130_fd_sc_hd__buf_2
Xoutput336 _1195_/Y vssd1 vssd1 vccd1 vccd1 sram_csb1[1] sky130_fd_sc_hd__buf_2
X_1525_ input31/X _1485_/A _1490_/X input88/X vssd1 vssd1 vccd1 vccd1 _1525_/X sky130_fd_sc_hd__a22o_1
Xoutput369 _1121_/Y vssd1 vssd1 vccd1 vccd1 sram_din0[8] sky130_fd_sc_hd__buf_2
Xoutput347 _1350_/X vssd1 vssd1 vccd1 vccd1 sram_din0[17] sky130_fd_sc_hd__buf_2
Xoutput358 _1372_/X vssd1 vssd1 vccd1 vccd1 sram_din0[27] sky130_fd_sc_hd__buf_2
XFILLER_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1456_ input68/X _1448_/X _1449_/X _1456_/B2 vssd1 vssd1 vccd1 vccd1 _1456_/X sky130_fd_sc_hd__a22o_1
X_1387_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2008_ _2018_/C vssd1 vssd1 vccd1 vccd1 _2142_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1310_ _1223_/X _1307_/X _1309_/X _1284_/X _1229_/X vssd1 vssd1 vccd1 vccd1 _1311_/B
+ sky130_fd_sc_hd__a221o_1
X_2290_ _2475_/A _2290_/D vssd1 vssd1 vccd1 vccd1 _2290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1241_ _1241_/A vssd1 vssd1 vccd1 vccd1 _1241_/X sky130_fd_sc_hd__buf_2
X_1172_ _1172_/A vssd1 vssd1 vccd1 vccd1 _2289_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1508_ input46/X _1505_/X _1501_/X _1507_/X vssd1 vssd1 vccd1 vccd1 _1508_/X sky130_fd_sc_hd__o211a_4
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1439_ input64/X _1409_/X _1410_/X input99/X vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 sram_dout0[110] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_2
X_1790_ _1790_/A _1790_/B _1789_/X vssd1 vssd1 vccd1 vccd1 _1790_/X sky130_fd_sc_hd__or3b_1
Xinput24 sram_dout0[120] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput46 sram_dout0[25] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
Xinput35 sram_dout0[15] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput79 sram_dout0[55] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
Xinput68 sram_dout0[45] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
Xinput57 sram_dout0[35] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2411_ _2472_/CLK _2411_/D vssd1 vssd1 vccd1 vccd1 _2411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2342_ _2472_/CLK _2342_/D vssd1 vssd1 vccd1 vccd1 _2342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2273_ _2273_/A _2273_/B _2275_/B vssd1 vssd1 vccd1 vccd1 _2274_/A sky130_fd_sc_hd__and3_1
X_1224_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1155_ _2342_/Q _2343_/Q vssd1 vssd1 vccd1 vccd1 _1182_/S sky130_fd_sc_hd__and2b_4
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1988_ _2366_/Q _1984_/X _1987_/Y vssd1 vssd1 vccd1 vccd1 _2366_/D sky130_fd_sc_hd__o21a_1
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ _2057_/A _1949_/B _1911_/C _1911_/D vssd1 vssd1 vccd1 vccd1 _1930_/B sky130_fd_sc_hd__nor4_4
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1842_ _1845_/A _1845_/C _1825_/X vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1773_ _2460_/Q vssd1 vssd1 vccd1 vccd1 _2238_/A sky130_fd_sc_hd__buf_2
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2325_ _2413_/CLK _2325_/D vssd1 vssd1 vccd1 vccd1 _2325_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ _2267_/D vssd1 vssd1 vccd1 vccd1 _2258_/B sky130_fd_sc_hd__clkinv_2
X_1207_ _1609_/A _2307_/Q _1602_/A vssd1 vssd1 vccd1 vccd1 _1234_/A sky130_fd_sc_hd__and3b_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2187_ _2438_/Q _2187_/A1 _2187_/S vssd1 vssd1 vccd1 vccd1 _2188_/A sky130_fd_sc_hd__mux2_1
X_1138_ _1366_/A vssd1 vssd1 vccd1 vccd1 _1379_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput236 sram_dout1[87] vssd1 vssd1 vccd1 vccd1 _1330_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput214 sram_dout1[67] vssd1 vssd1 vccd1 vccd1 _1283_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput225 sram_dout1[77] vssd1 vssd1 vccd1 vccd1 _1255_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput203 sram_dout1[55] vssd1 vssd1 vccd1 vccd1 _1330_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput247 sram_dout1[99] vssd1 vssd1 vccd1 vccd1 _1283_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput258 wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 _2225_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput269 wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 _2201_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2110_ _2112_/A vssd1 vssd1 vccd1 vccd1 _2121_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2041_ _2057_/C vssd1 vssd1 vccd1 vccd1 _2167_/B sky130_fd_sc_hd__buf_2
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1825_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1756_ _2431_/Q _2335_/Q vssd1 vssd1 vccd1 vccd1 _1756_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_116_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1687_ _1679_/Y _2332_/Q _1681_/X _2121_/A _1686_/X vssd1 vssd1 vccd1 vccd1 _1691_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 _1300_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2308_ _2316_/CLK _2308_/D vssd1 vssd1 vccd1 vccd1 _2308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_26 _1324_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_37 _1472_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2239_ _2239_/A _2243_/B _2239_/C vssd1 vssd1 vccd1 vccd1 _2240_/A sky130_fd_sc_hd__and3_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1610_ _1609_/B _1602_/A _1656_/B _1609_/A vssd1 vssd1 vccd1 vccd1 _1611_/C sky130_fd_sc_hd__a31o_1
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1541_ _1140_/A _1438_/A _1400_/X vssd1 vssd1 vccd1 vccd1 _1541_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1472_ input37/X _1463_/X _1459_/X _1471_/X vssd1 vssd1 vccd1 vccd1 _1472_/X sky130_fd_sc_hd__o211a_4
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2024_ _2378_/Q _2023_/X _2002_/X vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1808_ _1808_/A vssd1 vssd1 vccd1 vccd1 _2275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1739_ _1836_/A vssd1 vssd1 vccd1 vccd1 _1739_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput326 _2290_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[6] sky130_fd_sc_hd__buf_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput315 _1145_/X vssd1 vssd1 vccd1 vccd1 sram_addr0[4] sky130_fd_sc_hd__buf_2
Xoutput337 _1191_/Y vssd1 vssd1 vccd1 vccd1 sram_csb1[2] sky130_fd_sc_hd__buf_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1524_ input52/X _1442_/A _1518_/X _1523_/X vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__o211a_4
Xoutput348 _1352_/X vssd1 vssd1 vccd1 vccd1 sram_din0[18] sky130_fd_sc_hd__buf_2
Xoutput359 _1374_/X vssd1 vssd1 vccd1 vccd1 sram_din0[28] sky130_fd_sc_hd__buf_2
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1455_ input32/X _1442_/X _1438_/X _1454_/X vssd1 vssd1 vccd1 vccd1 _1455_/X sky130_fd_sc_hd__o211a_4
X_1386_ _1392_/C _1386_/B _1392_/B vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__and3_4
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2007_ _2040_/C _2438_/Q _1129_/Y vssd1 vssd1 vccd1 vccd1 _2018_/C sky130_fd_sc_hd__or3b_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1240_ _1240_/A _1240_/B vssd1 vssd1 vccd1 vccd1 _1241_/A sky130_fd_sc_hd__nor2_1
X_1171_ _2296_/Q _2314_/Q _1180_/S vssd1 vssd1 vccd1 vccd1 _1172_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1507_ input25/X _1473_/X _1478_/X _1506_/X vssd1 vssd1 vccd1 vccd1 _1507_/X sky130_fd_sc_hd__a211o_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1438_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__buf_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1369_ _1369_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1370_/A sky130_fd_sc_hd__and2_1
XFILLER_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput25 sram_dout0[121] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 sram_dout0[111] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput36 sram_dout0[16] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput69 sram_dout0[46] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
Xinput58 sram_dout0[36] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
Xinput47 sram_dout0[26] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2410_ _2446_/CLK _2410_/D vssd1 vssd1 vccd1 vccd1 _2410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2341_ _2468_/CLK _2341_/D vssd1 vssd1 vccd1 vccd1 _2341_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2272_ _2272_/A _2272_/B vssd1 vssd1 vccd1 vccd1 _2275_/B sky130_fd_sc_hd__nand2_1
X_1223_ _1235_/A vssd1 vssd1 vccd1 vccd1 _1223_/X sky130_fd_sc_hd__buf_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1154_ _2309_/Q vssd1 vssd1 vccd1 vccd1 _1621_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1987_ _1985_/X _1986_/X _1940_/X vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _2074_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _1911_/D sky130_fd_sc_hd__or2_1
X_1841_ _1845_/C _1841_/B vssd1 vssd1 vccd1 vccd1 _2337_/D sky130_fd_sc_hd__nor2_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1772_ _2373_/Q vssd1 vssd1 vccd1 vccd1 _1772_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2324_ _2425_/CLK _2324_/D vssd1 vssd1 vccd1 vccd1 _2324_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _2464_/Q _2465_/Q _2255_/C vssd1 vssd1 vccd1 vccd1 _2267_/D sky130_fd_sc_hd__and3_2
X_1206_ _1206_/A1 _1201_/X _1202_/X _1206_/B2 _1205_/X vssd1 vssd1 vccd1 vccd1 _1206_/X
+ sky130_fd_sc_hd__a221o_1
X_2186_ _2437_/Q _1898_/A _2185_/Y vssd1 vssd1 vccd1 vccd1 _2437_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1137_ _2074_/B vssd1 vssd1 vccd1 vccd1 _1935_/B sky130_fd_sc_hd__clkinv_2
XFILLER_26_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput226 sram_dout1[78] vssd1 vssd1 vccd1 vccd1 _1270_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput215 sram_dout1[68] vssd1 vssd1 vccd1 vccd1 _1315_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput204 sram_dout1[56] vssd1 vssd1 vccd1 vccd1 _1221_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput237 sram_dout1[88] vssd1 vssd1 vccd1 vccd1 _1221_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput248 sram_dout1[9] vssd1 vssd1 vccd1 vccd1 _1286_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput259 wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 _2227_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2040_ _2040_/A _2040_/B _2040_/C vssd1 vssd1 vccd1 vccd1 _2057_/C sky130_fd_sc_hd__or3_1
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1824_ _1824_/A _1846_/A vssd1 vssd1 vccd1 vccd1 _2331_/D sky130_fd_sc_hd__nor2_1
XFILLER_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1755_ _2430_/Q _1692_/Y _2340_/Q _2158_/A vssd1 vssd1 vccd1 vccd1 _1758_/B sky130_fd_sc_hd__a22o_1
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1686_ _2414_/Q _1683_/Y _1847_/A _2105_/A vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2316_/CLK _2307_/D vssd1 vssd1 vccd1 vccd1 _2307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_16 _1300_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_27 _1295_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_38 _1538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _2238_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2239_/C sky130_fd_sc_hd__or2_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2169_ _2429_/Q _2171_/B _1889_/X vssd1 vssd1 vccd1 vccd1 _2169_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _1140_/A _1518_/X _1402_/X vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_153_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1471_ _1471_/A1 _1432_/X _1470_/X _1435_/X vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__a211o_2
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2023_ _2136_/A _2052_/B _2142_/B vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__or3_2
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1807_ _2384_/Q vssd1 vssd1 vccd1 vccd1 _1807_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2425_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1738_ _1736_/Y _1831_/A _1692_/Y _2400_/Q _1737_/X vssd1 vssd1 vccd1 vccd1 _1738_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1669_ _2412_/Q _2334_/Q vssd1 vssd1 vccd1 vccd1 _1669_/X sky130_fd_sc_hd__xor2_1
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput316 _1147_/X vssd1 vssd1 vccd1 vccd1 sram_addr0[5] sky130_fd_sc_hd__buf_2
Xoutput327 _2291_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[7] sky130_fd_sc_hd__buf_2
Xoutput338 _1187_/Y vssd1 vssd1 vccd1 vccd1 sram_csb1[3] sky130_fd_sc_hd__buf_2
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1523_ input30/X _1443_/A _1492_/A _1522_/X vssd1 vssd1 vccd1 vccd1 _1523_/X sky130_fd_sc_hd__a211o_2
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput349 _1354_/X vssd1 vssd1 vccd1 vccd1 sram_din0[19] sky130_fd_sc_hd__buf_2
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1454_ _1454_/A1 _1432_/X _1453_/X _1435_/X vssd1 vssd1 vccd1 vccd1 _1454_/X sky130_fd_sc_hd__a211o_2
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1385_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1385_/X sky130_fd_sc_hd__buf_2
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2006_ _1098_/X _1986_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _2373_/D sky130_fd_sc_hd__a21o_1
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1170_ _1182_/S vssd1 vssd1 vccd1 vccd1 _1180_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1506_ input81/X _1479_/X _1480_/X _1506_/B2 vssd1 vssd1 vccd1 vccd1 _1506_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1437_ _1437_/A1 _1421_/X _1417_/X _1436_/X vssd1 vssd1 vccd1 vccd1 _1437_/X sky130_fd_sc_hd__o211a_4
X_1368_ _1368_/A vssd1 vssd1 vccd1 vccd1 _1368_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1299_ _1281_/X _1286_/X _1298_/X vssd1 vssd1 vccd1 vccd1 _1299_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 sram_dout0[122] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput15 sram_dout0[112] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
Xinput37 sram_dout0[17] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput59 sram_dout0[37] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
Xinput48 sram_dout0[27] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2340_ _2434_/CLK _2340_/D vssd1 vssd1 vccd1 vccd1 _2340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2271_ _2272_/A _2272_/B vssd1 vssd1 vccd1 vccd1 _2273_/B sky130_fd_sc_hd__or2_1
X_1222_ _2308_/Q _2306_/Q _2307_/Q vssd1 vssd1 vccd1 vccd1 _1235_/A sky130_fd_sc_hd__nor3b_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1153_ _1153_/A vssd1 vssd1 vccd1 vccd1 _1153_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1986_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__buf_2
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2469_ _2474_/A _2469_/D vssd1 vssd1 vccd1 vccd1 _2469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _1839_/A _1839_/B _1825_/X vssd1 vssd1 vccd1 vccd1 _1841_/B sky130_fd_sc_hd__o21ai_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1771_ _1768_/Y _2465_/Q _2267_/C _1770_/Y vssd1 vssd1 vccd1 vccd1 _1790_/B sky130_fd_sc_hd__a22o_1
XFILLER_155_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2413_/CLK _2323_/D vssd1 vssd1 vccd1 vccd1 _2323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2464_/D sky130_fd_sc_hd__clkbuf_1
X_1205_ _1303_/A _1303_/B _1205_/C vssd1 vssd1 vccd1 vccd1 _1205_/X sky130_fd_sc_hd__and3_1
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2185_ _2185_/A _2185_/B vssd1 vssd1 vccd1 vccd1 _2185_/Y sky130_fd_sc_hd__nor2_1
X_1136_ _2440_/Q _1136_/B vssd1 vssd1 vccd1 vccd1 _2074_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1969_ _2361_/Q _1950_/A _1966_/X vssd1 vssd1 vccd1 vccd1 _1969_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput216 sram_dout1[69] vssd1 vssd1 vccd1 vccd1 _1317_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput227 sram_dout1[79] vssd1 vssd1 vccd1 vccd1 _1294_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput205 sram_dout1[57] vssd1 vssd1 vccd1 vccd1 _1257_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput238 sram_dout1[89] vssd1 vssd1 vccd1 vccd1 _1257_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput249 wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 _2205_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1823_ _1766_/X _1790_/X _1796_/X _1822_/X vssd1 vssd1 vccd1 vccd1 _2330_/D sky130_fd_sc_hd__o31a_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1754_ _2426_/Q vssd1 vssd1 vccd1 vccd1 _2158_/A sky130_fd_sc_hd__inv_2
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1685_ _2406_/Q vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__inv_2
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2316_/CLK _2306_/D vssd1 vssd1 vccd1 vccd1 _2306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_17 _1300_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_28 _1336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _2238_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2243_/B sky130_fd_sc_hd__nand2_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _2168_/A vssd1 vssd1 vccd1 vccd1 _2171_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1119_ _1985_/A vssd1 vssd1 vccd1 vccd1 _1914_/A sky130_fd_sc_hd__inv_4
X_2099_ _2403_/Q _2084_/X _2098_/Y _2094_/X vssd1 vssd1 vccd1 vccd1 _2403_/D sky130_fd_sc_hd__a211o_1
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ input16/X _1425_/X _1433_/X input72/X vssd1 vssd1 vccd1 vccd1 _1470_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2022_ _2022_/A vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1806_ _2382_/Q _2243_/A _1794_/X _2380_/Q vssd1 vssd1 vccd1 vccd1 _1806_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1737_ _2396_/Q _1847_/A vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__xor2_1
XFILLER_171_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1668_ _2415_/Q _1824_/A vssd1 vssd1 vccd1 vccd1 _1668_/X sky130_fd_sc_hd__xor2_1
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1599_ _2341_/Q vssd1 vssd1 vccd1 vccd1 _1656_/A sky130_fd_sc_hd__inv_6
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput317 _1149_/X vssd1 vssd1 vccd1 vccd1 sram_addr0[6] sky130_fd_sc_hd__buf_2
Xoutput328 _2292_/Q vssd1 vssd1 vccd1 vccd1 sram_addr1[8] sky130_fd_sc_hd__buf_2
X_1522_ input87/X _1490_/A _1489_/A _1522_/B2 vssd1 vssd1 vccd1 vccd1 _1522_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput339 _1098_/X vssd1 vssd1 vccd1 vccd1 sram_din0[0] sky130_fd_sc_hd__buf_2
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1453_ input10/X _1425_/X _1433_/X input67/X vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__a22o_1
X_1384_ _1505_/A vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__buf_2
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2005_ _2373_/Q _1990_/X _2002_/X vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1505_ _1505_/A vssd1 vssd1 vccd1 vccd1 _1505_/X sky130_fd_sc_hd__buf_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1436_ input98/X _1432_/X _1434_/X _1435_/X vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__a211o_2
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1367_ _1367_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__and2_1
XFILLER_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1298_ _1298_/A _1298_/B vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__or2_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 sram_dout0[123] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput16 sram_dout0[113] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput49 sram_dout0[28] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
Xinput38 sram_dout0[18] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2270_ _2270_/A vssd1 vssd1 vccd1 vccd1 _2468_/D sky130_fd_sc_hd__clkbuf_1
X_1221_ _1221_/A1 _1216_/X _1217_/X _1221_/B2 _1220_/X vssd1 vssd1 vccd1 vccd1 _1221_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1152_ _2446_/Q _1537_/B vssd1 vssd1 vccd1 vccd1 _1153_/A sky130_fd_sc_hd__and2_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _1985_/A vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2468_ _2468_/CLK _2468_/D vssd1 vssd1 vccd1 vccd1 _2468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1419_ input93/X _1400_/X _1418_/X _1404_/X vssd1 vssd1 vccd1 vccd1 _1419_/X sky130_fd_sc_hd__a211o_1
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2399_ _2414_/CLK _2399_/D vssd1 vssd1 vccd1 vccd1 _2399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ _2365_/Q vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2322_ _2413_/CLK _2322_/D vssd1 vssd1 vccd1 vccd1 _2322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _2262_/A _2257_/B _2253_/C vssd1 vssd1 vccd1 vccd1 _2254_/A sky130_fd_sc_hd__and3_1
X_1204_ _1327_/B vssd1 vssd1 vccd1 vccd1 _1303_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2184_ _1544_/C _1544_/D _1537_/B vssd1 vssd1 vccd1 vccd1 _2185_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1135_ _2040_/B vssd1 vssd1 vccd1 vccd1 _1135_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1968_ _1105_/X _1957_/X _1967_/X vssd1 vssd1 vccd1 vccd1 _2360_/D sky130_fd_sc_hd__a21o_1
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1899_ _1899_/A _1949_/B _1911_/C _1899_/D vssd1 vssd1 vccd1 vccd1 _1904_/S sky130_fd_sc_hd__or4_2
XFILLER_174_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput206 sram_dout1[58] vssd1 vssd1 vccd1 vccd1 _1273_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput217 sram_dout1[6] vssd1 vssd1 vccd1 vccd1 _1237_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput239 sram_dout1[8] vssd1 vssd1 vccd1 vccd1 _1277_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput228 sram_dout1[7] vssd1 vssd1 vccd1 vccd1 _1261_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1822_ _1803_/X _1818_/X _1821_/Y _2330_/Q vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__a31o_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1753_ _2435_/Q _2331_/Q vssd1 vssd1 vccd1 vccd1 _1758_/A sky130_fd_sc_hd__xor2_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1684_ _2340_/Q vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__buf_2
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2316_/CLK _2305_/D vssd1 vssd1 vccd1 vccd1 _2305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_18 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_29 _1338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2236_/A vssd1 vssd1 vccd1 vccd1 _2460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2167_ _2167_/A _2167_/B _2167_/C vssd1 vssd1 vccd1 vccd1 _2168_/A sky130_fd_sc_hd__or3_2
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1118_ _1118_/A _1118_/B vssd1 vssd1 vccd1 vccd1 _1985_/A sky130_fd_sc_hd__nand2_4
XFILLER_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2098_ _2098_/A _2100_/B vssd1 vssd1 vccd1 vccd1 _2098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2021_ _1914_/A _2019_/X _2020_/Y _2016_/X vssd1 vssd1 vccd1 vccd1 _2377_/D sky130_fd_sc_hd__a211o_1
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1805_ _1805_/A vssd1 vssd1 vccd1 vccd1 _2243_/A sky130_fd_sc_hd__clkbuf_2
X_1736_ _2405_/Q vssd1 vssd1 vccd1 vccd1 _1736_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1667_ _1831_/A vssd1 vssd1 vccd1 vccd1 _1824_/A sky130_fd_sc_hd__buf_2
X_1598_ _1598_/A _1598_/B vssd1 vssd1 vccd1 vccd1 _2304_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2219_ _2219_/A vssd1 vssd1 vccd1 vccd1 _2452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1521_ input50/X _1505_/X _1518_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _1521_/X sky130_fd_sc_hd__o211a_4
Xoutput329 _2474_/X vssd1 vssd1 vccd1 vccd1 sram_clk0 sky130_fd_sc_hd__clkbuf_1
Xoutput318 _1151_/X vssd1 vssd1 vccd1 vccd1 sram_addr0[7] sky130_fd_sc_hd__buf_2
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1452_ input23/X _1442_/X _1438_/X _1451_/X vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__o211a_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1383_ _1392_/C _1386_/B _1392_/B vssd1 vssd1 vccd1 vccd1 _1505_/A sky130_fd_sc_hd__o21a_1
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2004_ _1102_/X _1986_/X _2003_/X vssd1 vssd1 vccd1 vccd1 _2372_/D sky130_fd_sc_hd__a21o_1
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1719_ _1719_/A _2326_/Q _2327_/Q vssd1 vssd1 vccd1 vccd1 _1725_/B sky130_fd_sc_hd__nand3_1
XFILLER_172_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1504_ input45/X _1484_/X _1501_/X _1503_/X vssd1 vssd1 vccd1 vccd1 _1504_/X sky130_fd_sc_hd__o211a_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1435_ _1492_/A vssd1 vssd1 vccd1 vccd1 _1435_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1366_ _1366_/A vssd1 vssd1 vccd1 vccd1 _1375_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1297_ _1235_/X _1294_/X _1296_/X _1284_/X _1232_/A vssd1 vssd1 vccd1 vccd1 _1298_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput28 sram_dout0[124] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 sram_dout0[114] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 sram_dout0[19] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1220_ _1308_/A _1308_/B _1220_/C vssd1 vssd1 vccd1 vccd1 _1220_/X sky130_fd_sc_hd__and3_1
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1151_ _1151_/A vssd1 vssd1 vccd1 vccd1 _1151_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__buf_2
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2467_ _2468_/CLK _2467_/D vssd1 vssd1 vccd1 vccd1 _2467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1418_ input2/X _1473_/A _1402_/X input58/X vssd1 vssd1 vccd1 vccd1 _1418_/X sky130_fd_sc_hd__a22o_1
X_2398_ _2414_/CLK _2398_/D vssd1 vssd1 vccd1 vccd1 _2398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1349_ _1349_/A _1353_/B vssd1 vssd1 vccd1 vccd1 _1350_/A sky130_fd_sc_hd__and2_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2321_ _2413_/CLK _2321_/D vssd1 vssd1 vccd1 vccd1 _2321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2464_/Q _2255_/C vssd1 vssd1 vccd1 vccd1 _2253_/C sky130_fd_sc_hd__or2_1
X_1203_ _1327_/A vssd1 vssd1 vccd1 vccd1 _1303_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ _1140_/A _1398_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _2436_/D sky130_fd_sc_hd__o21ba_4
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1134_ _2438_/Q _1531_/B vssd1 vssd1 vccd1 vccd1 _2040_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1967_ _2360_/Q _1950_/X _1966_/X vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1898_ _1898_/A _1909_/B _1898_/C vssd1 vssd1 vccd1 vccd1 _1899_/D sky130_fd_sc_hd__or3_1
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput207 sram_dout1[59] vssd1 vssd1 vccd1 vccd1 _1296_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput218 sram_dout1[70] vssd1 vssd1 vccd1 vccd1 _1206_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput229 sram_dout1[80] vssd1 vssd1 vccd1 vccd1 _1307_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1821_ _2381_/Q _2248_/A _2257_/A _2379_/Q _1820_/X vssd1 vssd1 vccd1 vccd1 _1821_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1752_ _1747_/X _1748_/Y _1749_/Y _1750_/X _1751_/X vssd1 vssd1 vccd1 vccd1 _1761_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1683_ _2332_/Q vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2316_/CLK _2304_/D vssd1 vssd1 vccd1 vccd1 _2304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_19 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2235_ _2235_/A _2239_/A vssd1 vssd1 vccd1 vccd1 _2236_/A sky130_fd_sc_hd__and2_1
X_2166_ _2428_/Q _2163_/X _2165_/Y vssd1 vssd1 vccd1 vccd1 _2428_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1117_ _1117_/A vssd1 vssd1 vccd1 vccd1 _1117_/X sky130_fd_sc_hd__buf_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2097_ _2402_/Q _2085_/Y _2096_/Y vssd1 vssd1 vccd1 vccd1 _2402_/D sky130_fd_sc_hd__o21a_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2020_ _2020_/A _2022_/A vssd1 vssd1 vccd1 vccd1 _2020_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1804_ _2462_/Q vssd1 vssd1 vccd1 vccd1 _1805_/A sky130_fd_sc_hd__clkinv_2
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1735_ _2401_/Q vssd1 vssd1 vccd1 vccd1 _1735_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1666_ _2331_/Q vssd1 vssd1 vccd1 vccd1 _1831_/A sky130_fd_sc_hd__clkbuf_2
X_1597_ _2304_/Q _1595_/A _1613_/A vssd1 vssd1 vccd1 vccd1 _1598_/B sky130_fd_sc_hd__o21ai_1
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2218_ _2452_/Q _2218_/A1 _2220_/S vssd1 vssd1 vccd1 vccd1 _2219_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2149_ _2422_/Q _2142_/X _2071_/X vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1520_ input29/X _1443_/A _1492_/A _1519_/X vssd1 vssd1 vccd1 vccd1 _1520_/X sky130_fd_sc_hd__a211o_2
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput319 _1153_/X vssd1 vssd1 vccd1 vccd1 sram_addr0[8] sky130_fd_sc_hd__buf_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1451_ input9/X _1443_/X _1447_/X _1450_/X vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__a211o_2
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1382_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _1386_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _2372_/Q _1990_/X _2002_/X vssd1 vssd1 vccd1 vccd1 _2003_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1718_ _1719_/A _2326_/Q _1717_/Y vssd1 vssd1 vccd1 vccd1 _2326_/D sky130_fd_sc_hd__a21oi_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1649_ _2319_/Q _1649_/B vssd1 vssd1 vccd1 vccd1 _1650_/B sky130_fd_sc_hd__xor2_1
XFILLER_144_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2452_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1503_ _1503_/A1 _1489_/X _1502_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1503_/X sky130_fd_sc_hd__a211o_2
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1434_ input6/X _1425_/X _1433_/X input63/X vssd1 vssd1 vccd1 vccd1 _1434_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1365_ _1365_/A vssd1 vssd1 vccd1 vccd1 _1365_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1296_ _1296_/A1 _1321_/B _1194_/A _1296_/B2 _1295_/X vssd1 vssd1 vccd1 vccd1 _1296_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput18 sram_dout0[115] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput29 sram_dout0[125] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ _2445_/Q _1150_/B vssd1 vssd1 vccd1 vccd1 _1151_/A sky130_fd_sc_hd__and2_2
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ _2167_/A _2052_/B _2109_/B vssd1 vssd1 vccd1 vccd1 _1986_/A sky130_fd_sc_hd__nor3_2
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2466_ _2468_/CLK _2466_/D vssd1 vssd1 vccd1 vccd1 _2466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1417_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1417_/X sky130_fd_sc_hd__buf_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2397_ _2452_/CLK _2397_/D vssd1 vssd1 vccd1 vccd1 _2397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1348_ _1348_/A vssd1 vssd1 vccd1 vccd1 _1348_/X sky130_fd_sc_hd__clkbuf_1
X_1279_ _1279_/A0 _1279_/A1 _1279_/A2 _1279_/A3 _1251_/B _1251_/A vssd1 vssd1 vccd1
+ vccd1 _1279_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2320_ _2413_/CLK _2320_/D vssd1 vssd1 vccd1 vccd1 _2320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _2464_/Q _2255_/C vssd1 vssd1 vccd1 vccd1 _2257_/B sky130_fd_sc_hd__nand2_1
X_1202_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1202_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2182_ _1098_/A _2164_/X _2181_/X vssd1 vssd1 vccd1 vccd1 _2435_/D sky130_fd_sc_hd__a21o_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1133_ _1136_/B vssd1 vssd1 vccd1 vccd1 _1531_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1966_ _2071_/A vssd1 vssd1 vccd1 vccd1 _1966_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1897_ _1909_/C _1907_/C _1897_/C vssd1 vssd1 vccd1 vccd1 _1898_/C sky130_fd_sc_hd__or3_1
XFILLER_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput208 sram_dout1[5] vssd1 vssd1 vccd1 vccd1 _1317_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput219 sram_dout1[71] vssd1 vssd1 vccd1 vccd1 _1252_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2449_ _2472_/CLK _2449_/D vssd1 vssd1 vccd1 vccd1 _2449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ _2383_/Q _1815_/Y _2267_/B _2020_/A _1819_/X vssd1 vssd1 vccd1 vccd1 _1820_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1751_ _2427_/Q _2339_/Q vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__xor2_1
XFILLER_144_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1682_ _2411_/Q vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__inv_2
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2316_/CLK _2303_/D vssd1 vssd1 vccd1 vccd1 _2303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2234_/A vssd1 vssd1 vccd1 vccd1 _2459_/D sky130_fd_sc_hd__clkbuf_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _1985_/X _2164_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1116_ _2089_/A vssd1 vssd1 vccd1 vccd1 _1117_/A sky130_fd_sc_hd__inv_2
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2096_ _1107_/A _2085_/Y _2079_/X vssd1 vssd1 vccd1 vccd1 _2096_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2434_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1949_ _2167_/A _1949_/B _2057_/B vssd1 vssd1 vccd1 vccd1 _1950_/A sky130_fd_sc_hd__or3_2
XFILLER_147_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1803_ _2380_/Q _1794_/X _2257_/A _2379_/Q _1802_/X vssd1 vssd1 vccd1 vccd1 _1803_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1734_ _2403_/Q _1740_/B _1733_/X vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__a21bo_1
XFILLER_156_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1665_ _1665_/A vssd1 vssd1 vccd1 vccd1 _2323_/D sky130_fd_sc_hd__clkbuf_1
X_1596_ _2304_/Q _2303_/Q _1596_/C vssd1 vssd1 vccd1 vccd1 _1598_/A sky130_fd_sc_hd__and3_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2217_ _2217_/A vssd1 vssd1 vccd1 vccd1 _2451_/D sky130_fd_sc_hd__clkbuf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2148_ _1111_/X _2137_/X _2147_/X vssd1 vssd1 vccd1 vccd1 _2421_/D sky130_fd_sc_hd__a21o_1
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ _2079_/A vssd1 vssd1 vccd1 vccd1 _2079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1450_ input66/X _1448_/X _1449_/X _1450_/B2 vssd1 vssd1 vccd1 vccd1 _1450_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1381_ _2448_/Q vssd1 vssd1 vccd1 vccd1 _1392_/C sky130_fd_sc_hd__buf_6
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2002_ _2071_/A vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1717_ _1719_/A _2326_/Q _1726_/A vssd1 vssd1 vccd1 vccd1 _1717_/Y sky130_fd_sc_hd__o21ai_1
X_1648_ _1648_/A _1648_/B _2318_/Q vssd1 vssd1 vccd1 vccd1 _1649_/B sky130_fd_sc_hd__or3b_1
XFILLER_144_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1579_ _1579_/A _1579_/B vssd1 vssd1 vccd1 vccd1 _2300_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1502_ input24/X _1485_/X _1490_/X input80/X vssd1 vssd1 vccd1 vccd1 _1502_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433_ _1490_/A vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1364_ _1364_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1365_/A sky130_fd_sc_hd__and2_1
X_1295_ _1329_/A _1329_/B _1295_/C vssd1 vssd1 vccd1 vccd1 _1295_/X sky130_fd_sc_hd__and3_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 sram_dout0[116] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ _1121_/Y _1976_/X _1981_/X _1944_/X vssd1 vssd1 vccd1 vccd1 _2365_/D sky130_fd_sc_hd__a211o_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2465_ _2468_/CLK _2465_/D vssd1 vssd1 vccd1 vccd1 _2465_/Q sky130_fd_sc_hd__dfxtp_2
X_2396_ _2452_/CLK _2396_/D vssd1 vssd1 vccd1 vccd1 _2396_/Q sky130_fd_sc_hd__dfxtp_1
X_1416_ input62/X _1385_/X _1398_/X _1415_/X vssd1 vssd1 vccd1 vccd1 _1416_/X sky130_fd_sc_hd__o211a_4
X_1347_ _1347_/A _1353_/B vssd1 vssd1 vccd1 vccd1 _1348_/A sky130_fd_sc_hd__and2_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1278_ _1314_/A _1278_/B vssd1 vssd1 vccd1 vccd1 _1278_/X sky130_fd_sc_hd__or2_1
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2250_/A vssd1 vssd1 vccd1 vccd1 _2463_/D sky130_fd_sc_hd__clkbuf_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ _1287_/A vssd1 vssd1 vccd1 vccd1 _1201_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2181_ _2435_/Q _2168_/A _1889_/X vssd1 vssd1 vccd1 vccd1 _2181_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1132_ _1132_/A vssd1 vssd1 vccd1 vccd1 _1935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1965_ _1108_/X _1957_/X _1964_/X vssd1 vssd1 vccd1 vccd1 _2359_/D sky130_fd_sc_hd__a21o_1
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1896_ _2448_/Q _2449_/Q _2450_/Q _2451_/Q vssd1 vssd1 vccd1 vccd1 _1897_/C sky130_fd_sc_hd__or4_1
XFILLER_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput209 sram_dout1[60] vssd1 vssd1 vccd1 vccd1 _1309_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2448_ _2472_/CLK _2448_/D vssd1 vssd1 vccd1 vccd1 _2448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2379_ _2474_/A _2379_/D vssd1 vssd1 vccd1 vccd1 _2379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _2428_/Q _2338_/Q vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__or2_1
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1681_ _1836_/A vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2302_ _2316_/CLK _2302_/D vssd1 vssd1 vccd1 vccd1 _2302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2233_ _2459_/Q _2233_/A1 _2233_/S vssd1 vssd1 vccd1 vccd1 _2234_/A sky130_fd_sc_hd__mux2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2164_ _2164_/A vssd1 vssd1 vccd1 vccd1 _2164_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1115_ _1115_/A _1366_/A vssd1 vssd1 vccd1 vccd1 _2089_/A sky130_fd_sc_hd__nand2_8
X_2095_ _2401_/Q _2084_/X _2093_/Y _2094_/X vssd1 vssd1 vccd1 vccd1 _2401_/D sky130_fd_sc_hd__a211o_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1948_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2167_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1879_ _2357_/Q _2257_/A _2267_/B _1877_/Y _1878_/X vssd1 vssd1 vccd1 vccd1 _1885_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1802_ _2381_/Q _2248_/A _1801_/Y _2375_/Q vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1733_ _2402_/Q _1699_/Y _1671_/X _2397_/Q vssd1 vssd1 vccd1 vccd1 _1733_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1664_ _1664_/A _1664_/B _1664_/C vssd1 vssd1 vccd1 vccd1 _1665_/A sky130_fd_sc_hd__and3_1
X_1595_ _1595_/A _1595_/B vssd1 vssd1 vccd1 vccd1 _2303_/D sky130_fd_sc_hd__nor2_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2216_ _2451_/Q _2216_/A1 _2220_/S vssd1 vssd1 vccd1 vccd1 _2217_/A sky130_fd_sc_hd__mux2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2147_ _2421_/Q _2142_/X _2071_/X vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _1124_/X _2076_/Y _2077_/X _2016_/X vssd1 vssd1 vccd1 vccd1 _2396_/D sky130_fd_sc_hd__a211o_1
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1380_ _1380_/A vssd1 vssd1 vccd1 vccd1 _1380_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2001_ _1105_/X _1986_/X _2000_/X vssd1 vssd1 vccd1 vccd1 _2371_/D sky130_fd_sc_hd__a21o_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1716_ _1716_/A vssd1 vssd1 vccd1 vccd1 _2325_/D sky130_fd_sc_hd__clkbuf_1
X_1647_ _2318_/Q _1644_/A _1646_/X vssd1 vssd1 vccd1 vccd1 _2318_/D sky130_fd_sc_hd__a21bo_1
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1578_ _2300_/Q _1576_/A _1714_/B vssd1 vssd1 vccd1 vccd1 _1579_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1501_ _1518_/A vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__buf_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1432_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1432_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1363_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1363_/X sky130_fd_sc_hd__clkbuf_1
X_1294_ _1294_/A1 _1190_/A _1194_/A _1294_/B2 _1293_/X vssd1 vssd1 vccd1 vccd1 _1294_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ _1976_/A _2365_/Q vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _2468_/CLK _2464_/D vssd1 vssd1 vccd1 vccd1 _2464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1415_ _1415_/A1 _1407_/X _1408_/X _1414_/X vssd1 vssd1 vccd1 vccd1 _1415_/X sky130_fd_sc_hd__a211o_2
X_2395_ _2435_/CLK _2395_/D vssd1 vssd1 vccd1 vccd1 _2395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1346_ _1346_/A vssd1 vssd1 vccd1 vccd1 _1346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1277_ _1277_/A1 _1233_/X _1234_/X _1277_/B2 _1276_/X vssd1 vssd1 vccd1 vccd1 _1278_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1200_/X sky130_fd_sc_hd__buf_2
X_2180_ _1930_/A _2164_/X _2179_/X vssd1 vssd1 vccd1 vccd1 _2434_/D sky130_fd_sc_hd__a21o_1
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ _2441_/Q _1136_/B vssd1 vssd1 vccd1 vccd1 _1132_/A sky130_fd_sc_hd__and2_1
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1964_ _2359_/Q _1950_/X _2185_/A vssd1 vssd1 vccd1 vccd1 _1964_/X sky130_fd_sc_hd__a21o_1
XFILLER_159_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1895_ _2453_/Q _2454_/Q _2455_/Q _2452_/Q vssd1 vssd1 vccd1 vccd1 _1907_/C sky130_fd_sc_hd__or4b_1
XFILLER_174_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2447_ _2472_/CLK _2447_/D vssd1 vssd1 vccd1 vccd1 _2447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2378_ _2474_/A _2378_/D vssd1 vssd1 vccd1 vccd1 _2378_/Q sky130_fd_sc_hd__dfxtp_1
X_1329_ _1329_/A _1329_/B _1329_/C vssd1 vssd1 vccd1 vccd1 _1329_/X sky130_fd_sc_hd__and3_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _2335_/Q vssd1 vssd1 vccd1 vccd1 _1836_/A sky130_fd_sc_hd__buf_2
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2301_ _2319_/CLK _2301_/D vssd1 vssd1 vccd1 vccd1 _2301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2232_ _2232_/A vssd1 vssd1 vccd1 vccd1 _2458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2163_ _2164_/A vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1114_ _1122_/B vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2094_ _2116_/A vssd1 vssd1 vccd1 vccd1 _2094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1947_ _1121_/Y _1943_/B _1946_/X _1944_/X vssd1 vssd1 vccd1 vccd1 _2354_/D sky130_fd_sc_hd__a211o_1
XFILLER_174_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1878_ _2362_/Q _2238_/A vssd1 vssd1 vccd1 vccd1 _1878_/X sky130_fd_sc_hd__xor2_1
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1801_ _2469_/Q vssd1 vssd1 vccd1 vccd1 _1801_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1732_ _2399_/Q _1728_/Y _1845_/A _1730_/Y _1731_/X vssd1 vssd1 vccd1 vccd1 _1732_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1663_ _1663_/A _1663_/B vssd1 vssd1 vccd1 vccd1 _1664_/C sky130_fd_sc_hd__or2_1
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1594_ _2303_/Q _1596_/C _1613_/A vssd1 vssd1 vccd1 vccd1 _1595_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2215_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2450_/D sky130_fd_sc_hd__clkbuf_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2146_ _1708_/Y _2142_/X _2145_/X vssd1 vssd1 vccd1 vccd1 _2420_/D sky130_fd_sc_hd__a21oi_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2077_ _2076_/Y _2396_/Q vssd1 vssd1 vccd1 vccd1 _2077_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _2371_/Q _1990_/X _1966_/X vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__a21o_1
XFILLER_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1715_ _1719_/A _1726_/A vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__and2b_1
XFILLER_172_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1646_ _2318_/Q _1646_/B _1650_/A _1648_/B vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__or4_1
X_1577_ _2300_/Q _2299_/Q _2298_/Q _1577_/D vssd1 vssd1 vccd1 vccd1 _1579_/A sky130_fd_sc_hd__and4_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2129_ _2102_/A _2121_/B _2118_/X vssd1 vssd1 vccd1 vccd1 _2129_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1500_ input44/X _1484_/X _1477_/X _1499_/X vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__o211a_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1431_ _1431_/A1 _1421_/X _1417_/X _1430_/X vssd1 vssd1 vccd1 vccd1 _1431_/X sky130_fd_sc_hd__o211a_4
XFILLER_141_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1362_ _1362_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__and2_1
X_1293_ _1327_/A _1327_/B _1293_/C vssd1 vssd1 vccd1 vccd1 _1293_/X sky130_fd_sc_hd__and3_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput190 sram_dout1[43] vssd1 vssd1 vccd1 vccd1 _1328_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1629_ _1629_/A _1634_/D vssd1 vssd1 vccd1 vccd1 _1631_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1980_ _1124_/X _1976_/X _1979_/X _1944_/X vssd1 vssd1 vccd1 vccd1 _2364_/D sky130_fd_sc_hd__a211o_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ _2474_/A _2463_/D vssd1 vssd1 vccd1 vccd1 _2463_/Q sky130_fd_sc_hd__dfxtp_1
X_1414_ input57/X _1409_/X _1410_/X input92/X vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__a22o_1
X_2394_ _2468_/CLK _2394_/D vssd1 vssd1 vccd1 vccd1 _2394_/Q sky130_fd_sc_hd__dfxtp_1
X_1345_ _1345_/A _1353_/B vssd1 vssd1 vccd1 vccd1 _1346_/A sky130_fd_sc_hd__and2_1
X_1276_ _1276_/A1 _1215_/A _1235_/A _1276_/B2 vssd1 vssd1 vccd1 vccd1 _1276_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2472_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1130_ _2472_/Q _2471_/Q vssd1 vssd1 vccd1 vccd1 _1136_/B sky130_fd_sc_hd__or2_1
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1963_ _1111_/X _1957_/X _1962_/X vssd1 vssd1 vccd1 vccd1 _2358_/D sky130_fd_sc_hd__a21o_1
XFILLER_159_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1894_ _2456_/Q _2457_/Q _2458_/Q _2459_/Q vssd1 vssd1 vccd1 vccd1 _1909_/C sky130_fd_sc_hd__or4_2
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2446_ _2446_/CLK _2446_/D vssd1 vssd1 vccd1 vccd1 _2446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2377_ _2474_/A _2377_/D vssd1 vssd1 vccd1 vccd1 _2377_/Q sky130_fd_sc_hd__dfxtp_1
X_1328_ _1328_/A1 _1287_/A _1224_/A _1328_/B2 _1327_/X vssd1 vssd1 vccd1 vccd1 _1328_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1259_ _1259_/A _1259_/B vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__or2_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2300_ _2319_/CLK _2300_/D vssd1 vssd1 vccd1 vccd1 _2300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2231_ _2458_/Q _2231_/A1 _2231_/S vssd1 vssd1 vccd1 vccd1 _2232_/A sky130_fd_sc_hd__mux2_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2162_ _2162_/A _2167_/B _2162_/C vssd1 vssd1 vccd1 vccd1 _2164_/A sky130_fd_sc_hd__nor3_2
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1113_ _2171_/A vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__clkinv_4
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2093_ _2093_/A _2100_/B vssd1 vssd1 vccd1 vccd1 _2093_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1946_ _1938_/A _2354_/Q vssd1 vssd1 vccd1 vccd1 _1946_/X sky130_fd_sc_hd__and2b_1
XFILLER_174_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1877_ _2355_/Q vssd1 vssd1 vccd1 vccd1 _1877_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2429_ _2434_/CLK _2429_/D vssd1 vssd1 vccd1 vccd1 _2429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1800_ _1800_/A vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__buf_2
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1731_ _2404_/Q _2332_/Q vssd1 vssd1 vccd1 vccd1 _1731_/X sky130_fd_sc_hd__xor2_1
X_1662_ _1663_/A _1663_/B vssd1 vssd1 vccd1 vccd1 _1664_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1593_ _2303_/Q _1596_/C vssd1 vssd1 vccd1 vccd1 _1595_/A sky130_fd_sc_hd__and2_1
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2450_/Q _2214_/A1 _2220_/S vssd1 vssd1 vccd1 vccd1 _2215_/A sky130_fd_sc_hd__mux2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2145_ _2171_/A _2138_/A _1952_/X vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2076_ _2157_/A _2085_/B _2157_/C vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__nor3_2
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1929_ _2349_/Q _1918_/X _1928_/Y vssd1 vssd1 vccd1 vccd1 _2349_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2337_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1714_ _1568_/D _1714_/B vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__and2b_1
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1645_ _1645_/A vssd1 vssd1 vccd1 vccd1 _2317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1576_ _1576_/A _1576_/B vssd1 vssd1 vccd1 vccd1 _2299_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _2414_/Q _2111_/X _2127_/Y vssd1 vssd1 vccd1 vccd1 _2414_/D sky130_fd_sc_hd__o21a_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2059_ _2089_/A _2053_/A _1952_/X vssd1 vssd1 vccd1 vccd1 _2059_/X sky130_fd_sc_hd__a21o_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1430_ input5/X _1407_/X _1408_/X _1429_/X vssd1 vssd1 vccd1 vccd1 _1430_/X sky130_fd_sc_hd__a211o_2
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1361_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1361_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1292_ _1234_/A _1289_/X _1291_/X _1233_/A vssd1 vssd1 vccd1 vccd1 _1298_/A sky130_fd_sc_hd__a22o_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput180 sram_dout1[34] vssd1 vssd1 vccd1 vccd1 _1279_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput191 sram_dout1[44] vssd1 vssd1 vccd1 vccd1 _1225_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1628_ _1629_/A _1634_/D vssd1 vssd1 vccd1 vccd1 _1628_/X sky130_fd_sc_hd__or2_1
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1559_ _1559_/A _1559_/B _1559_/C _1559_/D vssd1 vssd1 vccd1 vccd1 _1568_/D sky130_fd_sc_hd__and4_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2462_ _2474_/A _2462_/D vssd1 vssd1 vccd1 vccd1 _2462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2393_ _2468_/CLK _2393_/D vssd1 vssd1 vccd1 vccd1 _2393_/Q sky130_fd_sc_hd__dfxtp_1
X_1413_ input51/X _1385_/X _1398_/X _1412_/X vssd1 vssd1 vccd1 vccd1 _1413_/X sky130_fd_sc_hd__o211a_4
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1344_ _1379_/B vssd1 vssd1 vccd1 vccd1 _1353_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1275_ _1275_/A _1275_/B vssd1 vssd1 vccd1 vccd1 _1275_/X sky130_fd_sc_hd__or2_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1962_ _2358_/Q _1950_/X _2185_/A vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1893_ _2442_/Q _2443_/Q _2444_/Q _2445_/Q vssd1 vssd1 vccd1 vccd1 _1909_/B sky130_fd_sc_hd__or4_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2445_ _2446_/CLK _2445_/D vssd1 vssd1 vccd1 vccd1 _2445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _2459_/CLK _2376_/D vssd1 vssd1 vccd1 vccd1 _2376_/Q sky130_fd_sc_hd__dfxtp_1
X_1327_ _1327_/A _1327_/B _1327_/C vssd1 vssd1 vccd1 vccd1 _1327_/X sky130_fd_sc_hd__and3_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1258_ _1223_/X _1255_/X _1257_/X _1240_/A _1229_/X vssd1 vssd1 vccd1 vccd1 _1259_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1189_ _1287_/A vssd1 vssd1 vccd1 vccd1 _1190_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2230_ _2230_/A vssd1 vssd1 vccd1 vccd1 _2457_/D sky130_fd_sc_hd__clkbuf_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2161_ _2427_/Q _2158_/B _2160_/Y vssd1 vssd1 vccd1 vccd1 _2427_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1112_ _1112_/A _1118_/B vssd1 vssd1 vccd1 vccd1 _2171_/A sky130_fd_sc_hd__nand2_8
X_2092_ _2400_/Q _2085_/Y _2091_/Y vssd1 vssd1 vccd1 vccd1 _2400_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _1124_/X _1943_/B _1943_/Y _1944_/X vssd1 vssd1 vccd1 vccd1 _2353_/D sky130_fd_sc_hd__a211o_1
XFILLER_174_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1876_ _1874_/Y _2238_/B _1801_/Y _2353_/Q _1875_/X vssd1 vssd1 vccd1 vccd1 _1885_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2428_ _2434_/CLK _2428_/D vssd1 vssd1 vccd1 vccd1 _2428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2359_ _2435_/CLK _2359_/D vssd1 vssd1 vccd1 vccd1 _2359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1730_ _2398_/Q vssd1 vssd1 vccd1 vccd1 _1730_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1661_ _2323_/Q vssd1 vssd1 vccd1 vccd1 _1663_/A sky130_fd_sc_hd__inv_2
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ _1592_/A vssd1 vssd1 vccd1 vccd1 _2302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2213_ _2213_/A vssd1 vssd1 vccd1 vccd1 _2449_/D sky130_fd_sc_hd__clkbuf_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _1117_/X _2137_/X _2143_/X vssd1 vssd1 vccd1 vccd1 _2419_/D sky130_fd_sc_hd__a21o_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _2167_/C vssd1 vssd1 vccd1 vccd1 _2157_/C sky130_fd_sc_hd__buf_2
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1928_ _2098_/A _1922_/B _1919_/X vssd1 vssd1 vccd1 vccd1 _1928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ _2394_/Q _1815_/Y _1800_/A _2392_/Q vssd1 vssd1 vccd1 vccd1 _1859_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _2325_/Q vssd1 vssd1 vccd1 vccd1 _1719_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1644_ _1644_/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1645_/A sky130_fd_sc_hd__and2_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1575_ _2299_/Q _1573_/A _1714_/B vssd1 vssd1 vccd1 vccd1 _1576_/B sky130_fd_sc_hd__o21ai_1
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2127_ _2100_/A _2121_/B _2118_/X vssd1 vssd1 vccd1 vccd1 _2127_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2058_ _2058_/A vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__clkbuf_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1360_ _1360_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1361_/A sky130_fd_sc_hd__and2_1
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1291_ _1291_/A1 _1321_/B _1224_/X _1291_/B2 _1290_/X vssd1 vssd1 vccd1 vccd1 _1291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput181 sram_dout1[35] vssd1 vssd1 vccd1 vccd1 _1282_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput170 sram_dout1[23] vssd1 vssd1 vccd1 vccd1 _1320_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput192 sram_dout1[45] vssd1 vssd1 vccd1 vccd1 _1255_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1627_ _1615_/X _1625_/Y _1626_/X _1622_/X _2312_/Q vssd1 vssd1 vccd1 vccd1 _2312_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_160_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1558_ _2344_/Q _2328_/Q vssd1 vssd1 vccd1 vccd1 _1559_/D sky130_fd_sc_hd__xnor2_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1489_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1489_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2461_ _2468_/CLK _2461_/D vssd1 vssd1 vccd1 vccd1 _2461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1412_ _1412_/A1 _1407_/X _1408_/X _1411_/X vssd1 vssd1 vccd1 vccd1 _1412_/X sky130_fd_sc_hd__a211o_2
X_2392_ _2468_/CLK _2392_/D vssd1 vssd1 vccd1 vccd1 _2392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1343_ _1343_/A vssd1 vssd1 vccd1 vccd1 _1343_/X sky130_fd_sc_hd__clkbuf_1
X_1274_ _1223_/X _1271_/X _1273_/X _1240_/A _1229_/X vssd1 vssd1 vccd1 vccd1 _1275_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2185_/A sky130_fd_sc_hd__clkbuf_4
X_1892_ _2440_/Q _1898_/A _2441_/Q vssd1 vssd1 vccd1 vccd1 _1911_/C sky130_fd_sc_hd__or3b_2
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2444_ _2472_/CLK _2444_/D vssd1 vssd1 vccd1 vccd1 _2444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2375_ _2459_/CLK _2375_/D vssd1 vssd1 vccd1 vccd1 _2375_/Q sky130_fd_sc_hd__dfxtp_1
X_1326_ _1235_/X _1325_/X _1229_/X vssd1 vssd1 vccd1 vccd1 _1332_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1257_ _1257_/A1 _1201_/X _1202_/X _1257_/B2 _1256_/X vssd1 vssd1 vccd1 vccd1 _1257_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1188_ _2293_/Q _2294_/Q vssd1 vssd1 vccd1 vccd1 _1287_/A sky130_fd_sc_hd__and2b_1
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_0 _1147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2160_ _2049_/X _2158_/B _2139_/X vssd1 vssd1 vccd1 vccd1 _2160_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2091_ _1958_/X _2085_/Y _2079_/X vssd1 vssd1 vccd1 vccd1 _2091_/Y sky130_fd_sc_hd__a21oi_1
X_1111_ _1111_/A vssd1 vssd1 vccd1 vccd1 _1111_/X sky130_fd_sc_hd__buf_6
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _2116_/A vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1875_ _2354_/Q _2267_/C vssd1 vssd1 vccd1 vccd1 _1875_/X sky130_fd_sc_hd__xor2_1
XFILLER_174_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2427_ _2435_/CLK _2427_/D vssd1 vssd1 vccd1 vccd1 _2427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2358_ _2425_/CLK _2358_/D vssd1 vssd1 vccd1 vccd1 _2358_/Q sky130_fd_sc_hd__dfxtp_1
X_1309_ _1309_/A1 _1216_/X _1217_/X _1309_/B2 _1308_/X vssd1 vssd1 vccd1 vccd1 _1309_/X
+ sky130_fd_sc_hd__a221o_1
X_2289_ _2475_/A _2289_/D vssd1 vssd1 vccd1 vccd1 _2289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1660_ _1660_/A vssd1 vssd1 vccd1 vccd1 _2322_/D sky130_fd_sc_hd__clkbuf_1
X_1591_ _1596_/C _1613_/A _1591_/C vssd1 vssd1 vccd1 vccd1 _1592_/A sky130_fd_sc_hd__and3b_1
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2212_ _2449_/Q _2212_/A1 _2220_/S vssd1 vssd1 vccd1 vccd1 _2213_/A sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2143_ _2419_/Q _2142_/X _2071_/X vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2074_ _2441_/Q _2074_/B _2074_/C _2074_/D vssd1 vssd1 vccd1 vccd1 _2167_/C sky130_fd_sc_hd__or4_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1927_ _2348_/Q _1912_/Y _1926_/X _1916_/X vssd1 vssd1 vccd1 vccd1 _2348_/D sky130_fd_sc_hd__a211o_1
XFILLER_147_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1858_ _2394_/Q vssd1 vssd1 vccd1 vccd1 _1858_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1789_ _1779_/X _1784_/X _1789_/C _1789_/D vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__and4bb_1
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1712_ _1668_/X _1669_/X _1674_/X _1691_/X _1711_/X vssd1 vssd1 vccd1 vccd1 _2324_/D
+ sky130_fd_sc_hd__o41a_1
X_1643_ _1639_/A _1615_/A _1641_/C _2317_/Q vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__a31o_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1574_ _2299_/Q _2298_/Q _1577_/D vssd1 vssd1 vccd1 vccd1 _1576_/A sky130_fd_sc_hd__and3_1
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2126_ _2413_/Q _2111_/X _2125_/Y vssd1 vssd1 vccd1 vccd1 _2413_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2057_/A _2057_/B _2057_/C vssd1 vssd1 vccd1 vccd1 _2058_/A sky130_fd_sc_hd__or3_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1290_ _1308_/A _1308_/B _1290_/C vssd1 vssd1 vccd1 vccd1 _1290_/X sky130_fd_sc_hd__and3_1
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput171 sram_dout1[24] vssd1 vssd1 vccd1 vccd1 _1236_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput160 sram_dout1[14] vssd1 vssd1 vccd1 vccd1 _1276_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput193 sram_dout1[46] vssd1 vssd1 vccd1 vccd1 _1270_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput182 sram_dout1[36] vssd1 vssd1 vccd1 vccd1 _1315_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _1621_/A _1621_/B _1621_/C _2312_/Q vssd1 vssd1 vccd1 vccd1 _1626_/X sky130_fd_sc_hd__a31o_1
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1557_ _2347_/Q _2325_/Q vssd1 vssd1 vccd1 vccd1 _1559_/C sky130_fd_sc_hd__xnor2_1
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1488_ input41/X _1484_/X _1477_/X _1487_/X vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__o211a_4
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2109_ _2167_/A _2109_/B _2162_/C vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__nor3_2
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2460_ _2468_/CLK _2460_/D vssd1 vssd1 vccd1 vccd1 _2460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1411_ input56/X _1409_/X _1410_/X input91/X vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2391_ _2468_/CLK _2391_/D vssd1 vssd1 vccd1 vccd1 _2391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1342_ _1342_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _1343_/A sky130_fd_sc_hd__and2_1
X_1273_ _1273_/A1 _1216_/X _1217_/X _1273_/B2 _1272_/X vssd1 vssd1 vccd1 vccd1 _1273_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1609_ _1609_/A _1609_/B _1609_/C vssd1 vssd1 vccd1 vccd1 _1609_/X sky130_fd_sc_hd__and3_1
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ _2357_/Q _1957_/X _1959_/Y vssd1 vssd1 vccd1 vccd1 _2357_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1891_ _2439_/Q _2040_/C _2040_/B vssd1 vssd1 vccd1 vccd1 _1949_/B sky130_fd_sc_hd__or3b_4
XFILLER_174_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2443_ _2446_/CLK _2443_/D vssd1 vssd1 vccd1 vccd1 _2443_/Q sky130_fd_sc_hd__dfxtp_1
X_2374_ _2459_/CLK _2374_/D vssd1 vssd1 vccd1 vccd1 _2374_/Q sky130_fd_sc_hd__dfxtp_1
X_1325_ _1325_/A1 _1321_/B _1224_/X _1325_/B2 _1324_/X vssd1 vssd1 vccd1 vccd1 _1325_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1256_ _1301_/A _1301_/B _1256_/C vssd1 vssd1 vccd1 vccd1 _1256_/X sky130_fd_sc_hd__and3_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1187_ _1187_/A vssd1 vssd1 vccd1 vccd1 _1187_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1110_ _2093_/A vssd1 vssd1 vccd1 vccd1 _1111_/A sky130_fd_sc_hd__inv_2
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ _2399_/Q _2084_/X _2089_/Y _2016_/X vssd1 vssd1 vccd1 vccd1 _2399_/D sky130_fd_sc_hd__a211o_1
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2446_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ _1943_/A _1943_/B vssd1 vssd1 vccd1 vccd1 _1943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1874_ _2361_/Q vssd1 vssd1 vccd1 vccd1 _1874_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2426_ _2434_/CLK _2426_/D vssd1 vssd1 vccd1 vccd1 _2426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2357_ _2435_/CLK _2357_/D vssd1 vssd1 vccd1 vccd1 _2357_/Q sky130_fd_sc_hd__dfxtp_1
X_1308_ _1308_/A _1308_/B _1308_/C vssd1 vssd1 vccd1 vccd1 _1308_/X sky130_fd_sc_hd__and3_1
X_2288_ _2475_/A _2288_/D vssd1 vssd1 vccd1 vccd1 _2288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1239_ _1609_/A _1239_/B vssd1 vssd1 vccd1 vccd1 _1240_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1590_ _1240_/A _1656_/B _2302_/Q vssd1 vssd1 vccd1 vccd1 _1591_/C sky130_fd_sc_hd__a21o_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2211_ _2233_/S vssd1 vssd1 vccd1 vccd1 _2220_/S sky130_fd_sc_hd__clkbuf_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2142_ _2162_/A _2142_/B _2162_/C vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__or3_2
X_2073_ _1098_/X _2054_/A _2072_/X vssd1 vssd1 vccd1 vccd1 _2395_/D sky130_fd_sc_hd__a21o_1
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1926_ _1926_/A _1930_/B vssd1 vssd1 vccd1 vccd1 _1926_/X sky130_fd_sc_hd__and2_1
XFILLER_135_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1857_ _2395_/Q vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1788_ _1768_/Y _2465_/Q _2468_/Q _1770_/Y _1787_/X vssd1 vssd1 vccd1 vccd1 _1789_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2409_ _2425_/CLK _2409_/D vssd1 vssd1 vccd1 vccd1 _2409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1711_ _1693_/X _1695_/Y _1701_/X _1710_/X _2324_/Q vssd1 vssd1 vccd1 vccd1 _1711_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1642_ _1615_/A _1648_/B _1648_/A vssd1 vssd1 vccd1 vccd1 _1644_/A sky130_fd_sc_hd__a21o_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1573_ _1573_/A _1573_/B vssd1 vssd1 vccd1 vccd1 _2298_/D sky130_fd_sc_hd__nor2_1
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2125_ _2098_/A _2121_/B _2118_/X vssd1 vssd1 vccd1 vccd1 _2125_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2056_ _2388_/Q _2054_/X _2055_/Y vssd1 vssd1 vccd1 vccd1 _2388_/D sky130_fd_sc_hd__o21a_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1909_ _1909_/A _1909_/B _1909_/C _1909_/D vssd1 vssd1 vccd1 vccd1 _2074_/D sky130_fd_sc_hd__or4_1
XFILLER_163_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput150 sram_dout1[119] vssd1 vssd1 vccd1 vccd1 _1329_/C sky130_fd_sc_hd__clkbuf_2
Xinput172 sram_dout1[25] vssd1 vssd1 vccd1 vccd1 _1260_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput161 sram_dout1[15] vssd1 vssd1 vccd1 vccd1 _1285_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput183 sram_dout1[37] vssd1 vssd1 vccd1 vccd1 _1318_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput194 sram_dout1[47] vssd1 vssd1 vccd1 vccd1 _1294_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1625_ _1634_/D vssd1 vssd1 vccd1 vccd1 _1625_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1556_ _2346_/Q _2326_/Q vssd1 vssd1 vccd1 vccd1 _1559_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1487_ _1487_/A1 _1432_/X _1486_/X _1435_/X vssd1 vssd1 vccd1 vccd1 _1487_/X sky130_fd_sc_hd__a211o_2
XFILLER_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _2407_/Q _2105_/B _2107_/Y vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2039_ _1098_/X _2019_/X _2038_/X vssd1 vssd1 vccd1 vccd1 _2384_/D sky130_fd_sc_hd__a21o_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2414_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1410_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1410_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2390_ _2435_/CLK _2390_/D vssd1 vssd1 vccd1 vccd1 _2390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1341_ _1341_/A vssd1 vssd1 vccd1 vccd1 _1341_/X sky130_fd_sc_hd__clkbuf_1
X_1272_ _1301_/A _1301_/B _1272_/C vssd1 vssd1 vccd1 vccd1 _1272_/X sky130_fd_sc_hd__and3_1
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput410 _1416_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_172_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1608_ _1609_/B _1609_/C _1607_/Y vssd1 vssd1 vccd1 vccd1 _2307_/D sky130_fd_sc_hd__a21oi_1
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1539_ _1140_/A _1518_/X _1404_/X vssd1 vssd1 vccd1 vccd1 _1539_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1890_ _2446_/Q _2447_/Q _1099_/A vssd1 vssd1 vccd1 vccd1 _2040_/C sky130_fd_sc_hd__or3b_2
XFILLER_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2442_ _2446_/CLK _2442_/D vssd1 vssd1 vccd1 vccd1 _2442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2373_ _2474_/A _2373_/D vssd1 vssd1 vccd1 vccd1 _2373_/Q sky130_fd_sc_hd__dfxtp_1
X_1324_ _1329_/A _1329_/B _1324_/C vssd1 vssd1 vccd1 vccd1 _1324_/X sky130_fd_sc_hd__and3_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1255_ _1255_/A1 _1216_/X _1217_/X _1255_/B2 _1254_/X vssd1 vssd1 vccd1 vccd1 _1255_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1186_ _1327_/A _1327_/B vssd1 vssd1 vccd1 vccd1 _1187_/A sky130_fd_sc_hd__and2_2
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_2 _1238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1942_ _2352_/Q _1943_/B _1941_/Y vssd1 vssd1 vccd1 vccd1 _2352_/D sky130_fd_sc_hd__o21a_1
X_1873_ _1869_/Y _2261_/A _2272_/A _1943_/A _1872_/X vssd1 vssd1 vccd1 vccd1 _1873_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2425_ _2425_/CLK _2425_/D vssd1 vssd1 vccd1 vccd1 _2425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2356_ _2425_/CLK _2356_/D vssd1 vssd1 vccd1 vccd1 _2356_/Q sky130_fd_sc_hd__dfxtp_1
X_1307_ _1307_/A1 _1216_/X _1217_/X _1307_/B2 _1306_/X vssd1 vssd1 vccd1 vccd1 _1307_/X
+ sky130_fd_sc_hd__a221o_1
X_2287_ _2475_/A _2287_/D vssd1 vssd1 vccd1 vccd1 _2287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1238_ _1314_/A _1238_/B vssd1 vssd1 vccd1 vccd1 _1238_/X sky130_fd_sc_hd__or2_1
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1169_ _1169_/A vssd1 vssd1 vccd1 vccd1 _2288_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2210_ _2210_/A vssd1 vssd1 vccd1 vccd1 _2448_/D sky130_fd_sc_hd__clkbuf_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2141_ _2418_/Q _2137_/X _2140_/Y vssd1 vssd1 vccd1 vccd1 _2418_/D sky130_fd_sc_hd__o21a_1
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2072_ _2395_/Q _2058_/A _2071_/X vssd1 vssd1 vccd1 vccd1 _2072_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1925_ _2347_/Q _1918_/X _1924_/Y vssd1 vssd1 vccd1 vccd1 _2347_/D sky130_fd_sc_hd__o21a_1
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1856_ _2395_/Q _2235_/A _2470_/Q _2044_/A _1855_/X vssd1 vssd1 vccd1 vccd1 _1866_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1787_ _1775_/Y _2463_/Q _1794_/A _2369_/Q vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2408_ _2446_/CLK _2408_/D vssd1 vssd1 vccd1 vccd1 _2408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2339_ _2434_/CLK _2339_/D vssd1 vssd1 vccd1 vccd1 _2339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput310 wb_we_i vssd1 vssd1 vccd1 vccd1 _2279_/A1 sky130_fd_sc_hd__buf_2
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1710_ _1704_/X _1710_/B _1710_/C _1710_/D vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__and4b_1
X_1641_ _2316_/Q _2317_/Q _1641_/C vssd1 vssd1 vccd1 vccd1 _1648_/B sky130_fd_sc_hd__nand3_1
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1572_ _2298_/Q _1577_/D _1562_/X vssd1 vssd1 vccd1 vccd1 _1573_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2124_ _1108_/X _2112_/X _2123_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _2412_/D sky130_fd_sc_hd__a211o_1
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2055_ _1985_/X _2054_/A _2030_/X vssd1 vssd1 vccd1 vccd1 _2055_/Y sky130_fd_sc_hd__a21oi_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1908_ _2449_/Q _2450_/Q vssd1 vssd1 vccd1 vccd1 _1909_/D sky130_fd_sc_hd__or2_1
XFILLER_163_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1839_ _1839_/A _1839_/B vssd1 vssd1 vccd1 vccd1 _1845_/C sky130_fd_sc_hd__and2_1
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput151 sram_dout1[11] vssd1 vssd1 vccd1 vccd1 _1320_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput162 sram_dout1[16] vssd1 vssd1 vccd1 vccd1 _1312_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput140 sram_dout1[10] vssd1 vssd1 vccd1 vccd1 _1313_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput173 sram_dout1[26] vssd1 vssd1 vccd1 vccd1 _1276_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput195 sram_dout1[48] vssd1 vssd1 vccd1 vccd1 _1307_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput184 sram_dout1[38] vssd1 vssd1 vccd1 vccd1 _1206_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1624_ _2309_/Q _2310_/Q _2311_/Q _2312_/Q vssd1 vssd1 vccd1 vccd1 _1634_/D sky130_fd_sc_hd__and4_1
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1555_ _2345_/Q _2327_/Q vssd1 vssd1 vccd1 vccd1 _1559_/A sky130_fd_sc_hd__xnor2_1
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1486_ input19/X _1485_/X _1433_/X input76/X vssd1 vssd1 vccd1 vccd1 _1486_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2107_ _2049_/X _2105_/B _2079_/X vssd1 vssd1 vccd1 vccd1 _2107_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2384_/Q _2023_/X _2037_/X vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1340_ _1340_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _1341_/A sky130_fd_sc_hd__and2_1
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1271_ _1271_/A1 _1187_/A _1270_/X vssd1 vssd1 vccd1 vccd1 _1271_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput411 _1420_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[4] sky130_fd_sc_hd__buf_2
Xoutput400 _1500_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_173_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1607_ _1609_/B _1609_/C _1613_/A vssd1 vssd1 vccd1 vccd1 _1607_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1538_ _1538_/A vssd1 vssd1 vccd1 vccd1 _1538_/X sky130_fd_sc_hd__clkbuf_1
X_1469_ input36/X _1463_/X _1459_/X _1468_/X vssd1 vssd1 vccd1 vccd1 _1469_/X sky130_fd_sc_hd__o211a_4
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2441_ _2446_/CLK _2441_/D vssd1 vssd1 vccd1 vccd1 _2441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2372_ _2474_/A _2372_/D vssd1 vssd1 vccd1 vccd1 _2372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1323_ _1321_/X _1322_/X _1284_/X vssd1 vssd1 vccd1 vccd1 _1332_/A sky130_fd_sc_hd__o21a_1
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1254_ _1308_/A _1308_/B _1254_/C vssd1 vssd1 vccd1 vccd1 _1254_/X sky130_fd_sc_hd__and3_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1185_ _2293_/Q vssd1 vssd1 vccd1 vccd1 _1327_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_3 _1262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _1126_/A _1943_/B _1940_/X vssd1 vssd1 vccd1 vccd1 _1941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1872_ _2360_/Q _2243_/A _2275_/A _2352_/Q _1871_/X vssd1 vssd1 vccd1 vccd1 _1872_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2424_ _2435_/CLK _2424_/D vssd1 vssd1 vccd1 vccd1 _2424_/Q sky130_fd_sc_hd__dfxtp_1
X_2355_ _2435_/CLK _2355_/D vssd1 vssd1 vccd1 vccd1 _2355_/Q sky130_fd_sc_hd__dfxtp_1
X_1306_ _1308_/A _1308_/B _1306_/C vssd1 vssd1 vccd1 vccd1 _1306_/X sky130_fd_sc_hd__and3_1
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2286_ _2475_/A _2286_/D vssd1 vssd1 vccd1 vccd1 _2286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1237_ _1237_/A1 _1233_/X _1234_/X _1237_/B2 _1236_/X vssd1 vssd1 vccd1 vccd1 _1238_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1168_ _2295_/Q _1629_/A _1168_/S vssd1 vssd1 vccd1 vccd1 _1169_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1099_ _1099_/A vssd1 vssd1 vccd1 vccd1 _1122_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2140_ _1985_/X _2138_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__a21oi_1
X_2071_ _2071_/A vssd1 vssd1 vccd1 vccd1 _2071_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1924_ _2093_/A _1922_/B _1919_/X vssd1 vssd1 vccd1 vccd1 _1924_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1855_ _2391_/Q _1794_/A _1781_/A _2388_/Q vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__a22o_1
X_1786_ _2464_/Q vssd1 vssd1 vccd1 vccd1 _1794_/A sky130_fd_sc_hd__clkinv_2
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2407_ _2452_/CLK _2407_/D vssd1 vssd1 vccd1 vccd1 _2407_/Q sky130_fd_sc_hd__dfxtp_1
X_2338_ _2434_/CLK _2338_/D vssd1 vssd1 vccd1 vccd1 _2338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2269_ _2273_/A _2269_/B _2269_/C vssd1 vssd1 vccd1 vccd1 _2270_/A sky130_fd_sc_hd__and3_1
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput300 wb_data_i[6] vssd1 vssd1 vccd1 vccd1 _1115_/A sky130_fd_sc_hd__buf_2
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1640_ _1615_/A _1638_/Y _1639_/X _1622_/X _1639_/A vssd1 vssd1 vccd1 vccd1 _2316_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1571_ _2298_/Q _1577_/D vssd1 vssd1 vccd1 vccd1 _1573_/A sky130_fd_sc_hd__and2_1
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2123_ _2112_/A _2412_/Q vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__and2b_1
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2054_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1907_ _2448_/Q _2451_/Q _1907_/C vssd1 vssd1 vccd1 vccd1 _2074_/C sky130_fd_sc_hd__or3_1
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1838_ _1846_/A _1839_/B _1838_/C vssd1 vssd1 vccd1 vccd1 _2336_/D sky130_fd_sc_hd__nor3_1
XFILLER_163_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1769_ _2468_/Q vssd1 vssd1 vccd1 vccd1 _2267_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_173_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput152 sram_dout1[120] vssd1 vssd1 vccd1 vccd1 _1220_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 sram_dout1[110] vssd1 vssd1 vccd1 vccd1 _1271_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput130 sram_dout1[100] vssd1 vssd1 vccd1 vccd1 _1315_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 sram_dout1[17] vssd1 vssd1 vccd1 vccd1 _1319_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput185 sram_dout1[39] vssd1 vssd1 vccd1 vccd1 _1252_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput174 sram_dout1[27] vssd1 vssd1 vccd1 vccd1 _1285_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput196 sram_dout1[49] vssd1 vssd1 vccd1 vccd1 _1325_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1623_ _1615_/X _1620_/X _1621_/Y _1622_/X _1621_/C vssd1 vssd1 vccd1 vccd1 _2311_/D
+ sky130_fd_sc_hd__a32o_1
X_1554_ _1554_/A vssd1 vssd1 vccd1 vccd1 _2283_/D sky130_fd_sc_hd__clkbuf_1
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

