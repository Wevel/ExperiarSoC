VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 500.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 496.000 27.510 500.000 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 496.000 32.110 500.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 496.000 36.250 500.000 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 496.000 40.390 500.000 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 496.000 44.530 500.000 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 496.000 49.130 500.000 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 496.000 53.270 500.000 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 496.000 57.410 500.000 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 496.000 62.010 500.000 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 496.000 481.070 500.000 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 496.000 485.210 500.000 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 496.000 489.810 500.000 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 496.000 493.950 500.000 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 496.000 498.090 500.000 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 496.000 502.690 500.000 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 496.000 506.830 500.000 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 496.000 510.970 500.000 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 496.000 515.110 500.000 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 496.000 2.210 500.000 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 496.000 476.930 500.000 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 5.480 800.000 6.080 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 19.760 800.000 20.360 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 103.400 800.000 104.000 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 110.880 800.000 111.480 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 117.680 800.000 118.280 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 125.160 800.000 125.760 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 132.640 800.000 133.240 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 140.120 800.000 140.720 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 147.600 800.000 148.200 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 154.400 800.000 155.000 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 161.880 800.000 162.480 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 169.360 800.000 169.960 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 29.960 800.000 30.560 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 184.320 800.000 184.920 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 191.800 800.000 192.400 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 198.600 800.000 199.200 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 206.080 800.000 206.680 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 213.560 800.000 214.160 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 221.040 800.000 221.640 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 228.520 800.000 229.120 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 39.480 800.000 40.080 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 49.680 800.000 50.280 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 59.200 800.000 59.800 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 66.680 800.000 67.280 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 74.160 800.000 74.760 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 80.960 800.000 81.560 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 88.440 800.000 89.040 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 95.920 800.000 96.520 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 7.520 800.000 8.120 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 22.480 800.000 23.080 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 105.440 800.000 106.040 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 112.920 800.000 113.520 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 120.400 800.000 121.000 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 127.880 800.000 128.480 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 135.360 800.000 135.960 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 142.160 800.000 142.760 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 149.640 800.000 150.240 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 157.120 800.000 157.720 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 164.600 800.000 165.200 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 172.080 800.000 172.680 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 32.000 800.000 32.600 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 179.560 800.000 180.160 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 186.360 800.000 186.960 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 193.840 800.000 194.440 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 201.320 800.000 201.920 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 208.800 800.000 209.400 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 216.280 800.000 216.880 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 223.080 800.000 223.680 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 230.560 800.000 231.160 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 235.320 800.000 235.920 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 240.760 800.000 241.360 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 42.200 800.000 42.800 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 245.520 800.000 246.120 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 250.280 800.000 250.880 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.720 800.000 52.320 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 61.920 800.000 62.520 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 68.720 800.000 69.320 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 76.200 800.000 76.800 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 83.680 800.000 84.280 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 91.160 800.000 91.760 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 98.640 800.000 99.240 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 25.200 800.000 25.800 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 108.160 800.000 108.760 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 115.640 800.000 116.240 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 123.120 800.000 123.720 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 129.920 800.000 130.520 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 137.400 800.000 138.000 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 144.880 800.000 145.480 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 152.360 800.000 152.960 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 159.840 800.000 160.440 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 167.320 800.000 167.920 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 174.120 800.000 174.720 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 34.720 800.000 35.320 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 181.600 800.000 182.200 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 189.080 800.000 189.680 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 196.560 800.000 197.160 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 204.040 800.000 204.640 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 218.320 800.000 218.920 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 225.800 800.000 226.400 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 233.280 800.000 233.880 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 238.040 800.000 238.640 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 242.800 800.000 243.400 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 44.240 800.000 44.840 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 247.560 800.000 248.160 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 253.000 800.000 253.600 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 54.440 800.000 55.040 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 63.960 800.000 64.560 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 71.440 800.000 72.040 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 78.920 800.000 79.520 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 86.400 800.000 87.000 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 93.200 800.000 93.800 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 100.680 800.000 101.280 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 10.240 800.000 10.840 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 27.240 800.000 27.840 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 37.440 800.000 38.040 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 46.960 800.000 47.560 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 56.480 800.000 57.080 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 12.960 800.000 13.560 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 15.000 800.000 15.600 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 17.720 800.000 18.320 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 496.000 793.410 500.000 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 496.000 797.550 500.000 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 497.800 800.000 498.400 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 496.000 66.150 500.000 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 496.000 108.930 500.000 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 496.000 113.070 500.000 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 496.000 117.670 500.000 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 496.000 121.810 500.000 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 496.000 125.950 500.000 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 496.000 130.090 500.000 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 496.000 134.690 500.000 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 496.000 138.830 500.000 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 496.000 142.970 500.000 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 496.000 147.570 500.000 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 496.000 70.290 500.000 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 496.000 151.710 500.000 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 496.000 155.850 500.000 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 496.000 160.450 500.000 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 496.000 164.590 500.000 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 496.000 168.730 500.000 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 496.000 172.870 500.000 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 496.000 177.470 500.000 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 496.000 181.610 500.000 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 496.000 185.750 500.000 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 496.000 190.350 500.000 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 496.000 74.890 500.000 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 496.000 194.490 500.000 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 496.000 198.630 500.000 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 496.000 79.030 500.000 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 496.000 83.170 500.000 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 496.000 87.310 500.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 496.000 91.910 500.000 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 496.000 96.050 500.000 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 496.000 100.190 500.000 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 496.000 104.790 500.000 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 500.000 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 496.000 246.010 500.000 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 496.000 250.150 500.000 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 496.000 254.290 500.000 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 496.000 258.430 500.000 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 496.000 263.030 500.000 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 496.000 267.170 500.000 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 496.000 271.310 500.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 496.000 275.910 500.000 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 496.000 280.050 500.000 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 496.000 284.190 500.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 496.000 207.370 500.000 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 496.000 288.790 500.000 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 496.000 292.930 500.000 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 496.000 297.070 500.000 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 496.000 301.210 500.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 496.000 305.810 500.000 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 496.000 309.950 500.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 496.000 314.090 500.000 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 496.000 318.690 500.000 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 496.000 322.830 500.000 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 496.000 326.970 500.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 496.000 211.510 500.000 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 496.000 331.570 500.000 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 496.000 335.710 500.000 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 496.000 339.850 500.000 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 496.000 343.990 500.000 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 496.000 348.590 500.000 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 496.000 352.730 500.000 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 496.000 356.870 500.000 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 496.000 361.470 500.000 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 496.000 365.610 500.000 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 496.000 369.750 500.000 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 496.000 215.650 500.000 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 496.000 374.350 500.000 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 496.000 378.490 500.000 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 496.000 382.630 500.000 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 496.000 386.770 500.000 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 496.000 391.370 500.000 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 496.000 395.510 500.000 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 496.000 399.650 500.000 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 496.000 404.250 500.000 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 496.000 408.390 500.000 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 496.000 412.530 500.000 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 496.000 220.250 500.000 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 496.000 417.130 500.000 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 496.000 421.270 500.000 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 496.000 425.410 500.000 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 496.000 429.550 500.000 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 496.000 434.150 500.000 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 496.000 438.290 500.000 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 496.000 442.430 500.000 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 496.000 447.030 500.000 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 496.000 451.170 500.000 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 496.000 455.310 500.000 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 496.000 224.390 500.000 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 496.000 459.910 500.000 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 496.000 464.050 500.000 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 496.000 468.190 500.000 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 496.000 472.330 500.000 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 496.000 228.530 500.000 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 496.000 233.130 500.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 496.000 237.270 500.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 496.000 241.410 500.000 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 496.000 519.710 500.000 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 496.000 562.490 500.000 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 496.000 566.630 500.000 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 496.000 570.770 500.000 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 496.000 575.370 500.000 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 496.000 579.510 500.000 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 496.000 583.650 500.000 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 496.000 588.250 500.000 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 496.000 592.390 500.000 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 496.000 596.530 500.000 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 496.000 600.670 500.000 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 496.000 523.850 500.000 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 496.000 605.270 500.000 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 496.000 609.410 500.000 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 496.000 613.550 500.000 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 496.000 618.150 500.000 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 496.000 622.290 500.000 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 496.000 626.430 500.000 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 496.000 631.030 500.000 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 496.000 635.170 500.000 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 496.000 639.310 500.000 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 496.000 643.450 500.000 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 496.000 527.990 500.000 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 496.000 648.050 500.000 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 496.000 652.190 500.000 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 496.000 656.330 500.000 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 496.000 660.930 500.000 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 496.000 665.070 500.000 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 496.000 669.210 500.000 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 496.000 673.810 500.000 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 496.000 677.950 500.000 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 496.000 682.090 500.000 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 496.000 686.230 500.000 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 496.000 532.590 500.000 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 496.000 690.830 500.000 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 496.000 694.970 500.000 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 496.000 699.110 500.000 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 496.000 703.710 500.000 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 496.000 707.850 500.000 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 496.000 711.990 500.000 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 496.000 716.590 500.000 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 496.000 720.730 500.000 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 496.000 724.870 500.000 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 496.000 729.010 500.000 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 496.000 536.730 500.000 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 496.000 733.610 500.000 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 496.000 737.750 500.000 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 496.000 741.890 500.000 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 496.000 746.490 500.000 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 496.000 750.630 500.000 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 496.000 754.770 500.000 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 496.000 759.370 500.000 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 496.000 763.510 500.000 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 496.000 767.650 500.000 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 496.000 771.790 500.000 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 496.000 540.870 500.000 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 496.000 776.390 500.000 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 496.000 780.530 500.000 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 496.000 784.670 500.000 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 496.000 789.270 500.000 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 496.000 545.470 500.000 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 496.000 549.610 500.000 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 496.000 553.750 500.000 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 496.000 557.890 500.000 ;
    END
  END dout1[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 495.080 800.000 495.680 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 255.040 800.000 255.640 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 270.000 800.000 270.600 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 352.960 800.000 353.560 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 360.440 800.000 361.040 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 367.920 800.000 368.520 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 375.400 800.000 376.000 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 382.880 800.000 383.480 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 389.680 800.000 390.280 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 397.160 800.000 397.760 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 404.640 800.000 405.240 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 412.120 800.000 412.720 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 419.600 800.000 420.200 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 279.520 800.000 280.120 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 426.400 800.000 427.000 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 433.880 800.000 434.480 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 441.360 800.000 441.960 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 448.840 800.000 449.440 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 289.720 800.000 290.320 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.240 800.000 299.840 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 308.760 800.000 309.360 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.240 800.000 316.840 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 323.720 800.000 324.320 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 331.200 800.000 331.800 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 338.680 800.000 339.280 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 346.160 800.000 346.760 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 257.760 800.000 258.360 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 272.040 800.000 272.640 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 355.680 800.000 356.280 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 363.160 800.000 363.760 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 370.640 800.000 371.240 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 377.440 800.000 378.040 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.920 800.000 385.520 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 392.400 800.000 393.000 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 399.880 800.000 400.480 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 407.360 800.000 407.960 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 414.160 800.000 414.760 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 421.640 800.000 422.240 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 282.240 800.000 282.840 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 429.120 800.000 429.720 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 436.600 800.000 437.200 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 444.080 800.000 444.680 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 450.880 800.000 451.480 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 456.320 800.000 456.920 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 461.080 800.000 461.680 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 465.840 800.000 466.440 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 470.600 800.000 471.200 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 475.360 800.000 475.960 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 480.800 800.000 481.400 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 291.760 800.000 292.360 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 485.560 800.000 486.160 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 490.320 800.000 490.920 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 301.960 800.000 302.560 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 311.480 800.000 312.080 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 318.960 800.000 319.560 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 326.440 800.000 327.040 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 333.920 800.000 334.520 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 340.720 800.000 341.320 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 348.200 800.000 348.800 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 274.760 800.000 275.360 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 358.400 800.000 359.000 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 365.200 800.000 365.800 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 372.680 800.000 373.280 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 380.160 800.000 380.760 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 387.640 800.000 388.240 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 395.120 800.000 395.720 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 401.920 800.000 402.520 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 409.400 800.000 410.000 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 416.880 800.000 417.480 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 424.360 800.000 424.960 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 284.280 800.000 284.880 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 431.840 800.000 432.440 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 438.640 800.000 439.240 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 446.120 800.000 446.720 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 453.600 800.000 454.200 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 458.360 800.000 458.960 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 463.120 800.000 463.720 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 468.560 800.000 469.160 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 473.320 800.000 473.920 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 478.080 800.000 478.680 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 482.840 800.000 483.440 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 294.480 800.000 295.080 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 487.600 800.000 488.200 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.040 800.000 493.640 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 304.000 800.000 304.600 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 314.200 800.000 314.800 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 321.000 800.000 321.600 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 328.480 800.000 329.080 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 335.960 800.000 336.560 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 343.440 800.000 344.040 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.920 800.000 351.520 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 259.800 800.000 260.400 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 277.480 800.000 278.080 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 287.000 800.000 287.600 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 296.520 800.000 297.120 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 306.720 800.000 307.320 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 262.520 800.000 263.120 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 265.240 800.000 265.840 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 267.280 800.000 267.880 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END partID[9]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END probe_errorCode[1]
  PIN probe_errorCode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END probe_errorCode[2]
  PIN probe_errorCode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END probe_errorCode[3]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 487.120 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 0.720 800.000 1.320 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 2.760 800.000 3.360 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 496.000 6.350 500.000 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 496.000 10.490 500.000 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 496.000 14.630 500.000 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 496.000 19.230 500.000 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 496.000 23.370 500.000 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 486.965 ;
      LAYER met1 ;
        RECT 1.910 6.160 797.570 491.600 ;
      LAYER met2 ;
        RECT 2.490 495.720 5.790 498.285 ;
        RECT 6.630 495.720 9.930 498.285 ;
        RECT 10.770 495.720 14.070 498.285 ;
        RECT 14.910 495.720 18.670 498.285 ;
        RECT 19.510 495.720 22.810 498.285 ;
        RECT 23.650 495.720 26.950 498.285 ;
        RECT 27.790 495.720 31.550 498.285 ;
        RECT 32.390 495.720 35.690 498.285 ;
        RECT 36.530 495.720 39.830 498.285 ;
        RECT 40.670 495.720 43.970 498.285 ;
        RECT 44.810 495.720 48.570 498.285 ;
        RECT 49.410 495.720 52.710 498.285 ;
        RECT 53.550 495.720 56.850 498.285 ;
        RECT 57.690 495.720 61.450 498.285 ;
        RECT 62.290 495.720 65.590 498.285 ;
        RECT 66.430 495.720 69.730 498.285 ;
        RECT 70.570 495.720 74.330 498.285 ;
        RECT 75.170 495.720 78.470 498.285 ;
        RECT 79.310 495.720 82.610 498.285 ;
        RECT 83.450 495.720 86.750 498.285 ;
        RECT 87.590 495.720 91.350 498.285 ;
        RECT 92.190 495.720 95.490 498.285 ;
        RECT 96.330 495.720 99.630 498.285 ;
        RECT 100.470 495.720 104.230 498.285 ;
        RECT 105.070 495.720 108.370 498.285 ;
        RECT 109.210 495.720 112.510 498.285 ;
        RECT 113.350 495.720 117.110 498.285 ;
        RECT 117.950 495.720 121.250 498.285 ;
        RECT 122.090 495.720 125.390 498.285 ;
        RECT 126.230 495.720 129.530 498.285 ;
        RECT 130.370 495.720 134.130 498.285 ;
        RECT 134.970 495.720 138.270 498.285 ;
        RECT 139.110 495.720 142.410 498.285 ;
        RECT 143.250 495.720 147.010 498.285 ;
        RECT 147.850 495.720 151.150 498.285 ;
        RECT 151.990 495.720 155.290 498.285 ;
        RECT 156.130 495.720 159.890 498.285 ;
        RECT 160.730 495.720 164.030 498.285 ;
        RECT 164.870 495.720 168.170 498.285 ;
        RECT 169.010 495.720 172.310 498.285 ;
        RECT 173.150 495.720 176.910 498.285 ;
        RECT 177.750 495.720 181.050 498.285 ;
        RECT 181.890 495.720 185.190 498.285 ;
        RECT 186.030 495.720 189.790 498.285 ;
        RECT 190.630 495.720 193.930 498.285 ;
        RECT 194.770 495.720 198.070 498.285 ;
        RECT 198.910 495.720 202.670 498.285 ;
        RECT 203.510 495.720 206.810 498.285 ;
        RECT 207.650 495.720 210.950 498.285 ;
        RECT 211.790 495.720 215.090 498.285 ;
        RECT 215.930 495.720 219.690 498.285 ;
        RECT 220.530 495.720 223.830 498.285 ;
        RECT 224.670 495.720 227.970 498.285 ;
        RECT 228.810 495.720 232.570 498.285 ;
        RECT 233.410 495.720 236.710 498.285 ;
        RECT 237.550 495.720 240.850 498.285 ;
        RECT 241.690 495.720 245.450 498.285 ;
        RECT 246.290 495.720 249.590 498.285 ;
        RECT 250.430 495.720 253.730 498.285 ;
        RECT 254.570 495.720 257.870 498.285 ;
        RECT 258.710 495.720 262.470 498.285 ;
        RECT 263.310 495.720 266.610 498.285 ;
        RECT 267.450 495.720 270.750 498.285 ;
        RECT 271.590 495.720 275.350 498.285 ;
        RECT 276.190 495.720 279.490 498.285 ;
        RECT 280.330 495.720 283.630 498.285 ;
        RECT 284.470 495.720 288.230 498.285 ;
        RECT 289.070 495.720 292.370 498.285 ;
        RECT 293.210 495.720 296.510 498.285 ;
        RECT 297.350 495.720 300.650 498.285 ;
        RECT 301.490 495.720 305.250 498.285 ;
        RECT 306.090 495.720 309.390 498.285 ;
        RECT 310.230 495.720 313.530 498.285 ;
        RECT 314.370 495.720 318.130 498.285 ;
        RECT 318.970 495.720 322.270 498.285 ;
        RECT 323.110 495.720 326.410 498.285 ;
        RECT 327.250 495.720 331.010 498.285 ;
        RECT 331.850 495.720 335.150 498.285 ;
        RECT 335.990 495.720 339.290 498.285 ;
        RECT 340.130 495.720 343.430 498.285 ;
        RECT 344.270 495.720 348.030 498.285 ;
        RECT 348.870 495.720 352.170 498.285 ;
        RECT 353.010 495.720 356.310 498.285 ;
        RECT 357.150 495.720 360.910 498.285 ;
        RECT 361.750 495.720 365.050 498.285 ;
        RECT 365.890 495.720 369.190 498.285 ;
        RECT 370.030 495.720 373.790 498.285 ;
        RECT 374.630 495.720 377.930 498.285 ;
        RECT 378.770 495.720 382.070 498.285 ;
        RECT 382.910 495.720 386.210 498.285 ;
        RECT 387.050 495.720 390.810 498.285 ;
        RECT 391.650 495.720 394.950 498.285 ;
        RECT 395.790 495.720 399.090 498.285 ;
        RECT 399.930 495.720 403.690 498.285 ;
        RECT 404.530 495.720 407.830 498.285 ;
        RECT 408.670 495.720 411.970 498.285 ;
        RECT 412.810 495.720 416.570 498.285 ;
        RECT 417.410 495.720 420.710 498.285 ;
        RECT 421.550 495.720 424.850 498.285 ;
        RECT 425.690 495.720 428.990 498.285 ;
        RECT 429.830 495.720 433.590 498.285 ;
        RECT 434.430 495.720 437.730 498.285 ;
        RECT 438.570 495.720 441.870 498.285 ;
        RECT 442.710 495.720 446.470 498.285 ;
        RECT 447.310 495.720 450.610 498.285 ;
        RECT 451.450 495.720 454.750 498.285 ;
        RECT 455.590 495.720 459.350 498.285 ;
        RECT 460.190 495.720 463.490 498.285 ;
        RECT 464.330 495.720 467.630 498.285 ;
        RECT 468.470 495.720 471.770 498.285 ;
        RECT 472.610 495.720 476.370 498.285 ;
        RECT 477.210 495.720 480.510 498.285 ;
        RECT 481.350 495.720 484.650 498.285 ;
        RECT 485.490 495.720 489.250 498.285 ;
        RECT 490.090 495.720 493.390 498.285 ;
        RECT 494.230 495.720 497.530 498.285 ;
        RECT 498.370 495.720 502.130 498.285 ;
        RECT 502.970 495.720 506.270 498.285 ;
        RECT 507.110 495.720 510.410 498.285 ;
        RECT 511.250 495.720 514.550 498.285 ;
        RECT 515.390 495.720 519.150 498.285 ;
        RECT 519.990 495.720 523.290 498.285 ;
        RECT 524.130 495.720 527.430 498.285 ;
        RECT 528.270 495.720 532.030 498.285 ;
        RECT 532.870 495.720 536.170 498.285 ;
        RECT 537.010 495.720 540.310 498.285 ;
        RECT 541.150 495.720 544.910 498.285 ;
        RECT 545.750 495.720 549.050 498.285 ;
        RECT 549.890 495.720 553.190 498.285 ;
        RECT 554.030 495.720 557.330 498.285 ;
        RECT 558.170 495.720 561.930 498.285 ;
        RECT 562.770 495.720 566.070 498.285 ;
        RECT 566.910 495.720 570.210 498.285 ;
        RECT 571.050 495.720 574.810 498.285 ;
        RECT 575.650 495.720 578.950 498.285 ;
        RECT 579.790 495.720 583.090 498.285 ;
        RECT 583.930 495.720 587.690 498.285 ;
        RECT 588.530 495.720 591.830 498.285 ;
        RECT 592.670 495.720 595.970 498.285 ;
        RECT 596.810 495.720 600.110 498.285 ;
        RECT 600.950 495.720 604.710 498.285 ;
        RECT 605.550 495.720 608.850 498.285 ;
        RECT 609.690 495.720 612.990 498.285 ;
        RECT 613.830 495.720 617.590 498.285 ;
        RECT 618.430 495.720 621.730 498.285 ;
        RECT 622.570 495.720 625.870 498.285 ;
        RECT 626.710 495.720 630.470 498.285 ;
        RECT 631.310 495.720 634.610 498.285 ;
        RECT 635.450 495.720 638.750 498.285 ;
        RECT 639.590 495.720 642.890 498.285 ;
        RECT 643.730 495.720 647.490 498.285 ;
        RECT 648.330 495.720 651.630 498.285 ;
        RECT 652.470 495.720 655.770 498.285 ;
        RECT 656.610 495.720 660.370 498.285 ;
        RECT 661.210 495.720 664.510 498.285 ;
        RECT 665.350 495.720 668.650 498.285 ;
        RECT 669.490 495.720 673.250 498.285 ;
        RECT 674.090 495.720 677.390 498.285 ;
        RECT 678.230 495.720 681.530 498.285 ;
        RECT 682.370 495.720 685.670 498.285 ;
        RECT 686.510 495.720 690.270 498.285 ;
        RECT 691.110 495.720 694.410 498.285 ;
        RECT 695.250 495.720 698.550 498.285 ;
        RECT 699.390 495.720 703.150 498.285 ;
        RECT 703.990 495.720 707.290 498.285 ;
        RECT 708.130 495.720 711.430 498.285 ;
        RECT 712.270 495.720 716.030 498.285 ;
        RECT 716.870 495.720 720.170 498.285 ;
        RECT 721.010 495.720 724.310 498.285 ;
        RECT 725.150 495.720 728.450 498.285 ;
        RECT 729.290 495.720 733.050 498.285 ;
        RECT 733.890 495.720 737.190 498.285 ;
        RECT 738.030 495.720 741.330 498.285 ;
        RECT 742.170 495.720 745.930 498.285 ;
        RECT 746.770 495.720 750.070 498.285 ;
        RECT 750.910 495.720 754.210 498.285 ;
        RECT 755.050 495.720 758.810 498.285 ;
        RECT 759.650 495.720 762.950 498.285 ;
        RECT 763.790 495.720 767.090 498.285 ;
        RECT 767.930 495.720 771.230 498.285 ;
        RECT 772.070 495.720 775.830 498.285 ;
        RECT 776.670 495.720 779.970 498.285 ;
        RECT 780.810 495.720 784.110 498.285 ;
        RECT 784.950 495.720 788.710 498.285 ;
        RECT 789.550 495.720 792.850 498.285 ;
        RECT 793.690 495.720 796.990 498.285 ;
        RECT 1.940 4.280 797.540 495.720 ;
        RECT 1.940 0.835 9.470 4.280 ;
        RECT 10.310 0.835 28.790 4.280 ;
        RECT 29.630 0.835 48.110 4.280 ;
        RECT 48.950 0.835 67.890 4.280 ;
        RECT 68.730 0.835 87.210 4.280 ;
        RECT 88.050 0.835 106.990 4.280 ;
        RECT 107.830 0.835 126.310 4.280 ;
        RECT 127.150 0.835 145.630 4.280 ;
        RECT 146.470 0.835 165.410 4.280 ;
        RECT 166.250 0.835 184.730 4.280 ;
        RECT 185.570 0.835 204.510 4.280 ;
        RECT 205.350 0.835 223.830 4.280 ;
        RECT 224.670 0.835 243.150 4.280 ;
        RECT 243.990 0.835 262.930 4.280 ;
        RECT 263.770 0.835 282.250 4.280 ;
        RECT 283.090 0.835 302.030 4.280 ;
        RECT 302.870 0.835 321.350 4.280 ;
        RECT 322.190 0.835 341.130 4.280 ;
        RECT 341.970 0.835 360.450 4.280 ;
        RECT 361.290 0.835 379.770 4.280 ;
        RECT 380.610 0.835 399.550 4.280 ;
        RECT 400.390 0.835 418.870 4.280 ;
        RECT 419.710 0.835 438.650 4.280 ;
        RECT 439.490 0.835 457.970 4.280 ;
        RECT 458.810 0.835 477.290 4.280 ;
        RECT 478.130 0.835 497.070 4.280 ;
        RECT 497.910 0.835 516.390 4.280 ;
        RECT 517.230 0.835 536.170 4.280 ;
        RECT 537.010 0.835 555.490 4.280 ;
        RECT 556.330 0.835 575.270 4.280 ;
        RECT 576.110 0.835 594.590 4.280 ;
        RECT 595.430 0.835 613.910 4.280 ;
        RECT 614.750 0.835 633.690 4.280 ;
        RECT 634.530 0.835 653.010 4.280 ;
        RECT 653.850 0.835 672.790 4.280 ;
        RECT 673.630 0.835 692.110 4.280 ;
        RECT 692.950 0.835 711.430 4.280 ;
        RECT 712.270 0.835 731.210 4.280 ;
        RECT 732.050 0.835 750.530 4.280 ;
        RECT 751.370 0.835 770.310 4.280 ;
        RECT 771.150 0.835 789.630 4.280 ;
        RECT 790.470 0.835 797.540 4.280 ;
      LAYER met3 ;
        RECT 4.000 497.400 795.600 498.265 ;
        RECT 4.000 496.080 796.000 497.400 ;
        RECT 4.400 494.680 795.600 496.080 ;
        RECT 4.000 494.040 796.000 494.680 ;
        RECT 4.000 492.640 795.600 494.040 ;
        RECT 4.000 491.320 796.000 492.640 ;
        RECT 4.000 489.920 795.600 491.320 ;
        RECT 4.000 488.600 796.000 489.920 ;
        RECT 4.000 487.240 795.600 488.600 ;
        RECT 4.400 487.200 795.600 487.240 ;
        RECT 4.400 486.560 796.000 487.200 ;
        RECT 4.400 485.840 795.600 486.560 ;
        RECT 4.000 485.160 795.600 485.840 ;
        RECT 4.000 483.840 796.000 485.160 ;
        RECT 4.000 482.440 795.600 483.840 ;
        RECT 4.000 481.800 796.000 482.440 ;
        RECT 4.000 480.400 795.600 481.800 ;
        RECT 4.000 479.080 796.000 480.400 ;
        RECT 4.000 478.400 795.600 479.080 ;
        RECT 4.400 477.680 795.600 478.400 ;
        RECT 4.400 477.000 796.000 477.680 ;
        RECT 4.000 476.360 796.000 477.000 ;
        RECT 4.000 474.960 795.600 476.360 ;
        RECT 4.000 474.320 796.000 474.960 ;
        RECT 4.000 472.920 795.600 474.320 ;
        RECT 4.000 471.600 796.000 472.920 ;
        RECT 4.000 470.200 795.600 471.600 ;
        RECT 4.000 469.560 796.000 470.200 ;
        RECT 4.400 468.160 795.600 469.560 ;
        RECT 4.000 466.840 796.000 468.160 ;
        RECT 4.000 465.440 795.600 466.840 ;
        RECT 4.000 464.120 796.000 465.440 ;
        RECT 4.000 462.720 795.600 464.120 ;
        RECT 4.000 462.080 796.000 462.720 ;
        RECT 4.000 460.720 795.600 462.080 ;
        RECT 4.400 460.680 795.600 460.720 ;
        RECT 4.400 459.360 796.000 460.680 ;
        RECT 4.400 459.320 795.600 459.360 ;
        RECT 4.000 457.960 795.600 459.320 ;
        RECT 4.000 457.320 796.000 457.960 ;
        RECT 4.000 455.920 795.600 457.320 ;
        RECT 4.000 454.600 796.000 455.920 ;
        RECT 4.000 453.200 795.600 454.600 ;
        RECT 4.000 451.880 796.000 453.200 ;
        RECT 4.400 450.480 795.600 451.880 ;
        RECT 4.000 449.840 796.000 450.480 ;
        RECT 4.000 448.440 795.600 449.840 ;
        RECT 4.000 447.120 796.000 448.440 ;
        RECT 4.000 445.720 795.600 447.120 ;
        RECT 4.000 445.080 796.000 445.720 ;
        RECT 4.000 443.680 795.600 445.080 ;
        RECT 4.000 443.040 796.000 443.680 ;
        RECT 4.400 442.360 796.000 443.040 ;
        RECT 4.400 441.640 795.600 442.360 ;
        RECT 4.000 440.960 795.600 441.640 ;
        RECT 4.000 439.640 796.000 440.960 ;
        RECT 4.000 438.240 795.600 439.640 ;
        RECT 4.000 437.600 796.000 438.240 ;
        RECT 4.000 436.200 795.600 437.600 ;
        RECT 4.000 434.880 796.000 436.200 ;
        RECT 4.000 434.200 795.600 434.880 ;
        RECT 4.400 433.480 795.600 434.200 ;
        RECT 4.400 432.840 796.000 433.480 ;
        RECT 4.400 432.800 795.600 432.840 ;
        RECT 4.000 431.440 795.600 432.800 ;
        RECT 4.000 430.120 796.000 431.440 ;
        RECT 4.000 428.720 795.600 430.120 ;
        RECT 4.000 427.400 796.000 428.720 ;
        RECT 4.000 426.000 795.600 427.400 ;
        RECT 4.000 425.360 796.000 426.000 ;
        RECT 4.400 423.960 795.600 425.360 ;
        RECT 4.000 422.640 796.000 423.960 ;
        RECT 4.000 421.240 795.600 422.640 ;
        RECT 4.000 420.600 796.000 421.240 ;
        RECT 4.000 419.200 795.600 420.600 ;
        RECT 4.000 417.880 796.000 419.200 ;
        RECT 4.000 417.200 795.600 417.880 ;
        RECT 4.400 416.480 795.600 417.200 ;
        RECT 4.400 415.800 796.000 416.480 ;
        RECT 4.000 415.160 796.000 415.800 ;
        RECT 4.000 413.760 795.600 415.160 ;
        RECT 4.000 413.120 796.000 413.760 ;
        RECT 4.000 411.720 795.600 413.120 ;
        RECT 4.000 410.400 796.000 411.720 ;
        RECT 4.000 409.000 795.600 410.400 ;
        RECT 4.000 408.360 796.000 409.000 ;
        RECT 4.400 406.960 795.600 408.360 ;
        RECT 4.000 405.640 796.000 406.960 ;
        RECT 4.000 404.240 795.600 405.640 ;
        RECT 4.000 402.920 796.000 404.240 ;
        RECT 4.000 401.520 795.600 402.920 ;
        RECT 4.000 400.880 796.000 401.520 ;
        RECT 4.000 399.520 795.600 400.880 ;
        RECT 4.400 399.480 795.600 399.520 ;
        RECT 4.400 398.160 796.000 399.480 ;
        RECT 4.400 398.120 795.600 398.160 ;
        RECT 4.000 396.760 795.600 398.120 ;
        RECT 4.000 396.120 796.000 396.760 ;
        RECT 4.000 394.720 795.600 396.120 ;
        RECT 4.000 393.400 796.000 394.720 ;
        RECT 4.000 392.000 795.600 393.400 ;
        RECT 4.000 390.680 796.000 392.000 ;
        RECT 4.400 389.280 795.600 390.680 ;
        RECT 4.000 388.640 796.000 389.280 ;
        RECT 4.000 387.240 795.600 388.640 ;
        RECT 4.000 385.920 796.000 387.240 ;
        RECT 4.000 384.520 795.600 385.920 ;
        RECT 4.000 383.880 796.000 384.520 ;
        RECT 4.000 382.480 795.600 383.880 ;
        RECT 4.000 381.840 796.000 382.480 ;
        RECT 4.400 381.160 796.000 381.840 ;
        RECT 4.400 380.440 795.600 381.160 ;
        RECT 4.000 379.760 795.600 380.440 ;
        RECT 4.000 378.440 796.000 379.760 ;
        RECT 4.000 377.040 795.600 378.440 ;
        RECT 4.000 376.400 796.000 377.040 ;
        RECT 4.000 375.000 795.600 376.400 ;
        RECT 4.000 373.680 796.000 375.000 ;
        RECT 4.000 373.000 795.600 373.680 ;
        RECT 4.400 372.280 795.600 373.000 ;
        RECT 4.400 371.640 796.000 372.280 ;
        RECT 4.400 371.600 795.600 371.640 ;
        RECT 4.000 370.240 795.600 371.600 ;
        RECT 4.000 368.920 796.000 370.240 ;
        RECT 4.000 367.520 795.600 368.920 ;
        RECT 4.000 366.200 796.000 367.520 ;
        RECT 4.000 364.800 795.600 366.200 ;
        RECT 4.000 364.160 796.000 364.800 ;
        RECT 4.400 362.760 795.600 364.160 ;
        RECT 4.000 361.440 796.000 362.760 ;
        RECT 4.000 360.040 795.600 361.440 ;
        RECT 4.000 359.400 796.000 360.040 ;
        RECT 4.000 358.000 795.600 359.400 ;
        RECT 4.000 356.680 796.000 358.000 ;
        RECT 4.000 355.320 795.600 356.680 ;
        RECT 4.400 355.280 795.600 355.320 ;
        RECT 4.400 353.960 796.000 355.280 ;
        RECT 4.400 353.920 795.600 353.960 ;
        RECT 4.000 352.560 795.600 353.920 ;
        RECT 4.000 351.920 796.000 352.560 ;
        RECT 4.000 350.520 795.600 351.920 ;
        RECT 4.000 349.200 796.000 350.520 ;
        RECT 4.000 347.800 795.600 349.200 ;
        RECT 4.000 347.160 796.000 347.800 ;
        RECT 4.000 346.480 795.600 347.160 ;
        RECT 4.400 345.760 795.600 346.480 ;
        RECT 4.400 345.080 796.000 345.760 ;
        RECT 4.000 344.440 796.000 345.080 ;
        RECT 4.000 343.040 795.600 344.440 ;
        RECT 4.000 341.720 796.000 343.040 ;
        RECT 4.000 340.320 795.600 341.720 ;
        RECT 4.000 339.680 796.000 340.320 ;
        RECT 4.000 338.320 795.600 339.680 ;
        RECT 4.400 338.280 795.600 338.320 ;
        RECT 4.400 336.960 796.000 338.280 ;
        RECT 4.400 336.920 795.600 336.960 ;
        RECT 4.000 335.560 795.600 336.920 ;
        RECT 4.000 334.920 796.000 335.560 ;
        RECT 4.000 333.520 795.600 334.920 ;
        RECT 4.000 332.200 796.000 333.520 ;
        RECT 4.000 330.800 795.600 332.200 ;
        RECT 4.000 329.480 796.000 330.800 ;
        RECT 4.400 328.080 795.600 329.480 ;
        RECT 4.000 327.440 796.000 328.080 ;
        RECT 4.000 326.040 795.600 327.440 ;
        RECT 4.000 324.720 796.000 326.040 ;
        RECT 4.000 323.320 795.600 324.720 ;
        RECT 4.000 322.000 796.000 323.320 ;
        RECT 4.000 320.640 795.600 322.000 ;
        RECT 4.400 320.600 795.600 320.640 ;
        RECT 4.400 319.960 796.000 320.600 ;
        RECT 4.400 319.240 795.600 319.960 ;
        RECT 4.000 318.560 795.600 319.240 ;
        RECT 4.000 317.240 796.000 318.560 ;
        RECT 4.000 315.840 795.600 317.240 ;
        RECT 4.000 315.200 796.000 315.840 ;
        RECT 4.000 313.800 795.600 315.200 ;
        RECT 4.000 312.480 796.000 313.800 ;
        RECT 4.000 311.800 795.600 312.480 ;
        RECT 4.400 311.080 795.600 311.800 ;
        RECT 4.400 310.400 796.000 311.080 ;
        RECT 4.000 309.760 796.000 310.400 ;
        RECT 4.000 308.360 795.600 309.760 ;
        RECT 4.000 307.720 796.000 308.360 ;
        RECT 4.000 306.320 795.600 307.720 ;
        RECT 4.000 305.000 796.000 306.320 ;
        RECT 4.000 303.600 795.600 305.000 ;
        RECT 4.000 302.960 796.000 303.600 ;
        RECT 4.400 301.560 795.600 302.960 ;
        RECT 4.000 300.240 796.000 301.560 ;
        RECT 4.000 298.840 795.600 300.240 ;
        RECT 4.000 297.520 796.000 298.840 ;
        RECT 4.000 296.120 795.600 297.520 ;
        RECT 4.000 295.480 796.000 296.120 ;
        RECT 4.000 294.120 795.600 295.480 ;
        RECT 4.400 294.080 795.600 294.120 ;
        RECT 4.400 292.760 796.000 294.080 ;
        RECT 4.400 292.720 795.600 292.760 ;
        RECT 4.000 291.360 795.600 292.720 ;
        RECT 4.000 290.720 796.000 291.360 ;
        RECT 4.000 289.320 795.600 290.720 ;
        RECT 4.000 288.000 796.000 289.320 ;
        RECT 4.000 286.600 795.600 288.000 ;
        RECT 4.000 285.280 796.000 286.600 ;
        RECT 4.400 283.880 795.600 285.280 ;
        RECT 4.000 283.240 796.000 283.880 ;
        RECT 4.000 281.840 795.600 283.240 ;
        RECT 4.000 280.520 796.000 281.840 ;
        RECT 4.000 279.120 795.600 280.520 ;
        RECT 4.000 278.480 796.000 279.120 ;
        RECT 4.000 277.080 795.600 278.480 ;
        RECT 4.000 276.440 796.000 277.080 ;
        RECT 4.400 275.760 796.000 276.440 ;
        RECT 4.400 275.040 795.600 275.760 ;
        RECT 4.000 274.360 795.600 275.040 ;
        RECT 4.000 273.040 796.000 274.360 ;
        RECT 4.000 271.640 795.600 273.040 ;
        RECT 4.000 271.000 796.000 271.640 ;
        RECT 4.000 269.600 795.600 271.000 ;
        RECT 4.000 268.280 796.000 269.600 ;
        RECT 4.000 267.600 795.600 268.280 ;
        RECT 4.400 266.880 795.600 267.600 ;
        RECT 4.400 266.240 796.000 266.880 ;
        RECT 4.400 266.200 795.600 266.240 ;
        RECT 4.000 264.840 795.600 266.200 ;
        RECT 4.000 263.520 796.000 264.840 ;
        RECT 4.000 262.120 795.600 263.520 ;
        RECT 4.000 260.800 796.000 262.120 ;
        RECT 4.000 259.400 795.600 260.800 ;
        RECT 4.000 258.760 796.000 259.400 ;
        RECT 4.400 257.360 795.600 258.760 ;
        RECT 4.000 256.040 796.000 257.360 ;
        RECT 4.000 254.640 795.600 256.040 ;
        RECT 4.000 254.000 796.000 254.640 ;
        RECT 4.000 252.600 795.600 254.000 ;
        RECT 4.000 251.280 796.000 252.600 ;
        RECT 4.000 250.600 795.600 251.280 ;
        RECT 4.400 249.880 795.600 250.600 ;
        RECT 4.400 249.200 796.000 249.880 ;
        RECT 4.000 248.560 796.000 249.200 ;
        RECT 4.000 247.160 795.600 248.560 ;
        RECT 4.000 246.520 796.000 247.160 ;
        RECT 4.000 245.120 795.600 246.520 ;
        RECT 4.000 243.800 796.000 245.120 ;
        RECT 4.000 242.400 795.600 243.800 ;
        RECT 4.000 241.760 796.000 242.400 ;
        RECT 4.400 240.360 795.600 241.760 ;
        RECT 4.000 239.040 796.000 240.360 ;
        RECT 4.000 237.640 795.600 239.040 ;
        RECT 4.000 236.320 796.000 237.640 ;
        RECT 4.000 234.920 795.600 236.320 ;
        RECT 4.000 234.280 796.000 234.920 ;
        RECT 4.000 232.920 795.600 234.280 ;
        RECT 4.400 232.880 795.600 232.920 ;
        RECT 4.400 231.560 796.000 232.880 ;
        RECT 4.400 231.520 795.600 231.560 ;
        RECT 4.000 230.160 795.600 231.520 ;
        RECT 4.000 229.520 796.000 230.160 ;
        RECT 4.000 228.120 795.600 229.520 ;
        RECT 4.000 226.800 796.000 228.120 ;
        RECT 4.000 225.400 795.600 226.800 ;
        RECT 4.000 224.080 796.000 225.400 ;
        RECT 4.400 222.680 795.600 224.080 ;
        RECT 4.000 222.040 796.000 222.680 ;
        RECT 4.000 220.640 795.600 222.040 ;
        RECT 4.000 219.320 796.000 220.640 ;
        RECT 4.000 217.920 795.600 219.320 ;
        RECT 4.000 217.280 796.000 217.920 ;
        RECT 4.000 215.880 795.600 217.280 ;
        RECT 4.000 215.240 796.000 215.880 ;
        RECT 4.400 214.560 796.000 215.240 ;
        RECT 4.400 213.840 795.600 214.560 ;
        RECT 4.000 213.160 795.600 213.840 ;
        RECT 4.000 211.840 796.000 213.160 ;
        RECT 4.000 210.440 795.600 211.840 ;
        RECT 4.000 209.800 796.000 210.440 ;
        RECT 4.000 208.400 795.600 209.800 ;
        RECT 4.000 207.080 796.000 208.400 ;
        RECT 4.000 206.400 795.600 207.080 ;
        RECT 4.400 205.680 795.600 206.400 ;
        RECT 4.400 205.040 796.000 205.680 ;
        RECT 4.400 205.000 795.600 205.040 ;
        RECT 4.000 203.640 795.600 205.000 ;
        RECT 4.000 202.320 796.000 203.640 ;
        RECT 4.000 200.920 795.600 202.320 ;
        RECT 4.000 199.600 796.000 200.920 ;
        RECT 4.000 198.200 795.600 199.600 ;
        RECT 4.000 197.560 796.000 198.200 ;
        RECT 4.400 196.160 795.600 197.560 ;
        RECT 4.000 194.840 796.000 196.160 ;
        RECT 4.000 193.440 795.600 194.840 ;
        RECT 4.000 192.800 796.000 193.440 ;
        RECT 4.000 191.400 795.600 192.800 ;
        RECT 4.000 190.080 796.000 191.400 ;
        RECT 4.000 188.720 795.600 190.080 ;
        RECT 4.400 188.680 795.600 188.720 ;
        RECT 4.400 187.360 796.000 188.680 ;
        RECT 4.400 187.320 795.600 187.360 ;
        RECT 4.000 185.960 795.600 187.320 ;
        RECT 4.000 185.320 796.000 185.960 ;
        RECT 4.000 183.920 795.600 185.320 ;
        RECT 4.000 182.600 796.000 183.920 ;
        RECT 4.000 181.200 795.600 182.600 ;
        RECT 4.000 180.560 796.000 181.200 ;
        RECT 4.000 179.880 795.600 180.560 ;
        RECT 4.400 179.160 795.600 179.880 ;
        RECT 4.400 178.480 796.000 179.160 ;
        RECT 4.000 177.840 796.000 178.480 ;
        RECT 4.000 176.440 795.600 177.840 ;
        RECT 4.000 175.120 796.000 176.440 ;
        RECT 4.000 173.720 795.600 175.120 ;
        RECT 4.000 173.080 796.000 173.720 ;
        RECT 4.000 171.720 795.600 173.080 ;
        RECT 4.400 171.680 795.600 171.720 ;
        RECT 4.400 170.360 796.000 171.680 ;
        RECT 4.400 170.320 795.600 170.360 ;
        RECT 4.000 168.960 795.600 170.320 ;
        RECT 4.000 168.320 796.000 168.960 ;
        RECT 4.000 166.920 795.600 168.320 ;
        RECT 4.000 165.600 796.000 166.920 ;
        RECT 4.000 164.200 795.600 165.600 ;
        RECT 4.000 162.880 796.000 164.200 ;
        RECT 4.400 161.480 795.600 162.880 ;
        RECT 4.000 160.840 796.000 161.480 ;
        RECT 4.000 159.440 795.600 160.840 ;
        RECT 4.000 158.120 796.000 159.440 ;
        RECT 4.000 156.720 795.600 158.120 ;
        RECT 4.000 155.400 796.000 156.720 ;
        RECT 4.000 154.040 795.600 155.400 ;
        RECT 4.400 154.000 795.600 154.040 ;
        RECT 4.400 153.360 796.000 154.000 ;
        RECT 4.400 152.640 795.600 153.360 ;
        RECT 4.000 151.960 795.600 152.640 ;
        RECT 4.000 150.640 796.000 151.960 ;
        RECT 4.000 149.240 795.600 150.640 ;
        RECT 4.000 148.600 796.000 149.240 ;
        RECT 4.000 147.200 795.600 148.600 ;
        RECT 4.000 145.880 796.000 147.200 ;
        RECT 4.000 145.200 795.600 145.880 ;
        RECT 4.400 144.480 795.600 145.200 ;
        RECT 4.400 143.800 796.000 144.480 ;
        RECT 4.000 143.160 796.000 143.800 ;
        RECT 4.000 141.760 795.600 143.160 ;
        RECT 4.000 141.120 796.000 141.760 ;
        RECT 4.000 139.720 795.600 141.120 ;
        RECT 4.000 138.400 796.000 139.720 ;
        RECT 4.000 137.000 795.600 138.400 ;
        RECT 4.000 136.360 796.000 137.000 ;
        RECT 4.400 134.960 795.600 136.360 ;
        RECT 4.000 133.640 796.000 134.960 ;
        RECT 4.000 132.240 795.600 133.640 ;
        RECT 4.000 130.920 796.000 132.240 ;
        RECT 4.000 129.520 795.600 130.920 ;
        RECT 4.000 128.880 796.000 129.520 ;
        RECT 4.000 127.520 795.600 128.880 ;
        RECT 4.400 127.480 795.600 127.520 ;
        RECT 4.400 126.160 796.000 127.480 ;
        RECT 4.400 126.120 795.600 126.160 ;
        RECT 4.000 124.760 795.600 126.120 ;
        RECT 4.000 124.120 796.000 124.760 ;
        RECT 4.000 122.720 795.600 124.120 ;
        RECT 4.000 121.400 796.000 122.720 ;
        RECT 4.000 120.000 795.600 121.400 ;
        RECT 4.000 118.680 796.000 120.000 ;
        RECT 4.400 117.280 795.600 118.680 ;
        RECT 4.000 116.640 796.000 117.280 ;
        RECT 4.000 115.240 795.600 116.640 ;
        RECT 4.000 113.920 796.000 115.240 ;
        RECT 4.000 112.520 795.600 113.920 ;
        RECT 4.000 111.880 796.000 112.520 ;
        RECT 4.000 110.480 795.600 111.880 ;
        RECT 4.000 109.840 796.000 110.480 ;
        RECT 4.400 109.160 796.000 109.840 ;
        RECT 4.400 108.440 795.600 109.160 ;
        RECT 4.000 107.760 795.600 108.440 ;
        RECT 4.000 106.440 796.000 107.760 ;
        RECT 4.000 105.040 795.600 106.440 ;
        RECT 4.000 104.400 796.000 105.040 ;
        RECT 4.000 103.000 795.600 104.400 ;
        RECT 4.000 101.680 796.000 103.000 ;
        RECT 4.000 101.000 795.600 101.680 ;
        RECT 4.400 100.280 795.600 101.000 ;
        RECT 4.400 99.640 796.000 100.280 ;
        RECT 4.400 99.600 795.600 99.640 ;
        RECT 4.000 98.240 795.600 99.600 ;
        RECT 4.000 96.920 796.000 98.240 ;
        RECT 4.000 95.520 795.600 96.920 ;
        RECT 4.000 94.200 796.000 95.520 ;
        RECT 4.000 92.800 795.600 94.200 ;
        RECT 4.000 92.160 796.000 92.800 ;
        RECT 4.400 90.760 795.600 92.160 ;
        RECT 4.000 89.440 796.000 90.760 ;
        RECT 4.000 88.040 795.600 89.440 ;
        RECT 4.000 87.400 796.000 88.040 ;
        RECT 4.000 86.000 795.600 87.400 ;
        RECT 4.000 84.680 796.000 86.000 ;
        RECT 4.000 84.000 795.600 84.680 ;
        RECT 4.400 83.280 795.600 84.000 ;
        RECT 4.400 82.600 796.000 83.280 ;
        RECT 4.000 81.960 796.000 82.600 ;
        RECT 4.000 80.560 795.600 81.960 ;
        RECT 4.000 79.920 796.000 80.560 ;
        RECT 4.000 78.520 795.600 79.920 ;
        RECT 4.000 77.200 796.000 78.520 ;
        RECT 4.000 75.800 795.600 77.200 ;
        RECT 4.000 75.160 796.000 75.800 ;
        RECT 4.400 73.760 795.600 75.160 ;
        RECT 4.000 72.440 796.000 73.760 ;
        RECT 4.000 71.040 795.600 72.440 ;
        RECT 4.000 69.720 796.000 71.040 ;
        RECT 4.000 68.320 795.600 69.720 ;
        RECT 4.000 67.680 796.000 68.320 ;
        RECT 4.000 66.320 795.600 67.680 ;
        RECT 4.400 66.280 795.600 66.320 ;
        RECT 4.400 64.960 796.000 66.280 ;
        RECT 4.400 64.920 795.600 64.960 ;
        RECT 4.000 63.560 795.600 64.920 ;
        RECT 4.000 62.920 796.000 63.560 ;
        RECT 4.000 61.520 795.600 62.920 ;
        RECT 4.000 60.200 796.000 61.520 ;
        RECT 4.000 58.800 795.600 60.200 ;
        RECT 4.000 57.480 796.000 58.800 ;
        RECT 4.400 56.080 795.600 57.480 ;
        RECT 4.000 55.440 796.000 56.080 ;
        RECT 4.000 54.040 795.600 55.440 ;
        RECT 4.000 52.720 796.000 54.040 ;
        RECT 4.000 51.320 795.600 52.720 ;
        RECT 4.000 50.680 796.000 51.320 ;
        RECT 4.000 49.280 795.600 50.680 ;
        RECT 4.000 48.640 796.000 49.280 ;
        RECT 4.400 47.960 796.000 48.640 ;
        RECT 4.400 47.240 795.600 47.960 ;
        RECT 4.000 46.560 795.600 47.240 ;
        RECT 4.000 45.240 796.000 46.560 ;
        RECT 4.000 43.840 795.600 45.240 ;
        RECT 4.000 43.200 796.000 43.840 ;
        RECT 4.000 41.800 795.600 43.200 ;
        RECT 4.000 40.480 796.000 41.800 ;
        RECT 4.000 39.800 795.600 40.480 ;
        RECT 4.400 39.080 795.600 39.800 ;
        RECT 4.400 38.440 796.000 39.080 ;
        RECT 4.400 38.400 795.600 38.440 ;
        RECT 4.000 37.040 795.600 38.400 ;
        RECT 4.000 35.720 796.000 37.040 ;
        RECT 4.000 34.320 795.600 35.720 ;
        RECT 4.000 33.000 796.000 34.320 ;
        RECT 4.000 31.600 795.600 33.000 ;
        RECT 4.000 30.960 796.000 31.600 ;
        RECT 4.400 29.560 795.600 30.960 ;
        RECT 4.000 28.240 796.000 29.560 ;
        RECT 4.000 26.840 795.600 28.240 ;
        RECT 4.000 26.200 796.000 26.840 ;
        RECT 4.000 24.800 795.600 26.200 ;
        RECT 4.000 23.480 796.000 24.800 ;
        RECT 4.000 22.120 795.600 23.480 ;
        RECT 4.400 22.080 795.600 22.120 ;
        RECT 4.400 20.760 796.000 22.080 ;
        RECT 4.400 20.720 795.600 20.760 ;
        RECT 4.000 19.360 795.600 20.720 ;
        RECT 4.000 18.720 796.000 19.360 ;
        RECT 4.000 17.320 795.600 18.720 ;
        RECT 4.000 16.000 796.000 17.320 ;
        RECT 4.000 14.600 795.600 16.000 ;
        RECT 4.000 13.960 796.000 14.600 ;
        RECT 4.000 13.280 795.600 13.960 ;
        RECT 4.400 12.560 795.600 13.280 ;
        RECT 4.400 11.880 796.000 12.560 ;
        RECT 4.000 11.240 796.000 11.880 ;
        RECT 4.000 9.840 795.600 11.240 ;
        RECT 4.000 8.520 796.000 9.840 ;
        RECT 4.000 7.120 795.600 8.520 ;
        RECT 4.000 6.480 796.000 7.120 ;
        RECT 4.000 5.120 795.600 6.480 ;
        RECT 4.400 5.080 795.600 5.120 ;
        RECT 4.400 3.760 796.000 5.080 ;
        RECT 4.400 3.720 795.600 3.760 ;
        RECT 4.000 2.360 795.600 3.720 ;
        RECT 4.000 1.720 796.000 2.360 ;
        RECT 4.000 0.855 795.600 1.720 ;
      LAYER met4 ;
        RECT 781.375 285.095 785.385 471.745 ;
  END
END ExperiarCore
END LIBRARY

