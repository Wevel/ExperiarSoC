magic
tech sky130A
magscale 1 2
timestamp 1651190804
<< viali >>
rect 38025 37417 38059 37451
rect 16773 37281 16807 37315
rect 22293 37213 22327 37247
rect 30021 37213 30055 37247
rect 37841 37213 37875 37247
rect 30205 37077 30239 37111
rect 37381 37077 37415 37111
rect 29929 36873 29963 36907
rect 13369 36805 13403 36839
rect 22201 36737 22235 36771
rect 2697 36669 2731 36703
rect 2881 36669 2915 36703
rect 4169 36669 4203 36703
rect 13185 36669 13219 36703
rect 13829 36669 13863 36703
rect 22385 36669 22419 36703
rect 22661 36669 22695 36703
rect 4997 36533 5031 36567
rect 9045 36533 9079 36567
rect 17417 36533 17451 36567
rect 25513 36533 25547 36567
rect 2329 36329 2363 36363
rect 12909 36329 12943 36363
rect 5273 36193 5307 36227
rect 9413 36193 9447 36227
rect 13553 36193 13587 36227
rect 15945 36193 15979 36227
rect 18705 36193 18739 36227
rect 22109 36193 22143 36227
rect 24409 36193 24443 36227
rect 25421 36193 25455 36227
rect 2789 36125 2823 36159
rect 4353 36125 4387 36159
rect 4813 36125 4847 36159
rect 8401 36125 8435 36159
rect 8953 36125 8987 36159
rect 12081 36125 12115 36159
rect 21189 36125 21223 36159
rect 21649 36125 21683 36159
rect 30941 36125 30975 36159
rect 4997 36057 5031 36091
rect 9137 36057 9171 36091
rect 14105 36057 14139 36091
rect 15761 36057 15795 36091
rect 16865 36057 16899 36091
rect 18521 36057 18555 36091
rect 21833 36057 21867 36091
rect 25605 36057 25639 36091
rect 27261 36057 27295 36091
rect 30674 36057 30708 36091
rect 29561 35989 29595 36023
rect 4997 35785 5031 35819
rect 21833 35785 21867 35819
rect 29745 35785 29779 35819
rect 2697 35649 2731 35683
rect 5181 35649 5215 35683
rect 13645 35649 13679 35683
rect 16773 35649 16807 35683
rect 19349 35649 19383 35683
rect 22017 35649 22051 35683
rect 22477 35649 22511 35683
rect 23489 35649 23523 35683
rect 28834 35649 28868 35683
rect 29561 35649 29595 35683
rect 2881 35581 2915 35615
rect 3157 35581 3191 35615
rect 7297 35581 7331 35615
rect 7481 35581 7515 35615
rect 9137 35581 9171 35615
rect 11805 35581 11839 35615
rect 13461 35581 13495 35615
rect 16957 35581 16991 35615
rect 17233 35581 17267 35615
rect 19073 35581 19107 35615
rect 23673 35581 23707 35615
rect 23949 35581 23983 35615
rect 29101 35581 29135 35615
rect 22661 35513 22695 35547
rect 10977 35445 11011 35479
rect 15485 35445 15519 35479
rect 25973 35445 26007 35479
rect 27721 35445 27755 35479
rect 7389 35241 7423 35275
rect 19441 35241 19475 35275
rect 19625 35241 19659 35275
rect 20545 35241 20579 35275
rect 21281 35241 21315 35275
rect 21741 35241 21775 35275
rect 22385 35241 22419 35275
rect 28457 35241 28491 35275
rect 20361 35173 20395 35207
rect 2973 35105 3007 35139
rect 4629 35105 4663 35139
rect 5549 35105 5583 35139
rect 8953 35105 8987 35139
rect 9413 35105 9447 35139
rect 11805 35105 11839 35139
rect 13553 35105 13587 35139
rect 14381 35105 14415 35139
rect 15485 35105 15519 35139
rect 16865 35105 16899 35139
rect 18429 35105 18463 35139
rect 18705 35105 18739 35139
rect 19809 35105 19843 35139
rect 20637 35105 20671 35139
rect 21373 35105 21407 35139
rect 26249 35105 26283 35139
rect 3249 35037 3283 35071
rect 3985 35037 4019 35071
rect 14105 35037 14139 35071
rect 19625 35037 19659 35071
rect 20545 35037 20579 35071
rect 21557 35037 21591 35071
rect 22201 35037 22235 35071
rect 28273 35037 28307 35071
rect 4813 34969 4847 35003
rect 9137 34969 9171 35003
rect 13369 34969 13403 35003
rect 15669 34969 15703 35003
rect 19901 34969 19935 35003
rect 20821 34969 20855 35003
rect 21281 34969 21315 35003
rect 24409 34969 24443 35003
rect 26065 34969 26099 35003
rect 4169 34901 4203 34935
rect 4721 34697 4755 34731
rect 7573 34697 7607 34731
rect 8585 34697 8619 34731
rect 15577 34697 15611 34731
rect 17601 34697 17635 34731
rect 21189 34697 21223 34731
rect 28365 34697 28399 34731
rect 29653 34697 29687 34731
rect 10885 34629 10919 34663
rect 18245 34629 18279 34663
rect 3985 34561 4019 34595
rect 4905 34561 4939 34595
rect 5181 34561 5215 34595
rect 7389 34561 7423 34595
rect 8401 34561 8435 34595
rect 13277 34561 13311 34595
rect 14565 34561 14599 34595
rect 15393 34561 15427 34595
rect 17417 34561 17451 34595
rect 20729 34561 20763 34595
rect 21005 34561 21039 34595
rect 23857 34561 23891 34595
rect 25145 34561 25179 34595
rect 28549 34561 28583 34595
rect 29469 34561 29503 34595
rect 31309 34561 31343 34595
rect 31493 34561 31527 34595
rect 32137 34561 32171 34595
rect 4261 34493 4295 34527
rect 4997 34493 5031 34527
rect 9045 34493 9079 34527
rect 9229 34493 9263 34527
rect 13553 34493 13587 34527
rect 14841 34493 14875 34527
rect 18061 34493 18095 34527
rect 18521 34493 18555 34527
rect 20821 34493 20855 34527
rect 23581 34493 23615 34527
rect 24869 34493 24903 34527
rect 28733 34493 28767 34527
rect 29285 34493 29319 34527
rect 31125 34493 31159 34527
rect 4905 34357 4939 34391
rect 5733 34357 5767 34391
rect 20729 34357 20763 34391
rect 32321 34357 32355 34391
rect 4721 34153 4755 34187
rect 4905 34153 4939 34187
rect 5549 34153 5583 34187
rect 9137 34153 9171 34187
rect 9597 34153 9631 34187
rect 15669 34153 15703 34187
rect 16129 34153 16163 34187
rect 18429 34153 18463 34187
rect 5365 34085 5399 34119
rect 18613 34085 18647 34119
rect 5641 34017 5675 34051
rect 16037 34017 16071 34051
rect 26341 34017 26375 34051
rect 32597 34017 32631 34051
rect 1409 33949 1443 33983
rect 2513 33949 2547 33983
rect 3985 33949 4019 33983
rect 4629 33949 4663 33983
rect 4721 33949 4755 33983
rect 5549 33949 5583 33983
rect 8953 33949 8987 33983
rect 9781 33949 9815 33983
rect 12725 33949 12759 33983
rect 15853 33949 15887 33983
rect 18337 33949 18371 33983
rect 18429 33949 18463 33983
rect 25421 33949 25455 33983
rect 32330 33949 32364 33983
rect 37473 33949 37507 33983
rect 38117 33949 38151 33983
rect 4445 33881 4479 33915
rect 5825 33881 5859 33915
rect 16129 33881 16163 33915
rect 18153 33881 18187 33915
rect 25605 33881 25639 33915
rect 29009 33881 29043 33915
rect 1593 33813 1627 33847
rect 3801 33813 3835 33847
rect 6377 33813 6411 33847
rect 29653 33813 29687 33847
rect 30481 33813 30515 33847
rect 31217 33813 31251 33847
rect 37933 33813 37967 33847
rect 4721 33609 4755 33643
rect 5733 33609 5767 33643
rect 23121 33609 23155 33643
rect 28273 33609 28307 33643
rect 29285 33609 29319 33643
rect 31309 33609 31343 33643
rect 1409 33541 1443 33575
rect 2605 33541 2639 33575
rect 14105 33541 14139 33575
rect 22661 33541 22695 33575
rect 28641 33541 28675 33575
rect 29561 33541 29595 33575
rect 29653 33541 29687 33575
rect 30941 33541 30975 33575
rect 31033 33541 31067 33575
rect 2421 33473 2455 33507
rect 4905 33473 4939 33507
rect 5181 33473 5215 33507
rect 9045 33473 9079 33507
rect 14289 33473 14323 33507
rect 15301 33473 15335 33507
rect 18153 33473 18187 33507
rect 20361 33473 20395 33507
rect 22937 33473 22971 33507
rect 25421 33473 25455 33507
rect 28457 33473 28491 33507
rect 28549 33473 28583 33507
rect 28825 33473 28859 33507
rect 29469 33473 29503 33507
rect 29837 33473 29871 33507
rect 30757 33473 30791 33507
rect 31125 33473 31159 33507
rect 2881 33405 2915 33439
rect 5089 33405 5123 33439
rect 12449 33405 12483 33439
rect 15577 33405 15611 33439
rect 20637 33405 20671 33439
rect 22753 33405 22787 33439
rect 5181 33269 5215 33303
rect 22845 33269 22879 33303
rect 27813 33269 27847 33303
rect 4077 33065 4111 33099
rect 4537 33065 4571 33099
rect 8125 33065 8159 33099
rect 8401 33065 8435 33099
rect 8953 33065 8987 33099
rect 9137 33065 9171 33099
rect 16129 33065 16163 33099
rect 16589 33065 16623 33099
rect 16773 33065 16807 33099
rect 19993 33065 20027 33099
rect 20637 33065 20671 33099
rect 21925 33065 21959 33099
rect 22109 33065 22143 33099
rect 22569 33065 22603 33099
rect 23029 33065 23063 33099
rect 15669 32997 15703 33031
rect 4445 32929 4479 32963
rect 8125 32929 8159 32963
rect 9321 32929 9355 32963
rect 14933 32929 14967 32963
rect 16037 32929 16071 32963
rect 16957 32929 16991 32963
rect 21741 32929 21775 32963
rect 22661 32929 22695 32963
rect 27169 32929 27203 32963
rect 28365 32929 28399 32963
rect 4261 32861 4295 32895
rect 5641 32861 5675 32895
rect 8217 32861 8251 32895
rect 9137 32861 9171 32895
rect 12725 32861 12759 32895
rect 14657 32861 14691 32895
rect 15853 32861 15887 32895
rect 16129 32861 16163 32895
rect 16773 32861 16807 32895
rect 19809 32861 19843 32895
rect 20453 32861 20487 32895
rect 21925 32861 21959 32895
rect 22845 32861 22879 32895
rect 24869 32861 24903 32895
rect 4537 32793 4571 32827
rect 7941 32793 7975 32827
rect 9413 32793 9447 32827
rect 17049 32793 17083 32827
rect 21649 32793 21683 32827
rect 22569 32793 22603 32827
rect 25053 32793 25087 32827
rect 26709 32793 26743 32827
rect 27353 32793 27387 32827
rect 30021 32793 30055 32827
rect 30665 32725 30699 32759
rect 5365 32521 5399 32555
rect 7389 32521 7423 32555
rect 8677 32521 8711 32555
rect 17141 32521 17175 32555
rect 18337 32521 18371 32555
rect 20729 32521 20763 32555
rect 22017 32521 22051 32555
rect 23489 32521 23523 32555
rect 25329 32521 25363 32555
rect 6929 32453 6963 32487
rect 8217 32453 8251 32487
rect 14105 32453 14139 32487
rect 1409 32385 1443 32419
rect 2053 32385 2087 32419
rect 4721 32385 4755 32419
rect 5181 32385 5215 32419
rect 7205 32385 7239 32419
rect 8493 32385 8527 32419
rect 14289 32385 14323 32419
rect 16957 32385 16991 32419
rect 17601 32385 17635 32419
rect 18521 32385 18555 32419
rect 19165 32385 19199 32419
rect 19809 32385 19843 32419
rect 20545 32385 20579 32419
rect 21189 32385 21223 32419
rect 22201 32385 22235 32419
rect 23029 32385 23063 32419
rect 23305 32385 23339 32419
rect 24685 32385 24719 32419
rect 25513 32385 25547 32419
rect 25973 32385 26007 32419
rect 28457 32385 28491 32419
rect 32321 32385 32355 32419
rect 33057 32385 33091 32419
rect 33324 32385 33358 32419
rect 7021 32317 7055 32351
rect 8401 32317 8435 32351
rect 12725 32317 12759 32351
rect 15301 32317 15335 32351
rect 15577 32317 15611 32351
rect 23213 32317 23247 32351
rect 28641 32317 28675 32351
rect 29009 32317 29043 32351
rect 32137 32317 32171 32351
rect 24869 32249 24903 32283
rect 1593 32181 1627 32215
rect 7205 32181 7239 32215
rect 8217 32181 8251 32215
rect 18981 32181 19015 32215
rect 19625 32181 19659 32215
rect 23305 32181 23339 32215
rect 23949 32181 23983 32215
rect 32505 32181 32539 32215
rect 34437 32181 34471 32215
rect 4997 31977 5031 32011
rect 15761 31977 15795 32011
rect 16221 31977 16255 32011
rect 19625 31977 19659 32011
rect 22109 31977 22143 32011
rect 33241 31977 33275 32011
rect 21005 31909 21039 31943
rect 5641 31841 5675 31875
rect 6101 31841 6135 31875
rect 12449 31841 12483 31875
rect 13369 31841 13403 31875
rect 16037 31841 16071 31875
rect 19625 31841 19659 31875
rect 30757 31841 30791 31875
rect 30941 31841 30975 31875
rect 31585 31841 31619 31875
rect 5181 31773 5215 31807
rect 13553 31773 13587 31807
rect 14289 31773 14323 31807
rect 15945 31773 15979 31807
rect 16221 31773 16255 31807
rect 19441 31773 19475 31807
rect 19717 31773 19751 31807
rect 20545 31773 20579 31807
rect 22293 31773 22327 31807
rect 22753 31773 22787 31807
rect 23029 31773 23063 31807
rect 33057 31773 33091 31807
rect 5825 31705 5859 31739
rect 19257 31637 19291 31671
rect 20361 31637 20395 31671
rect 5549 31433 5583 31467
rect 6377 31433 6411 31467
rect 19901 31433 19935 31467
rect 24317 31433 24351 31467
rect 32689 31433 32723 31467
rect 35081 31433 35115 31467
rect 2513 31365 2547 31399
rect 7297 31365 7331 31399
rect 14749 31365 14783 31399
rect 21833 31365 21867 31399
rect 32321 31365 32355 31399
rect 35173 31365 35207 31399
rect 1409 31297 1443 31331
rect 2789 31297 2823 31331
rect 5733 31297 5767 31331
rect 6561 31297 6595 31331
rect 7481 31297 7515 31331
rect 8033 31297 8067 31331
rect 12357 31297 12391 31331
rect 14933 31297 14967 31331
rect 22017 31297 22051 31331
rect 22569 31297 22603 31331
rect 22845 31297 22879 31331
rect 23857 31297 23891 31331
rect 24133 31297 24167 31331
rect 27261 31297 27295 31331
rect 30113 31297 30147 31331
rect 32137 31297 32171 31331
rect 32413 31297 32447 31331
rect 32505 31297 32539 31331
rect 2605 31229 2639 31263
rect 13093 31229 13127 31263
rect 24041 31229 24075 31263
rect 26985 31229 27019 31263
rect 29837 31229 29871 31263
rect 34897 31229 34931 31263
rect 1593 31161 1627 31195
rect 34253 31161 34287 31195
rect 2513 31093 2547 31127
rect 2973 31093 3007 31127
rect 8953 31093 8987 31127
rect 21281 31093 21315 31127
rect 23857 31093 23891 31127
rect 24777 31093 24811 31127
rect 31493 31093 31527 31127
rect 35541 31093 35575 31127
rect 6193 30889 6227 30923
rect 6377 30889 6411 30923
rect 21097 30889 21131 30923
rect 21925 30889 21959 30923
rect 25605 30889 25639 30923
rect 32045 30889 32079 30923
rect 1409 30821 1443 30855
rect 22109 30821 22143 30855
rect 22845 30821 22879 30855
rect 26065 30821 26099 30855
rect 6101 30753 6135 30787
rect 8953 30753 8987 30787
rect 21741 30753 21775 30787
rect 25697 30753 25731 30787
rect 27353 30753 27387 30787
rect 27629 30753 27663 30787
rect 31401 30753 31435 30787
rect 2789 30685 2823 30719
rect 6193 30685 6227 30719
rect 12909 30685 12943 30719
rect 17693 30685 17727 30719
rect 18705 30685 18739 30719
rect 21925 30685 21959 30719
rect 25881 30685 25915 30719
rect 5917 30617 5951 30651
rect 9137 30617 9171 30651
rect 10793 30617 10827 30651
rect 21649 30617 21683 30651
rect 22661 30617 22695 30651
rect 23305 30617 23339 30651
rect 25605 30617 25639 30651
rect 29561 30617 29595 30651
rect 31217 30617 31251 30651
rect 18521 30549 18555 30583
rect 5089 30345 5123 30379
rect 17785 30277 17819 30311
rect 25513 30277 25547 30311
rect 26985 30277 27019 30311
rect 31401 30277 31435 30311
rect 2789 30209 2823 30243
rect 5273 30209 5307 30243
rect 5733 30209 5767 30243
rect 14473 30209 14507 30243
rect 17601 30209 17635 30243
rect 21833 30209 21867 30243
rect 25789 30209 25823 30243
rect 27261 30209 27295 30243
rect 28549 30209 28583 30243
rect 29745 30209 29779 30243
rect 33793 30209 33827 30243
rect 34060 30209 34094 30243
rect 2973 30141 3007 30175
rect 3249 30141 3283 30175
rect 7021 30141 7055 30175
rect 7297 30141 7331 30175
rect 7757 30141 7791 30175
rect 8493 30141 8527 30175
rect 8953 30141 8987 30175
rect 9137 30141 9171 30175
rect 9413 30141 9447 30175
rect 13093 30141 13127 30175
rect 14289 30141 14323 30175
rect 18245 30141 18279 30175
rect 22109 30141 22143 30175
rect 25605 30141 25639 30175
rect 27077 30141 27111 30175
rect 28273 30141 28307 30175
rect 30021 30141 30055 30175
rect 25973 30073 26007 30107
rect 27445 30073 27479 30107
rect 2329 30005 2363 30039
rect 16681 30005 16715 30039
rect 20913 30005 20947 30039
rect 25053 30005 25087 30039
rect 25513 30005 25547 30039
rect 26985 30005 27019 30039
rect 35173 30005 35207 30039
rect 38117 30005 38151 30039
rect 1593 29801 1627 29835
rect 6837 29801 6871 29835
rect 9137 29801 9171 29835
rect 14473 29801 14507 29835
rect 14933 29801 14967 29835
rect 3801 29665 3835 29699
rect 4629 29665 4663 29699
rect 13277 29665 13311 29699
rect 14841 29665 14875 29699
rect 16681 29665 16715 29699
rect 18521 29665 18555 29699
rect 20729 29665 20763 29699
rect 22293 29665 22327 29699
rect 22477 29665 22511 29699
rect 25237 29665 25271 29699
rect 26709 29665 26743 29699
rect 36369 29665 36403 29699
rect 1409 29597 1443 29631
rect 2053 29597 2087 29631
rect 3065 29597 3099 29631
rect 6653 29597 6687 29631
rect 7297 29597 7331 29631
rect 8953 29597 8987 29631
rect 9597 29597 9631 29631
rect 12265 29597 12299 29631
rect 13553 29597 13587 29631
rect 14657 29597 14691 29631
rect 19441 29597 19475 29631
rect 23121 29597 23155 29631
rect 23581 29597 23615 29631
rect 24593 29597 24627 29631
rect 3985 29529 4019 29563
rect 14933 29529 14967 29563
rect 16865 29529 16899 29563
rect 25421 29529 25455 29563
rect 36614 29529 36648 29563
rect 3249 29461 3283 29495
rect 22937 29461 22971 29495
rect 24777 29461 24811 29495
rect 35725 29461 35759 29495
rect 37749 29461 37783 29495
rect 2881 29257 2915 29291
rect 8401 29257 8435 29291
rect 15393 29257 15427 29291
rect 16865 29257 16899 29291
rect 22937 29257 22971 29291
rect 24501 29257 24535 29291
rect 29285 29257 29319 29291
rect 35173 29257 35207 29291
rect 36461 29257 36495 29291
rect 14933 29189 14967 29223
rect 22477 29189 22511 29223
rect 2697 29121 2731 29155
rect 8217 29121 8251 29155
rect 8861 29121 8895 29155
rect 12265 29121 12299 29155
rect 15209 29121 15243 29155
rect 16681 29121 16715 29155
rect 20545 29121 20579 29155
rect 21833 29121 21867 29155
rect 22753 29121 22787 29155
rect 24041 29121 24075 29155
rect 24317 29121 24351 29155
rect 29101 29121 29135 29155
rect 34989 29121 35023 29155
rect 35817 29121 35851 29155
rect 36001 29121 36035 29155
rect 36093 29121 36127 29155
rect 36185 29121 36219 29155
rect 2237 29053 2271 29087
rect 3341 29053 3375 29087
rect 3525 29053 3559 29087
rect 3893 29053 3927 29087
rect 9045 29053 9079 29087
rect 10701 29053 10735 29087
rect 12449 29053 12483 29087
rect 12725 29053 12759 29087
rect 15025 29053 15059 29087
rect 19165 29053 19199 29087
rect 20361 29053 20395 29087
rect 22569 29053 22603 29087
rect 24133 29053 24167 29087
rect 35357 29053 35391 29087
rect 22017 28985 22051 29019
rect 15209 28917 15243 28951
rect 22477 28917 22511 28951
rect 24041 28917 24075 28951
rect 34805 28917 34839 28951
rect 3249 28713 3283 28747
rect 3801 28713 3835 28747
rect 4261 28713 4295 28747
rect 7941 28713 7975 28747
rect 8401 28713 8435 28747
rect 9137 28713 9171 28747
rect 15485 28713 15519 28747
rect 28457 28713 28491 28747
rect 37197 28713 37231 28747
rect 15853 28645 15887 28679
rect 4077 28577 4111 28611
rect 8033 28577 8067 28611
rect 13277 28577 13311 28611
rect 14381 28577 14415 28611
rect 15485 28577 15519 28611
rect 18245 28577 18279 28611
rect 20177 28577 20211 28611
rect 35265 28577 35299 28611
rect 37105 28577 37139 28611
rect 1409 28509 1443 28543
rect 2053 28509 2087 28543
rect 3065 28509 3099 28543
rect 3985 28509 4019 28543
rect 4261 28509 4295 28543
rect 7941 28509 7975 28543
rect 8217 28509 8251 28543
rect 8953 28509 8987 28543
rect 13553 28509 13587 28543
rect 14105 28509 14139 28543
rect 15669 28509 15703 28543
rect 16865 28509 16899 28543
rect 20453 28509 20487 28543
rect 37289 28509 37323 28543
rect 37381 28509 37415 28543
rect 15393 28441 15427 28475
rect 17049 28441 17083 28475
rect 28089 28441 28123 28475
rect 28273 28441 28307 28475
rect 35532 28441 35566 28475
rect 1593 28373 1627 28407
rect 29009 28373 29043 28407
rect 36645 28373 36679 28407
rect 3709 28169 3743 28203
rect 8401 28169 8435 28203
rect 13737 28169 13771 28203
rect 15301 28169 15335 28203
rect 20637 28169 20671 28203
rect 21097 28169 21131 28203
rect 34069 28169 34103 28203
rect 4169 28101 4203 28135
rect 7941 28101 7975 28135
rect 9229 28101 9263 28135
rect 14197 28101 14231 28135
rect 14841 28101 14875 28135
rect 30297 28101 30331 28135
rect 31585 28101 31619 28135
rect 3893 28033 3927 28067
rect 3985 28033 4019 28067
rect 8217 28033 8251 28067
rect 13921 28033 13955 28067
rect 15117 28033 15151 28067
rect 16957 28033 16991 28067
rect 27629 28033 27663 28067
rect 27896 28033 27930 28067
rect 30481 28033 30515 28067
rect 31033 28033 31067 28067
rect 31125 28033 31159 28067
rect 31309 28033 31343 28067
rect 31401 28033 31435 28067
rect 32137 28033 32171 28067
rect 32321 28033 32355 28067
rect 34253 28033 34287 28067
rect 34989 28033 35023 28067
rect 36461 28033 36495 28067
rect 8033 27965 8067 27999
rect 14105 27965 14139 27999
rect 14933 27965 14967 27999
rect 32505 27965 32539 27999
rect 34529 27965 34563 27999
rect 35265 27965 35299 27999
rect 36645 27965 36679 27999
rect 9413 27897 9447 27931
rect 29009 27897 29043 27931
rect 4169 27829 4203 27863
rect 7941 27829 7975 27863
rect 14197 27829 14231 27863
rect 15117 27829 15151 27863
rect 21833 27829 21867 27863
rect 34437 27829 34471 27863
rect 36277 27829 36311 27863
rect 4261 27625 4295 27659
rect 7481 27625 7515 27659
rect 7941 27625 7975 27659
rect 8401 27625 8435 27659
rect 14105 27625 14139 27659
rect 14289 27625 14323 27659
rect 20085 27625 20119 27659
rect 20269 27625 20303 27659
rect 21281 27625 21315 27659
rect 28181 27625 28215 27659
rect 31493 27625 31527 27659
rect 33885 27625 33919 27659
rect 35633 27625 35667 27659
rect 3801 27557 3835 27591
rect 21741 27557 21775 27591
rect 35265 27557 35299 27591
rect 4077 27489 4111 27523
rect 8033 27489 8067 27523
rect 9597 27489 9631 27523
rect 16497 27489 16531 27523
rect 20453 27489 20487 27523
rect 21373 27489 21407 27523
rect 26525 27489 26559 27523
rect 27537 27489 27571 27523
rect 3985 27421 4019 27455
rect 4261 27421 4295 27455
rect 4905 27421 4939 27455
rect 7297 27421 7331 27455
rect 7941 27421 7975 27455
rect 8217 27421 8251 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 16221 27421 16255 27455
rect 20269 27421 20303 27455
rect 20545 27421 20579 27455
rect 21281 27421 21315 27455
rect 21557 27421 21591 27455
rect 22385 27421 22419 27455
rect 22845 27421 22879 27455
rect 28365 27421 28399 27455
rect 31401 27421 31435 27455
rect 31585 27421 31619 27455
rect 34161 27421 34195 27455
rect 35173 27421 35207 27455
rect 35449 27421 35483 27455
rect 36093 27421 36127 27455
rect 9413 27353 9447 27387
rect 14565 27353 14599 27387
rect 27445 27353 27479 27387
rect 33885 27353 33919 27387
rect 4721 27285 4755 27319
rect 5365 27285 5399 27319
rect 22201 27285 22235 27319
rect 26985 27285 27019 27319
rect 27353 27285 27387 27319
rect 28825 27285 28859 27319
rect 29837 27285 29871 27319
rect 33333 27285 33367 27319
rect 34069 27285 34103 27319
rect 5181 27081 5215 27115
rect 7389 27081 7423 27115
rect 13737 27081 13771 27115
rect 15025 27081 15059 27115
rect 15485 27081 15519 27115
rect 26065 27081 26099 27115
rect 29653 27081 29687 27115
rect 34161 27081 34195 27115
rect 9137 27013 9171 27047
rect 14197 27013 14231 27047
rect 22017 27013 22051 27047
rect 25605 27013 25639 27047
rect 26249 27013 26283 27047
rect 26433 27013 26467 27047
rect 30472 27013 30506 27047
rect 1409 26945 1443 26979
rect 2053 26945 2087 26979
rect 4629 26945 4663 26979
rect 7205 26945 7239 26979
rect 7849 26945 7883 26979
rect 9321 26945 9355 26979
rect 10057 26945 10091 26979
rect 13921 26945 13955 26979
rect 14841 26945 14875 26979
rect 15669 26945 15703 26979
rect 20821 26945 20855 26979
rect 21005 26945 21039 26979
rect 21097 26945 21131 26979
rect 21833 26945 21867 26979
rect 23673 26945 23707 26979
rect 29377 26945 29411 26979
rect 30205 26945 30239 26979
rect 34069 26945 34103 26979
rect 34253 26945 34287 26979
rect 34713 26945 34747 26979
rect 34805 26945 34839 26979
rect 34989 26945 35023 26979
rect 35725 26945 35759 26979
rect 8125 26877 8159 26911
rect 14013 26877 14047 26911
rect 26985 26877 27019 26911
rect 27169 26877 27203 26911
rect 27445 26877 27479 26911
rect 36001 26877 36035 26911
rect 20269 26809 20303 26843
rect 34989 26809 35023 26843
rect 1593 26741 1627 26775
rect 4445 26741 4479 26775
rect 9873 26741 9907 26775
rect 10701 26741 10735 26775
rect 14197 26741 14231 26775
rect 20821 26741 20855 26775
rect 21281 26741 21315 26775
rect 31585 26741 31619 26775
rect 33609 26741 33643 26775
rect 7941 26537 7975 26571
rect 15117 26537 15151 26571
rect 15301 26537 15335 26571
rect 20177 26537 20211 26571
rect 20821 26537 20855 26571
rect 21189 26537 21223 26571
rect 30481 26537 30515 26571
rect 14197 26469 14231 26503
rect 38025 26469 38059 26503
rect 3985 26401 4019 26435
rect 4813 26401 4847 26435
rect 10333 26401 10367 26435
rect 10609 26401 10643 26435
rect 10793 26401 10827 26435
rect 14933 26401 14967 26435
rect 20913 26401 20947 26435
rect 22017 26401 22051 26435
rect 23857 26401 23891 26435
rect 26985 26401 27019 26435
rect 27997 26401 28031 26435
rect 3249 26333 3283 26367
rect 3801 26333 3835 26367
rect 6653 26333 6687 26367
rect 6929 26333 6963 26367
rect 8033 26333 8067 26367
rect 8125 26333 8159 26367
rect 12081 26333 12115 26367
rect 14381 26333 14415 26367
rect 15117 26333 15151 26367
rect 18061 26333 18095 26367
rect 20729 26333 20763 26367
rect 21005 26333 21039 26367
rect 24409 26333 24443 26367
rect 30297 26333 30331 26367
rect 37841 26333 37875 26367
rect 7849 26265 7883 26299
rect 14841 26265 14875 26299
rect 22201 26265 22235 26299
rect 27813 26265 27847 26299
rect 8309 26197 8343 26231
rect 3065 25993 3099 26027
rect 3525 25993 3559 26027
rect 24961 25993 24995 26027
rect 27721 25993 27755 26027
rect 29377 25993 29411 26027
rect 30389 25993 30423 26027
rect 3985 25925 4019 25959
rect 7021 25925 7055 25959
rect 10793 25925 10827 25959
rect 22385 25925 22419 25959
rect 27353 25925 27387 25959
rect 28273 25925 28307 25959
rect 1409 25857 1443 25891
rect 2053 25857 2087 25891
rect 2881 25857 2915 25891
rect 3709 25857 3743 25891
rect 7849 25857 7883 25891
rect 8125 25857 8159 25891
rect 12081 25857 12115 25891
rect 15117 25857 15151 25891
rect 15761 25857 15795 25891
rect 17969 25857 18003 25891
rect 24225 25857 24259 25891
rect 24777 25857 24811 25891
rect 25697 25857 25731 25891
rect 27261 25857 27295 25891
rect 30297 25857 30331 25891
rect 34345 25857 34379 25891
rect 34437 25857 34471 25891
rect 34621 25857 34655 25891
rect 35173 25857 35207 25891
rect 35357 25857 35391 25891
rect 3893 25789 3927 25823
rect 8033 25789 8067 25823
rect 8953 25789 8987 25823
rect 9137 25789 9171 25823
rect 12265 25789 12299 25823
rect 13461 25789 13495 25823
rect 18153 25789 18187 25823
rect 19441 25789 19475 25823
rect 24041 25789 24075 25823
rect 25421 25789 25455 25823
rect 27077 25789 27111 25823
rect 30481 25789 30515 25823
rect 35265 25789 35299 25823
rect 14933 25721 14967 25755
rect 15577 25721 15611 25755
rect 33701 25721 33735 25755
rect 34529 25721 34563 25755
rect 1593 25653 1627 25687
rect 3893 25653 3927 25687
rect 7849 25653 7883 25687
rect 8309 25653 8343 25687
rect 29929 25653 29963 25687
rect 34161 25653 34195 25687
rect 2513 25449 2547 25483
rect 4077 25449 4111 25483
rect 9137 25449 9171 25483
rect 9597 25449 9631 25483
rect 14473 25449 14507 25483
rect 15209 25449 15243 25483
rect 17693 25449 17727 25483
rect 21925 25449 21959 25483
rect 22569 25449 22603 25483
rect 23673 25449 23707 25483
rect 23857 25449 23891 25483
rect 24409 25449 24443 25483
rect 30297 25449 30331 25483
rect 2789 25313 2823 25347
rect 3985 25313 4019 25347
rect 15301 25313 15335 25347
rect 24501 25313 24535 25347
rect 1961 25245 1995 25279
rect 2881 25245 2915 25279
rect 4077 25245 4111 25279
rect 4905 25245 4939 25279
rect 7941 25245 7975 25279
rect 8953 25245 8987 25279
rect 14289 25245 14323 25279
rect 15393 25245 15427 25279
rect 16865 25245 16899 25279
rect 17509 25245 17543 25279
rect 18153 25245 18187 25279
rect 21741 25245 21775 25279
rect 22385 25245 22419 25279
rect 23581 25245 23615 25279
rect 23673 25245 23707 25279
rect 24685 25245 24719 25279
rect 29929 25245 29963 25279
rect 30113 25245 30147 25279
rect 2421 25177 2455 25211
rect 3801 25177 3835 25211
rect 15117 25177 15151 25211
rect 23397 25177 23431 25211
rect 24409 25177 24443 25211
rect 3065 25109 3099 25143
rect 4261 25109 4295 25143
rect 4721 25109 4755 25143
rect 7757 25109 7791 25143
rect 15577 25109 15611 25143
rect 17049 25109 17083 25143
rect 24869 25109 24903 25143
rect 26893 25109 26927 25143
rect 27445 25109 27479 25143
rect 8033 24905 8067 24939
rect 29101 24905 29135 24939
rect 15117 24837 15151 24871
rect 17877 24837 17911 24871
rect 24685 24837 24719 24871
rect 2697 24769 2731 24803
rect 4537 24769 4571 24803
rect 5181 24769 5215 24803
rect 7849 24769 7883 24803
rect 13277 24769 13311 24803
rect 15393 24769 15427 24803
rect 23765 24769 23799 24803
rect 24041 24769 24075 24803
rect 28917 24769 28951 24803
rect 30573 24769 30607 24803
rect 35909 24769 35943 24803
rect 36001 24769 36035 24803
rect 36277 24769 36311 24803
rect 2881 24701 2915 24735
rect 13553 24701 13587 24735
rect 15301 24701 15335 24735
rect 17693 24701 17727 24735
rect 18245 24701 18279 24735
rect 23857 24701 23891 24735
rect 4997 24633 5031 24667
rect 8585 24633 8619 24667
rect 15577 24633 15611 24667
rect 24225 24633 24259 24667
rect 5825 24565 5859 24599
rect 15209 24565 15243 24599
rect 23765 24565 23799 24599
rect 28365 24565 28399 24599
rect 30757 24565 30791 24599
rect 34805 24565 34839 24599
rect 35725 24565 35759 24599
rect 36185 24565 36219 24599
rect 1593 24361 1627 24395
rect 14473 24361 14507 24395
rect 30205 24361 30239 24395
rect 15117 24293 15151 24327
rect 29009 24293 29043 24327
rect 36093 24225 36127 24259
rect 36737 24225 36771 24259
rect 1409 24157 1443 24191
rect 2053 24157 2087 24191
rect 7297 24157 7331 24191
rect 12817 24157 12851 24191
rect 14657 24157 14691 24191
rect 15301 24157 15335 24191
rect 19441 24157 19475 24191
rect 29929 24157 29963 24191
rect 30021 24157 30055 24191
rect 30849 24157 30883 24191
rect 31105 24157 31139 24191
rect 33057 24157 33091 24191
rect 33241 24157 33275 24191
rect 34989 24157 35023 24191
rect 35173 24157 35207 24191
rect 35817 24157 35851 24191
rect 35909 24157 35943 24191
rect 36185 24157 36219 24191
rect 36829 24157 36863 24191
rect 28825 24089 28859 24123
rect 33793 24089 33827 24123
rect 35633 24089 35667 24123
rect 12633 24021 12667 24055
rect 22109 24021 22143 24055
rect 32229 24021 32263 24055
rect 33149 24021 33183 24055
rect 35081 24021 35115 24055
rect 37289 24021 37323 24055
rect 13921 23817 13955 23851
rect 29009 23817 29043 23851
rect 29929 23817 29963 23851
rect 30297 23817 30331 23851
rect 37381 23817 37415 23851
rect 11805 23749 11839 23783
rect 14381 23749 14415 23783
rect 14841 23749 14875 23783
rect 18613 23749 18647 23783
rect 29837 23749 29871 23783
rect 35602 23749 35636 23783
rect 6377 23681 6411 23715
rect 7205 23681 7239 23715
rect 14105 23681 14139 23715
rect 15117 23681 15151 23715
rect 20453 23681 20487 23715
rect 22293 23681 22327 23715
rect 27169 23681 27203 23715
rect 32229 23681 32263 23715
rect 32496 23681 32530 23715
rect 34713 23681 34747 23715
rect 34897 23681 34931 23715
rect 35357 23681 35391 23715
rect 37289 23681 37323 23715
rect 7389 23613 7423 23647
rect 9045 23613 9079 23647
rect 11621 23613 11655 23647
rect 13461 23613 13495 23647
rect 14289 23613 14323 23647
rect 15025 23613 15059 23647
rect 20269 23613 20303 23647
rect 29653 23613 29687 23647
rect 34253 23613 34287 23647
rect 22477 23545 22511 23579
rect 36737 23545 36771 23579
rect 6561 23477 6595 23511
rect 14105 23477 14139 23511
rect 14841 23477 14875 23511
rect 15301 23477 15335 23511
rect 16957 23477 16991 23511
rect 22937 23477 22971 23511
rect 26985 23477 27019 23511
rect 33609 23477 33643 23511
rect 34897 23477 34931 23511
rect 6561 23273 6595 23307
rect 7941 23273 7975 23307
rect 11713 23273 11747 23307
rect 13185 23273 13219 23307
rect 14105 23273 14139 23307
rect 14289 23273 14323 23307
rect 27537 23273 27571 23307
rect 36921 23273 36955 23307
rect 5641 23205 5675 23239
rect 15025 23205 15059 23239
rect 6377 23137 6411 23171
rect 14473 23137 14507 23171
rect 16865 23137 16899 23171
rect 22017 23137 22051 23171
rect 23857 23137 23891 23171
rect 1409 23069 1443 23103
rect 2053 23069 2087 23103
rect 2881 23069 2915 23103
rect 3985 23069 4019 23103
rect 5825 23069 5859 23103
rect 6285 23069 6319 23103
rect 6561 23069 6595 23103
rect 7297 23069 7331 23103
rect 8125 23069 8159 23103
rect 8953 23069 8987 23103
rect 12909 23069 12943 23103
rect 13001 23069 13035 23103
rect 13185 23069 13219 23103
rect 14289 23069 14323 23103
rect 14565 23069 14599 23103
rect 15209 23069 15243 23103
rect 16037 23069 16071 23103
rect 26810 23069 26844 23103
rect 27077 23069 27111 23103
rect 27721 23069 27755 23103
rect 27905 23069 27939 23103
rect 35541 23069 35575 23103
rect 35797 23069 35831 23103
rect 17049 23001 17083 23035
rect 18705 23001 18739 23035
rect 22201 23001 22235 23035
rect 1593 22933 1627 22967
rect 3801 22933 3835 22967
rect 5181 22933 5215 22967
rect 6745 22933 6779 22967
rect 7481 22933 7515 22967
rect 12725 22933 12759 22967
rect 16221 22933 16255 22967
rect 25697 22933 25731 22967
rect 5365 22729 5399 22763
rect 6837 22729 6871 22763
rect 14565 22729 14599 22763
rect 27537 22729 27571 22763
rect 30481 22729 30515 22763
rect 36185 22729 36219 22763
rect 2973 22661 3007 22695
rect 5825 22661 5859 22695
rect 6377 22661 6411 22695
rect 7849 22661 7883 22695
rect 9505 22661 9539 22695
rect 19993 22661 20027 22695
rect 27261 22661 27295 22695
rect 34069 22661 34103 22695
rect 2789 22593 2823 22627
rect 4629 22593 4663 22627
rect 5549 22593 5583 22627
rect 6653 22593 6687 22627
rect 7665 22593 7699 22627
rect 14749 22593 14783 22627
rect 24685 22593 24719 22627
rect 26985 22593 27019 22627
rect 27169 22593 27203 22627
rect 27353 22593 27387 22627
rect 30573 22593 30607 22627
rect 33885 22593 33919 22627
rect 35633 22593 35667 22627
rect 36277 22593 36311 22627
rect 5733 22525 5767 22559
rect 6561 22525 6595 22559
rect 10977 22525 11011 22559
rect 11529 22525 11563 22559
rect 11713 22525 11747 22559
rect 13277 22525 13311 22559
rect 18153 22525 18187 22559
rect 18337 22525 18371 22559
rect 24225 22525 24259 22559
rect 24501 22525 24535 22559
rect 26341 22457 26375 22491
rect 5825 22389 5859 22423
rect 6561 22389 6595 22423
rect 6469 22185 6503 22219
rect 13185 22185 13219 22219
rect 18245 22185 18279 22219
rect 6377 22049 6411 22083
rect 13001 22049 13035 22083
rect 20821 22049 20855 22083
rect 22753 22049 22787 22083
rect 25697 22049 25731 22083
rect 26433 22049 26467 22083
rect 29929 22049 29963 22083
rect 36277 22049 36311 22083
rect 6469 21981 6503 22015
rect 7297 21981 7331 22015
rect 10425 21981 10459 22015
rect 11713 21981 11747 22015
rect 12909 21981 12943 22015
rect 13185 21981 13219 22015
rect 19257 21981 19291 22015
rect 22477 21981 22511 22015
rect 27721 21981 27755 22015
rect 31953 21981 31987 22015
rect 36185 21981 36219 22015
rect 37841 21981 37875 22015
rect 6193 21913 6227 21947
rect 20637 21913 20671 21947
rect 26249 21913 26283 21947
rect 30113 21913 30147 21947
rect 36093 21913 36127 21947
rect 6653 21845 6687 21879
rect 7113 21845 7147 21879
rect 11529 21845 11563 21879
rect 12725 21845 12759 21879
rect 19441 21845 19475 21879
rect 27537 21845 27571 21879
rect 32045 21845 32079 21879
rect 35725 21845 35759 21879
rect 37381 21845 37415 21879
rect 38025 21845 38059 21879
rect 11897 21641 11931 21675
rect 13553 21641 13587 21675
rect 17141 21641 17175 21675
rect 28825 21641 28859 21675
rect 36277 21641 36311 21675
rect 6837 21573 6871 21607
rect 27252 21573 27286 21607
rect 1409 21505 1443 21539
rect 2053 21505 2087 21539
rect 6561 21505 6595 21539
rect 6653 21505 6687 21539
rect 7481 21505 7515 21539
rect 12081 21505 12115 21539
rect 13737 21505 13771 21539
rect 14565 21505 14599 21539
rect 17233 21505 17267 21539
rect 20269 21505 20303 21539
rect 20821 21505 20855 21539
rect 22109 21505 22143 21539
rect 26985 21505 27019 21539
rect 29009 21505 29043 21539
rect 29193 21505 29227 21539
rect 32689 21505 32723 21539
rect 36369 21505 36403 21539
rect 14289 21437 14323 21471
rect 21833 21437 21867 21471
rect 30021 21437 30055 21471
rect 30297 21437 30331 21471
rect 36461 21437 36495 21471
rect 21005 21369 21039 21403
rect 1593 21301 1627 21335
rect 5825 21301 5859 21335
rect 6377 21301 6411 21335
rect 6561 21301 6595 21335
rect 7297 21301 7331 21335
rect 28365 21301 28399 21335
rect 32597 21301 32631 21335
rect 35909 21301 35943 21335
rect 2513 21097 2547 21131
rect 14197 21097 14231 21131
rect 21097 21097 21131 21131
rect 21373 21097 21407 21131
rect 28549 21097 28583 21131
rect 29745 21097 29779 21131
rect 31953 21097 31987 21131
rect 6561 20961 6595 20995
rect 6745 20961 6779 20995
rect 10333 20961 10367 20995
rect 10517 20961 10551 20995
rect 15025 20961 15059 20995
rect 16313 20961 16347 20995
rect 16589 20961 16623 20995
rect 18153 20961 18187 20995
rect 21005 20961 21039 20995
rect 24685 20961 24719 20995
rect 30573 20961 30607 20995
rect 2513 20893 2547 20927
rect 2605 20893 2639 20927
rect 5641 20893 5675 20927
rect 15301 20893 15335 20927
rect 18429 20893 18463 20927
rect 19625 20893 19659 20927
rect 19901 20893 19935 20927
rect 21189 20893 21223 20927
rect 21833 20893 21867 20927
rect 24409 20893 24443 20927
rect 27997 20893 28031 20927
rect 28365 20893 28399 20927
rect 29561 20893 29595 20927
rect 8401 20825 8435 20859
rect 12173 20825 12207 20859
rect 20913 20825 20947 20859
rect 28181 20825 28215 20859
rect 28273 20825 28307 20859
rect 30840 20825 30874 20859
rect 1409 20757 1443 20791
rect 2881 20757 2915 20791
rect 5457 20757 5491 20791
rect 22017 20757 22051 20791
rect 27445 20757 27479 20791
rect 17141 20553 17175 20587
rect 19441 20553 19475 20587
rect 20729 20553 20763 20587
rect 31033 20553 31067 20587
rect 3525 20485 3559 20519
rect 3709 20485 3743 20519
rect 16681 20485 16715 20519
rect 24501 20485 24535 20519
rect 34437 20485 34471 20519
rect 1409 20417 1443 20451
rect 2421 20417 2455 20451
rect 2789 20417 2823 20451
rect 2881 20417 2915 20451
rect 7849 20417 7883 20451
rect 14657 20417 14691 20451
rect 16957 20417 16991 20451
rect 19533 20417 19567 20451
rect 20269 20417 20303 20451
rect 20545 20417 20579 20451
rect 24685 20417 24719 20451
rect 30389 20417 30423 20451
rect 30573 20417 30607 20451
rect 31217 20417 31251 20451
rect 34621 20417 34655 20451
rect 34713 20417 34747 20451
rect 35265 20417 35299 20451
rect 35449 20417 35483 20451
rect 14381 20349 14415 20383
rect 15853 20349 15887 20383
rect 16129 20349 16163 20383
rect 16773 20349 16807 20383
rect 20361 20349 20395 20383
rect 24225 20349 24259 20383
rect 30205 20349 30239 20383
rect 1593 20281 1627 20315
rect 21925 20281 21959 20315
rect 2513 20213 2547 20247
rect 3065 20213 3099 20247
rect 3893 20213 3927 20247
rect 4721 20213 4755 20247
rect 7665 20213 7699 20247
rect 10517 20213 10551 20247
rect 16681 20213 16715 20247
rect 18797 20213 18831 20247
rect 20545 20213 20579 20247
rect 35357 20213 35391 20247
rect 3801 20009 3835 20043
rect 13369 20009 13403 20043
rect 18061 20009 18095 20043
rect 18521 20009 18555 20043
rect 20913 20009 20947 20043
rect 37657 20009 37691 20043
rect 3157 19941 3191 19975
rect 19441 19941 19475 19975
rect 20269 19941 20303 19975
rect 37013 19941 37047 19975
rect 3893 19873 3927 19907
rect 4721 19873 4755 19907
rect 4905 19873 4939 19907
rect 12081 19873 12115 19907
rect 13185 19873 13219 19907
rect 15025 19873 15059 19907
rect 16037 19873 16071 19907
rect 16773 19873 16807 19907
rect 18153 19873 18187 19907
rect 23857 19873 23891 19907
rect 30297 19873 30331 19907
rect 1869 19805 1903 19839
rect 2973 19805 3007 19839
rect 3249 19805 3283 19839
rect 3801 19805 3835 19839
rect 4077 19805 4111 19839
rect 13093 19805 13127 19839
rect 13369 19805 13403 19839
rect 14749 19805 14783 19839
rect 16313 19805 16347 19839
rect 17049 19805 17083 19839
rect 18337 19805 18371 19839
rect 19257 19805 19291 19839
rect 21465 19805 21499 19839
rect 22109 19805 22143 19839
rect 27445 19805 27479 19839
rect 30481 19805 30515 19839
rect 35449 19805 35483 19839
rect 35679 19805 35713 19839
rect 35817 19805 35851 19839
rect 35909 19805 35943 19839
rect 36369 19805 36403 19839
rect 37013 19805 37047 19839
rect 37197 19805 37231 19839
rect 6561 19737 6595 19771
rect 10241 19737 10275 19771
rect 11897 19737 11931 19771
rect 18061 19737 18095 19771
rect 20085 19737 20119 19771
rect 20821 19737 20855 19771
rect 25605 19737 25639 19771
rect 27261 19737 27295 19771
rect 30665 19737 30699 19771
rect 35541 19737 35575 19771
rect 1961 19669 1995 19703
rect 2789 19669 2823 19703
rect 4261 19669 4295 19703
rect 12909 19669 12943 19703
rect 21649 19669 21683 19703
rect 27997 19669 28031 19703
rect 31309 19669 31343 19703
rect 35265 19669 35299 19703
rect 36461 19669 36495 19703
rect 3525 19465 3559 19499
rect 11805 19465 11839 19499
rect 18797 19465 18831 19499
rect 23305 19465 23339 19499
rect 24501 19465 24535 19499
rect 25145 19465 25179 19499
rect 29745 19465 29779 19499
rect 30389 19465 30423 19499
rect 34535 19465 34569 19499
rect 35357 19465 35391 19499
rect 3065 19397 3099 19431
rect 9137 19397 9171 19431
rect 10149 19397 10183 19431
rect 10333 19397 10367 19431
rect 13369 19397 13403 19431
rect 14013 19397 14047 19431
rect 16681 19397 16715 19431
rect 19441 19397 19475 19431
rect 19533 19397 19567 19431
rect 22845 19397 22879 19431
rect 29469 19397 29503 19431
rect 30849 19397 30883 19431
rect 32229 19397 32263 19431
rect 34621 19397 34655 19431
rect 3341 19329 3375 19363
rect 11621 19329 11655 19363
rect 13093 19329 13127 19363
rect 13185 19329 13219 19363
rect 14933 19329 14967 19363
rect 16129 19329 16163 19363
rect 16865 19329 16899 19363
rect 16957 19329 16991 19363
rect 18613 19329 18647 19363
rect 19625 19329 19659 19363
rect 20177 19329 20211 19363
rect 22201 19329 22235 19363
rect 23121 19329 23155 19363
rect 24317 19329 24351 19363
rect 24961 19329 24995 19363
rect 29193 19329 29227 19363
rect 29377 19329 29411 19363
rect 29561 19329 29595 19363
rect 30757 19329 30791 19363
rect 32137 19329 32171 19363
rect 32321 19329 32355 19363
rect 32781 19329 32815 19363
rect 34437 19329 34471 19363
rect 34713 19329 34747 19363
rect 35173 19329 35207 19363
rect 35357 19329 35391 19363
rect 3157 19261 3191 19295
rect 14657 19261 14691 19295
rect 19993 19261 20027 19295
rect 23029 19261 23063 19295
rect 30941 19261 30975 19295
rect 28733 19193 28767 19227
rect 33885 19193 33919 19227
rect 3065 19125 3099 19159
rect 6469 19125 6503 19159
rect 9045 19125 9079 19159
rect 12909 19125 12943 19159
rect 13369 19125 13403 19159
rect 14105 19125 14139 19159
rect 15945 19125 15979 19159
rect 16681 19125 16715 19159
rect 17141 19125 17175 19159
rect 17969 19125 18003 19159
rect 22385 19125 22419 19159
rect 22845 19125 22879 19159
rect 1593 18921 1627 18955
rect 4077 18921 4111 18955
rect 21465 18921 21499 18955
rect 22109 18921 22143 18955
rect 22937 18921 22971 18955
rect 23397 18921 23431 18955
rect 31585 18921 31619 18955
rect 35449 18921 35483 18955
rect 37749 18921 37783 18955
rect 4261 18853 4295 18887
rect 5549 18853 5583 18887
rect 4169 18785 4203 18819
rect 4390 18785 4424 18819
rect 15025 18785 15059 18819
rect 22201 18785 22235 18819
rect 23029 18785 23063 18819
rect 25789 18785 25823 18819
rect 26985 18785 27019 18819
rect 30941 18785 30975 18819
rect 33241 18785 33275 18819
rect 34069 18785 34103 18819
rect 34805 18785 34839 18819
rect 1409 18717 1443 18751
rect 2053 18717 2087 18751
rect 4537 18717 4571 18751
rect 5365 18717 5399 18751
rect 6837 18717 6871 18751
rect 7297 18717 7331 18751
rect 10333 18717 10367 18751
rect 10793 18717 10827 18751
rect 15301 18717 15335 18751
rect 16405 18717 16439 18751
rect 18705 18717 18739 18751
rect 19533 18717 19567 18751
rect 22017 18717 22051 18751
rect 22293 18717 22327 18751
rect 23213 18717 23247 18751
rect 27169 18717 27203 18751
rect 27629 18717 27663 18751
rect 32045 18717 32079 18751
rect 36369 18717 36403 18751
rect 36625 18717 36659 18751
rect 6653 18649 6687 18683
rect 10977 18649 11011 18683
rect 12633 18649 12667 18683
rect 16589 18649 16623 18683
rect 22937 18649 22971 18683
rect 31217 18649 31251 18683
rect 32689 18649 32723 18683
rect 7481 18581 7515 18615
rect 14473 18581 14507 18615
rect 19349 18581 19383 18615
rect 20085 18581 20119 18615
rect 22477 18581 22511 18615
rect 30389 18581 30423 18615
rect 31125 18581 31159 18615
rect 32229 18581 32263 18615
rect 34989 18581 35023 18615
rect 35081 18581 35115 18615
rect 5733 18377 5767 18411
rect 7113 18377 7147 18411
rect 11989 18377 12023 18411
rect 17601 18377 17635 18411
rect 22109 18377 22143 18411
rect 23305 18377 23339 18411
rect 26341 18377 26375 18411
rect 27445 18377 27479 18411
rect 28273 18377 28307 18411
rect 33609 18377 33643 18411
rect 36001 18377 36035 18411
rect 36737 18377 36771 18411
rect 18245 18309 18279 18343
rect 18429 18309 18463 18343
rect 22845 18309 22879 18343
rect 23765 18309 23799 18343
rect 6377 18241 6411 18275
rect 7205 18241 7239 18275
rect 7757 18241 7791 18275
rect 8401 18241 8435 18275
rect 12173 18241 12207 18275
rect 13737 18241 13771 18275
rect 14013 18241 14047 18275
rect 14657 18241 14691 18275
rect 14933 18241 14967 18275
rect 21925 18241 21959 18275
rect 23029 18241 23063 18275
rect 23121 18241 23155 18275
rect 24777 18241 24811 18275
rect 32229 18241 32263 18275
rect 32485 18241 32519 18275
rect 35541 18241 35575 18275
rect 36553 18241 36587 18275
rect 37841 18241 37875 18275
rect 13921 18173 13955 18207
rect 14749 18173 14783 18207
rect 25053 18173 25087 18207
rect 27169 18173 27203 18207
rect 27353 18173 27387 18207
rect 35633 18173 35667 18207
rect 8585 18105 8619 18139
rect 4721 18037 4755 18071
rect 6561 18037 6595 18071
rect 7941 18037 7975 18071
rect 9045 18037 9079 18071
rect 13553 18037 13587 18071
rect 13829 18037 13863 18071
rect 14473 18037 14507 18071
rect 14657 18037 14691 18071
rect 22937 18037 22971 18071
rect 27813 18037 27847 18071
rect 35357 18037 35391 18071
rect 37289 18037 37323 18071
rect 38025 18037 38059 18071
rect 7481 17833 7515 17867
rect 7941 17833 7975 17867
rect 14657 17833 14691 17867
rect 21833 17833 21867 17867
rect 22937 17833 22971 17867
rect 29561 17833 29595 17867
rect 1593 17765 1627 17799
rect 18337 17765 18371 17799
rect 7573 17697 7607 17731
rect 8953 17697 8987 17731
rect 9137 17697 9171 17731
rect 9689 17697 9723 17731
rect 14749 17697 14783 17731
rect 22937 17697 22971 17731
rect 26525 17697 26559 17731
rect 27721 17697 27755 17731
rect 30113 17697 30147 17731
rect 1409 17629 1443 17663
rect 2053 17629 2087 17663
rect 7757 17629 7791 17663
rect 12357 17629 12391 17663
rect 13369 17629 13403 17663
rect 14933 17629 14967 17663
rect 17601 17629 17635 17663
rect 22753 17629 22787 17663
rect 23029 17629 23063 17663
rect 26341 17629 26375 17663
rect 28641 17629 28675 17663
rect 28825 17629 28859 17663
rect 7481 17561 7515 17595
rect 14657 17561 14691 17595
rect 18153 17561 18187 17595
rect 30297 17561 30331 17595
rect 31953 17561 31987 17595
rect 6929 17493 6963 17527
rect 13185 17493 13219 17527
rect 15117 17493 15151 17527
rect 23213 17493 23247 17527
rect 29009 17493 29043 17527
rect 8769 17289 8803 17323
rect 22661 17289 22695 17323
rect 30113 17289 30147 17323
rect 4629 17221 4663 17255
rect 6837 17221 6871 17255
rect 12541 17221 12575 17255
rect 28825 17221 28859 17255
rect 7113 17153 7147 17187
rect 7757 17153 7791 17187
rect 8033 17153 8067 17187
rect 12357 17153 12391 17187
rect 23765 17153 23799 17187
rect 26985 17153 27019 17187
rect 27252 17153 27286 17187
rect 34621 17153 34655 17187
rect 35081 17153 35115 17187
rect 35244 17156 35278 17190
rect 35360 17156 35394 17190
rect 35449 17153 35483 17187
rect 2789 17085 2823 17119
rect 2973 17085 3007 17119
rect 7021 17085 7055 17119
rect 7849 17085 7883 17119
rect 14013 17085 14047 17119
rect 17785 17085 17819 17119
rect 17969 17085 18003 17119
rect 19349 17085 19383 17119
rect 24041 17085 24075 17119
rect 29653 17085 29687 17119
rect 28365 17017 28399 17051
rect 29929 17017 29963 17051
rect 7113 16949 7147 16983
rect 7297 16949 7331 16983
rect 7757 16949 7791 16983
rect 8217 16949 8251 16983
rect 35725 16949 35759 16983
rect 2881 16745 2915 16779
rect 6929 16745 6963 16779
rect 7573 16745 7607 16779
rect 9045 16745 9079 16779
rect 17877 16745 17911 16779
rect 27353 16745 27387 16779
rect 6745 16609 6779 16643
rect 7665 16609 7699 16643
rect 13553 16609 13587 16643
rect 26065 16609 26099 16643
rect 26341 16609 26375 16643
rect 35633 16609 35667 16643
rect 3801 16541 3835 16575
rect 6653 16541 6687 16575
rect 6929 16541 6963 16575
rect 7573 16541 7607 16575
rect 7849 16541 7883 16575
rect 14657 16541 14691 16575
rect 15577 16541 15611 16575
rect 27537 16541 27571 16575
rect 35900 16541 35934 16575
rect 7113 16405 7147 16439
rect 8033 16405 8067 16439
rect 14473 16405 14507 16439
rect 15761 16405 15795 16439
rect 20177 16405 20211 16439
rect 37013 16405 37047 16439
rect 2881 16201 2915 16235
rect 3341 16201 3375 16235
rect 17877 16201 17911 16235
rect 18981 16201 19015 16235
rect 22845 16201 22879 16235
rect 23765 16201 23799 16235
rect 30757 16201 30791 16235
rect 3801 16133 3835 16167
rect 14105 16133 14139 16167
rect 18521 16133 18555 16167
rect 23305 16133 23339 16167
rect 26157 16133 26191 16167
rect 1409 16065 1443 16099
rect 2053 16065 2087 16099
rect 2697 16065 2731 16099
rect 3525 16065 3559 16099
rect 4261 16065 4295 16099
rect 13093 16065 13127 16099
rect 13921 16065 13955 16099
rect 18061 16065 18095 16099
rect 18797 16065 18831 16099
rect 20729 16065 20763 16099
rect 21833 16065 21867 16099
rect 23489 16065 23523 16099
rect 23581 16065 23615 16099
rect 32873 16065 32907 16099
rect 33885 16065 33919 16099
rect 3709 15997 3743 16031
rect 7665 15997 7699 16031
rect 7849 15997 7883 16031
rect 9505 15997 9539 16031
rect 15761 15997 15795 16031
rect 18613 15997 18647 16031
rect 20453 15997 20487 16031
rect 24685 15997 24719 16031
rect 26341 15997 26375 16031
rect 34069 15997 34103 16031
rect 34529 15997 34563 16031
rect 33057 15929 33091 15963
rect 1593 15861 1627 15895
rect 3801 15861 3835 15895
rect 4445 15861 4479 15895
rect 4905 15861 4939 15895
rect 12081 15861 12115 15895
rect 12909 15861 12943 15895
rect 18705 15861 18739 15895
rect 19901 15861 19935 15895
rect 22017 15861 22051 15895
rect 23305 15861 23339 15895
rect 29561 15861 29595 15895
rect 32137 15861 32171 15895
rect 7205 15657 7239 15691
rect 7849 15657 7883 15691
rect 18245 15657 18279 15691
rect 18705 15657 18739 15691
rect 23397 15657 23431 15691
rect 29009 15657 29043 15691
rect 34897 15657 34931 15691
rect 37749 15657 37783 15691
rect 32321 15589 32355 15623
rect 3801 15521 3835 15555
rect 4261 15521 4295 15555
rect 11713 15521 11747 15555
rect 11897 15521 11931 15555
rect 13553 15521 13587 15555
rect 15669 15521 15703 15555
rect 16681 15521 16715 15555
rect 19257 15521 19291 15555
rect 19533 15521 19567 15555
rect 21281 15521 21315 15555
rect 22109 15521 22143 15555
rect 23581 15521 23615 15555
rect 24685 15521 24719 15555
rect 26525 15521 26559 15555
rect 30113 15521 30147 15555
rect 30205 15521 30239 15555
rect 30941 15521 30975 15555
rect 32873 15521 32907 15555
rect 34805 15521 34839 15555
rect 34989 15521 35023 15555
rect 3065 15453 3099 15487
rect 7665 15453 7699 15487
rect 9137 15453 9171 15487
rect 11253 15453 11287 15487
rect 15485 15453 15519 15487
rect 18429 15453 18463 15487
rect 18521 15453 18555 15487
rect 20545 15453 20579 15487
rect 20637 15453 20671 15487
rect 20821 15453 20855 15487
rect 22385 15453 22419 15487
rect 23673 15453 23707 15487
rect 31125 15453 31159 15487
rect 31217 15453 31251 15487
rect 33149 15453 33183 15487
rect 34713 15453 34747 15487
rect 36369 15453 36403 15487
rect 3985 15385 4019 15419
rect 18705 15385 18739 15419
rect 23397 15385 23431 15419
rect 26341 15385 26375 15419
rect 35909 15385 35943 15419
rect 36614 15385 36648 15419
rect 3249 15317 3283 15351
rect 8953 15317 8987 15351
rect 23857 15317 23891 15351
rect 29653 15317 29687 15351
rect 30021 15317 30055 15351
rect 31585 15317 31619 15351
rect 13829 15113 13863 15147
rect 22753 15113 22787 15147
rect 34621 15113 34655 15147
rect 35633 15113 35667 15147
rect 4721 15045 4755 15079
rect 8677 15045 8711 15079
rect 13369 15045 13403 15079
rect 22293 15045 22327 15079
rect 23857 15045 23891 15079
rect 1409 14977 1443 15011
rect 2053 14977 2087 15011
rect 4905 14977 4939 15011
rect 7757 14977 7791 15011
rect 11529 14977 11563 15011
rect 14013 14977 14047 15011
rect 14289 14977 14323 15011
rect 15485 14977 15519 15011
rect 20545 14977 20579 15011
rect 21097 14977 21131 15011
rect 22569 14977 22603 15011
rect 23213 14977 23247 15011
rect 28181 14977 28215 15011
rect 28641 14977 28675 15011
rect 30490 14977 30524 15011
rect 30757 14977 30791 15011
rect 32137 14977 32171 15011
rect 32321 14977 32355 15011
rect 32505 14977 32539 15011
rect 35449 14977 35483 15011
rect 3341 14909 3375 14943
rect 8493 14909 8527 14943
rect 10333 14909 10367 14943
rect 11713 14909 11747 14943
rect 14105 14909 14139 14943
rect 18797 14909 18831 14943
rect 19073 14909 19107 14943
rect 22385 14909 22419 14943
rect 28825 14841 28859 14875
rect 29377 14841 29411 14875
rect 1593 14773 1627 14807
rect 7297 14773 7331 14807
rect 7941 14773 7975 14807
rect 14289 14773 14323 14807
rect 17969 14773 18003 14807
rect 21281 14773 21315 14807
rect 22385 14773 22419 14807
rect 23397 14773 23431 14807
rect 31493 14773 31527 14807
rect 2513 14569 2547 14603
rect 3801 14569 3835 14603
rect 4169 14569 4203 14603
rect 8953 14569 8987 14603
rect 21925 14569 21959 14603
rect 22201 14569 22235 14603
rect 22845 14569 22879 14603
rect 28733 14569 28767 14603
rect 30573 14569 30607 14603
rect 34805 14569 34839 14603
rect 2605 14433 2639 14467
rect 4077 14433 4111 14467
rect 13093 14433 13127 14467
rect 15025 14433 15059 14467
rect 15301 14433 15335 14467
rect 21925 14433 21959 14467
rect 24685 14433 24719 14467
rect 25697 14433 25731 14467
rect 2513 14365 2547 14399
rect 2789 14365 2823 14399
rect 3985 14365 4019 14399
rect 8033 14365 8067 14399
rect 13369 14365 13403 14399
rect 18245 14365 18279 14399
rect 19257 14365 19291 14399
rect 19533 14365 19567 14399
rect 21097 14365 21131 14399
rect 21741 14365 21775 14399
rect 22017 14365 22051 14399
rect 22661 14365 22695 14399
rect 24409 14365 24443 14399
rect 25973 14365 26007 14399
rect 28181 14365 28215 14399
rect 29561 14365 29595 14399
rect 29745 14365 29779 14399
rect 29929 14365 29963 14399
rect 30389 14365 30423 14399
rect 34713 14365 34747 14399
rect 35357 14365 35391 14399
rect 4261 14297 4295 14331
rect 17417 14297 17451 14331
rect 37381 14297 37415 14331
rect 38025 14297 38059 14331
rect 2973 14229 3007 14263
rect 7849 14229 7883 14263
rect 17509 14229 17543 14263
rect 18061 14229 18095 14263
rect 21281 14229 21315 14263
rect 28089 14229 28123 14263
rect 37933 14229 37967 14263
rect 3433 14025 3467 14059
rect 5089 14025 5123 14059
rect 13277 14025 13311 14059
rect 14657 14025 14691 14059
rect 22109 14025 22143 14059
rect 32597 14025 32631 14059
rect 3893 13957 3927 13991
rect 4353 13957 4387 13991
rect 7941 13957 7975 13991
rect 13737 13957 13771 13991
rect 34069 13957 34103 13991
rect 3617 13889 3651 13923
rect 4537 13889 4571 13923
rect 7757 13889 7791 13923
rect 12357 13889 12391 13923
rect 13461 13889 13495 13923
rect 14841 13889 14875 13923
rect 17509 13889 17543 13923
rect 20545 13889 20579 13923
rect 20821 13889 20855 13923
rect 24593 13889 24627 13923
rect 30573 13889 30607 13923
rect 32413 13889 32447 13923
rect 3801 13821 3835 13855
rect 8309 13821 8343 13855
rect 13645 13821 13679 13855
rect 17233 13821 17267 13855
rect 20637 13821 20671 13855
rect 24869 13821 24903 13855
rect 30021 13821 30055 13855
rect 33885 13821 33919 13855
rect 35541 13821 35575 13855
rect 30757 13753 30791 13787
rect 3893 13685 3927 13719
rect 12541 13685 12575 13719
rect 13737 13685 13771 13719
rect 20361 13685 20395 13719
rect 20821 13685 20855 13719
rect 1593 13481 1627 13515
rect 4445 13481 4479 13515
rect 17417 13481 17451 13515
rect 21097 13481 21131 13515
rect 21925 13481 21959 13515
rect 30113 13481 30147 13515
rect 5089 13413 5123 13447
rect 17877 13413 17911 13447
rect 22201 13413 22235 13447
rect 16497 13345 16531 13379
rect 17601 13345 17635 13379
rect 20177 13345 20211 13379
rect 21005 13345 21039 13379
rect 21833 13345 21867 13379
rect 25605 13345 25639 13379
rect 26893 13345 26927 13379
rect 28549 13345 28583 13379
rect 1409 13277 1443 13311
rect 2053 13277 2087 13311
rect 3985 13277 4019 13311
rect 4629 13277 4663 13311
rect 5273 13277 5307 13311
rect 5733 13277 5767 13311
rect 7757 13277 7791 13311
rect 16773 13277 16807 13311
rect 17693 13277 17727 13311
rect 19901 13277 19935 13311
rect 20821 13277 20855 13311
rect 21097 13277 21131 13311
rect 21741 13277 21775 13311
rect 22017 13277 22051 13311
rect 25881 13277 25915 13311
rect 28733 13277 28767 13311
rect 34805 13277 34839 13311
rect 34989 13277 35023 13311
rect 17417 13209 17451 13243
rect 30021 13209 30055 13243
rect 21281 13141 21315 13175
rect 34897 13141 34931 13175
rect 29745 12937 29779 12971
rect 34621 12937 34655 12971
rect 7941 12869 7975 12903
rect 9597 12869 9631 12903
rect 12633 12869 12667 12903
rect 13553 12869 13587 12903
rect 18153 12869 18187 12903
rect 19809 12869 19843 12903
rect 21925 12869 21959 12903
rect 22937 12869 22971 12903
rect 23857 12869 23891 12903
rect 27445 12869 27479 12903
rect 7757 12801 7791 12835
rect 12357 12801 12391 12835
rect 13277 12801 13311 12835
rect 22201 12801 22235 12835
rect 23213 12801 23247 12835
rect 24133 12801 24167 12835
rect 35081 12801 35115 12835
rect 35265 12801 35299 12835
rect 35357 12801 35391 12835
rect 35449 12801 35483 12835
rect 2973 12733 3007 12767
rect 3433 12733 3467 12767
rect 3617 12733 3651 12767
rect 5273 12733 5307 12767
rect 12541 12733 12575 12767
rect 13369 12733 13403 12767
rect 19993 12733 20027 12767
rect 22109 12733 22143 12767
rect 23029 12733 23063 12767
rect 23949 12733 23983 12767
rect 29101 12733 29135 12767
rect 29285 12733 29319 12767
rect 17693 12665 17727 12699
rect 10241 12597 10275 12631
rect 12173 12597 12207 12631
rect 12633 12597 12667 12631
rect 13093 12597 13127 12631
rect 13553 12597 13587 12631
rect 21925 12597 21959 12631
rect 22385 12597 22419 12631
rect 22937 12597 22971 12631
rect 23397 12597 23431 12631
rect 23857 12597 23891 12631
rect 24317 12597 24351 12631
rect 35725 12597 35759 12631
rect 3249 12393 3283 12427
rect 4077 12393 4111 12427
rect 6285 12393 6319 12427
rect 12633 12393 12667 12427
rect 17049 12393 17083 12427
rect 21649 12393 21683 12427
rect 22477 12393 22511 12427
rect 32597 12393 32631 12427
rect 37381 12393 37415 12427
rect 11253 12257 11287 12291
rect 11713 12257 11747 12291
rect 12541 12257 12575 12291
rect 17141 12257 17175 12291
rect 18153 12257 18187 12291
rect 22293 12257 22327 12291
rect 25973 12257 26007 12291
rect 27261 12257 27295 12291
rect 29837 12257 29871 12291
rect 1409 12189 1443 12223
rect 2053 12189 2087 12223
rect 3065 12189 3099 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4261 12189 4295 12223
rect 4905 12189 4939 12223
rect 9229 12189 9263 12223
rect 12449 12189 12483 12223
rect 13369 12189 13403 12223
rect 16957 12189 16991 12223
rect 17233 12189 17267 12223
rect 17877 12189 17911 12223
rect 22201 12189 22235 12223
rect 22477 12189 22511 12223
rect 25237 12189 25271 12223
rect 25789 12189 25823 12223
rect 33057 12189 33091 12223
rect 33241 12189 33275 12223
rect 33333 12189 33367 12223
rect 33425 12189 33459 12223
rect 36001 12189 36035 12223
rect 36257 12189 36291 12223
rect 11529 12121 11563 12155
rect 12725 12121 12759 12155
rect 14197 12121 14231 12155
rect 25053 12121 25087 12155
rect 30082 12121 30116 12155
rect 1593 12053 1627 12087
rect 3801 12053 3835 12087
rect 4721 12053 4755 12087
rect 12265 12053 12299 12087
rect 13185 12053 13219 12087
rect 17417 12053 17451 12087
rect 22661 12053 22695 12087
rect 31217 12053 31251 12087
rect 33701 12053 33735 12087
rect 35449 12053 35483 12087
rect 6561 11849 6595 11883
rect 8309 11849 8343 11883
rect 17785 11849 17819 11883
rect 28365 11849 28399 11883
rect 33241 11849 33275 11883
rect 35173 11849 35207 11883
rect 4169 11781 4203 11815
rect 10977 11781 11011 11815
rect 13185 11781 13219 11815
rect 17325 11781 17359 11815
rect 29929 11781 29963 11815
rect 30849 11781 30883 11815
rect 31033 11781 31067 11815
rect 34038 11781 34072 11815
rect 6377 11713 6411 11747
rect 8033 11713 8067 11747
rect 9137 11713 9171 11747
rect 12081 11713 12115 11747
rect 12357 11713 12391 11747
rect 13461 11713 13495 11747
rect 15945 11713 15979 11747
rect 17049 11713 17083 11747
rect 17141 11713 17175 11747
rect 24593 11713 24627 11747
rect 29377 11713 29411 11747
rect 29469 11713 29503 11747
rect 29653 11713 29687 11747
rect 29745 11713 29779 11747
rect 30665 11713 30699 11747
rect 32597 11713 32631 11747
rect 33793 11713 33827 11747
rect 3985 11645 4019 11679
rect 5825 11645 5859 11679
rect 9321 11645 9355 11679
rect 13277 11645 13311 11679
rect 24869 11645 24903 11679
rect 16865 11577 16899 11611
rect 13461 11509 13495 11543
rect 13645 11509 13679 11543
rect 16129 11509 16163 11543
rect 17049 11509 17083 11543
rect 20361 11509 20395 11543
rect 28825 11509 28859 11543
rect 32689 11509 32723 11543
rect 3985 11305 4019 11339
rect 4261 11305 4295 11339
rect 6837 11305 6871 11339
rect 7573 11305 7607 11339
rect 10609 11305 10643 11339
rect 13461 11305 13495 11339
rect 19349 11305 19383 11339
rect 20637 11305 20671 11339
rect 21649 11305 21683 11339
rect 29561 11305 29595 11339
rect 30481 11305 30515 11339
rect 19901 11237 19935 11271
rect 27077 11237 27111 11271
rect 12265 11169 12299 11203
rect 13369 11169 13403 11203
rect 16221 11169 16255 11203
rect 16681 11169 16715 11203
rect 22201 11169 22235 11203
rect 29929 11169 29963 11203
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 5273 11101 5307 11135
rect 5549 11101 5583 11135
rect 6653 11101 6687 11135
rect 7389 11101 7423 11135
rect 8401 11101 8435 11135
rect 10793 11101 10827 11135
rect 11989 11101 12023 11135
rect 13277 11101 13311 11135
rect 13553 11101 13587 11135
rect 14105 11101 14139 11135
rect 15577 11101 15611 11135
rect 16037 11101 16071 11135
rect 18521 11101 18555 11135
rect 22477 11101 22511 11135
rect 25237 11101 25271 11135
rect 25697 11101 25731 11135
rect 29745 11101 29779 11135
rect 34897 11101 34931 11135
rect 34989 11101 35023 11135
rect 35173 11101 35207 11135
rect 35265 11101 35299 11135
rect 35910 11101 35944 11135
rect 36093 11101 36127 11135
rect 3801 11033 3835 11067
rect 25964 11033 25998 11067
rect 34713 11033 34747 11067
rect 35725 11033 35759 11067
rect 8217 10965 8251 10999
rect 13093 10965 13127 10999
rect 14289 10965 14323 10999
rect 18337 10965 18371 10999
rect 21097 10965 21131 10999
rect 3617 10761 3651 10795
rect 5365 10761 5399 10795
rect 7113 10761 7147 10795
rect 8033 10761 8067 10795
rect 26985 10761 27019 10795
rect 27353 10761 27387 10795
rect 30573 10761 30607 10795
rect 33609 10761 33643 10795
rect 35081 10761 35115 10795
rect 17417 10693 17451 10727
rect 19073 10693 19107 10727
rect 19901 10693 19935 10727
rect 24685 10693 24719 10727
rect 28733 10693 28767 10727
rect 28917 10693 28951 10727
rect 29653 10693 29687 10727
rect 34253 10693 34287 10727
rect 1409 10625 1443 10659
rect 2053 10625 2087 10659
rect 3157 10625 3191 10659
rect 3433 10625 3467 10659
rect 4445 10625 4479 10659
rect 5181 10625 5215 10659
rect 6377 10625 6411 10659
rect 13093 10625 13127 10659
rect 19533 10625 19567 10659
rect 19717 10625 19751 10659
rect 20821 10625 20855 10659
rect 22017 10625 22051 10659
rect 22109 10625 22143 10659
rect 22385 10625 22419 10659
rect 27169 10625 27203 10659
rect 27445 10625 27479 10659
rect 29469 10625 29503 10659
rect 35081 10625 35115 10659
rect 35265 10625 35299 10659
rect 3249 10557 3283 10591
rect 17233 10557 17267 10591
rect 20913 10557 20947 10591
rect 21833 10557 21867 10591
rect 24409 10557 24443 10591
rect 24869 10557 24903 10591
rect 34529 10557 34563 10591
rect 6561 10489 6595 10523
rect 1593 10421 1627 10455
rect 3157 10421 3191 10455
rect 10425 10421 10459 10455
rect 12909 10421 12943 10455
rect 13737 10421 13771 10455
rect 20821 10421 20855 10455
rect 21189 10421 21223 10455
rect 2973 10217 3007 10251
rect 6009 10217 6043 10251
rect 17325 10217 17359 10251
rect 20821 10217 20855 10251
rect 28181 10217 28215 10251
rect 2789 10149 2823 10183
rect 6653 10149 6687 10183
rect 19533 10149 19567 10183
rect 20269 10149 20303 10183
rect 21741 10149 21775 10183
rect 4537 10081 4571 10115
rect 14105 10081 14139 10115
rect 14289 10081 14323 10115
rect 15945 10081 15979 10115
rect 20913 10081 20947 10115
rect 27353 10081 27387 10115
rect 30757 10081 30791 10115
rect 2973 10013 3007 10047
rect 3065 10013 3099 10047
rect 4813 10013 4847 10047
rect 5825 10013 5859 10047
rect 7665 10013 7699 10047
rect 10425 10013 10459 10047
rect 12265 10013 12299 10047
rect 12725 10013 12759 10047
rect 20085 10013 20119 10047
rect 20821 10013 20855 10047
rect 22293 10013 22327 10047
rect 23121 10013 23155 10047
rect 27537 10013 27571 10047
rect 29653 10013 29687 10047
rect 29837 10013 29871 10047
rect 29929 10013 29963 10047
rect 30021 10013 30055 10047
rect 38117 10013 38151 10047
rect 3249 9945 3283 9979
rect 7849 9945 7883 9979
rect 10609 9945 10643 9979
rect 25697 9945 25731 9979
rect 28089 9945 28123 9979
rect 31002 9945 31036 9979
rect 16497 9877 16531 9911
rect 18613 9877 18647 9911
rect 21189 9877 21223 9911
rect 22477 9877 22511 9911
rect 22937 9877 22971 9911
rect 30297 9877 30331 9911
rect 32137 9877 32171 9911
rect 19349 9673 19383 9707
rect 21005 9673 21039 9707
rect 26985 9673 27019 9707
rect 29653 9673 29687 9707
rect 7481 9605 7515 9639
rect 12449 9605 12483 9639
rect 14105 9605 14139 9639
rect 17601 9605 17635 9639
rect 18613 9605 18647 9639
rect 19257 9605 19291 9639
rect 22109 9605 22143 9639
rect 26341 9605 26375 9639
rect 30113 9605 30147 9639
rect 30297 9605 30331 9639
rect 32137 9605 32171 9639
rect 1409 9537 1443 9571
rect 2237 9537 2271 9571
rect 2329 9537 2363 9571
rect 3157 9537 3191 9571
rect 3341 9537 3375 9571
rect 3709 9537 3743 9571
rect 4077 9537 4111 9571
rect 4813 9537 4847 9571
rect 6377 9537 6411 9571
rect 15669 9537 15703 9571
rect 15945 9537 15979 9571
rect 16681 9537 16715 9571
rect 16957 9537 16991 9571
rect 19441 9537 19475 9571
rect 26157 9537 26191 9571
rect 26433 9537 26467 9571
rect 27169 9537 27203 9571
rect 27353 9537 27387 9571
rect 27445 9537 27479 9571
rect 29285 9537 29319 9571
rect 29469 9537 29503 9571
rect 35613 9537 35647 9571
rect 5089 9469 5123 9503
rect 12265 9469 12299 9503
rect 15209 9469 15243 9503
rect 15761 9469 15795 9503
rect 16865 9469 16899 9503
rect 19809 9469 19843 9503
rect 19993 9469 20027 9503
rect 22661 9469 22695 9503
rect 22845 9469 22879 9503
rect 23673 9469 23707 9503
rect 25421 9469 25455 9503
rect 28549 9469 28583 9503
rect 35357 9469 35391 9503
rect 4261 9401 4295 9435
rect 20453 9401 20487 9435
rect 27905 9401 27939 9435
rect 32413 9401 32447 9435
rect 1593 9333 1627 9367
rect 15945 9333 15979 9367
rect 16129 9333 16163 9367
rect 16681 9333 16715 9367
rect 17141 9333 17175 9367
rect 22017 9333 22051 9367
rect 25973 9333 26007 9367
rect 30481 9333 30515 9367
rect 32597 9333 32631 9367
rect 34805 9333 34839 9367
rect 36737 9333 36771 9367
rect 2513 9129 2547 9163
rect 2973 9129 3007 9163
rect 4905 9129 4939 9163
rect 8217 9129 8251 9163
rect 16589 9129 16623 9163
rect 20545 9129 20579 9163
rect 26985 9129 27019 9163
rect 29009 9129 29043 9163
rect 29653 9129 29687 9163
rect 35357 9129 35391 9163
rect 1409 9061 1443 9095
rect 19349 9061 19383 9095
rect 2605 8993 2639 9027
rect 2789 8925 2823 8959
rect 4445 8925 4479 8959
rect 4997 8925 5031 8959
rect 7389 8925 7423 8959
rect 7665 8925 7699 8959
rect 26157 8925 26191 8959
rect 26433 8925 26467 8959
rect 31033 8925 31067 8959
rect 34713 8925 34747 8959
rect 34897 8925 34931 8959
rect 34989 8925 35023 8959
rect 35081 8925 35115 8959
rect 2513 8857 2547 8891
rect 5549 8857 5583 8891
rect 30766 8857 30800 8891
rect 25973 8789 26007 8823
rect 26341 8789 26375 8823
rect 5825 8585 5859 8619
rect 8861 8585 8895 8619
rect 10425 8585 10459 8619
rect 29101 8585 29135 8619
rect 29653 8585 29687 8619
rect 30757 8585 30791 8619
rect 34437 8585 34471 8619
rect 9413 8517 9447 8551
rect 22477 8517 22511 8551
rect 24133 8517 24167 8551
rect 4445 8449 4479 8483
rect 7205 8449 7239 8483
rect 7665 8449 7699 8483
rect 8309 8449 8343 8483
rect 9689 8449 9723 8483
rect 17141 8449 17175 8483
rect 25605 8449 25639 8483
rect 30113 8449 30147 8483
rect 30297 8449 30331 8483
rect 30389 8449 30423 8483
rect 30481 8449 30515 8483
rect 34713 8449 34747 8483
rect 37289 8449 37323 8483
rect 6929 8381 6963 8415
rect 9505 8381 9539 8415
rect 22293 8381 22327 8415
rect 25881 8381 25915 8415
rect 34437 8381 34471 8415
rect 9873 8313 9907 8347
rect 34621 8313 34655 8347
rect 37473 8313 37507 8347
rect 3709 8245 3743 8279
rect 7849 8245 7883 8279
rect 9413 8245 9447 8279
rect 17325 8245 17359 8279
rect 1593 8041 1627 8075
rect 6653 8041 6687 8075
rect 8217 8041 8251 8075
rect 9229 8041 9263 8075
rect 26709 8041 26743 8075
rect 3801 7905 3835 7939
rect 5641 7905 5675 7939
rect 8033 7905 8067 7939
rect 9045 7905 9079 7939
rect 11069 7905 11103 7939
rect 24869 7905 24903 7939
rect 25329 7905 25363 7939
rect 1409 7837 1443 7871
rect 2053 7837 2087 7871
rect 7205 7837 7239 7871
rect 7941 7837 7975 7871
rect 8217 7837 8251 7871
rect 9229 7837 9263 7871
rect 11345 7837 11379 7871
rect 14289 7837 14323 7871
rect 16589 7837 16623 7871
rect 20729 7837 20763 7871
rect 21465 7837 21499 7871
rect 25596 7837 25630 7871
rect 3985 7769 4019 7803
rect 8953 7769 8987 7803
rect 7389 7701 7423 7735
rect 8401 7701 8435 7735
rect 9413 7701 9447 7735
rect 14105 7701 14139 7735
rect 16773 7701 16807 7735
rect 20913 7701 20947 7735
rect 3617 7497 3651 7531
rect 8861 7497 8895 7531
rect 7757 7429 7791 7463
rect 9689 7429 9723 7463
rect 14013 7429 14047 7463
rect 17601 7429 17635 7463
rect 28917 7429 28951 7463
rect 3433 7361 3467 7395
rect 4077 7361 4111 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 23213 7361 23247 7395
rect 30573 7361 30607 7395
rect 30757 7361 30791 7395
rect 30849 7361 30883 7395
rect 30941 7361 30975 7395
rect 34161 7361 34195 7395
rect 34345 7361 34379 7395
rect 5273 7293 5307 7327
rect 5549 7293 5583 7327
rect 6377 7293 6411 7327
rect 13737 7293 13771 7327
rect 14197 7293 14231 7327
rect 17417 7293 17451 7327
rect 18889 7293 18923 7327
rect 23305 7293 23339 7327
rect 23397 7293 23431 7327
rect 27261 7293 27295 7327
rect 29101 7293 29135 7327
rect 24133 7225 24167 7259
rect 4261 7157 4295 7191
rect 7849 7157 7883 7191
rect 8217 7157 8251 7191
rect 9781 7157 9815 7191
rect 22845 7157 22879 7191
rect 30021 7157 30055 7191
rect 31217 7157 31251 7191
rect 34253 7157 34287 7191
rect 4261 6953 4295 6987
rect 4721 6953 4755 6987
rect 5181 6953 5215 6987
rect 7849 6953 7883 6987
rect 30297 6953 30331 6987
rect 33885 6953 33919 6987
rect 4169 6817 4203 6851
rect 4997 6817 5031 6851
rect 7849 6817 7883 6851
rect 10609 6817 10643 6851
rect 16773 6817 16807 6851
rect 18429 6817 18463 6851
rect 19441 6817 19475 6851
rect 20729 6817 20763 6851
rect 23121 6817 23155 6851
rect 24501 6817 24535 6851
rect 35817 6817 35851 6851
rect 36369 6817 36403 6851
rect 1409 6749 1443 6783
rect 2053 6749 2087 6783
rect 3985 6749 4019 6783
rect 4905 6749 4939 6783
rect 8033 6749 8067 6783
rect 8953 6749 8987 6783
rect 10885 6749 10919 6783
rect 14105 6749 14139 6783
rect 14473 6749 14507 6783
rect 16589 6749 16623 6783
rect 19257 6749 19291 6783
rect 23213 6749 23247 6783
rect 30205 6749 30239 6783
rect 30389 6749 30423 6783
rect 34161 6749 34195 6783
rect 34989 6749 35023 6783
rect 35081 6749 35115 6783
rect 35173 6749 35207 6783
rect 35357 6749 35391 6783
rect 4261 6681 4295 6715
rect 5181 6681 5215 6715
rect 7757 6681 7791 6715
rect 14289 6681 14323 6715
rect 14381 6681 14415 6715
rect 23305 6681 23339 6715
rect 33885 6681 33919 6715
rect 36614 6681 36648 6715
rect 1593 6613 1627 6647
rect 3801 6613 3835 6647
rect 8217 6613 8251 6647
rect 9137 6613 9171 6647
rect 14657 6613 14691 6647
rect 15117 6613 15151 6647
rect 23673 6613 23707 6647
rect 34069 6613 34103 6647
rect 34713 6613 34747 6647
rect 37749 6613 37783 6647
rect 14565 6409 14599 6443
rect 16773 6409 16807 6443
rect 20637 6409 20671 6443
rect 22477 6409 22511 6443
rect 23949 6409 23983 6443
rect 33057 6409 33091 6443
rect 5641 6341 5675 6375
rect 12992 6341 13026 6375
rect 22385 6341 22419 6375
rect 27537 6341 27571 6375
rect 35642 6341 35676 6375
rect 5365 6273 5399 6307
rect 8401 6273 8435 6307
rect 14749 6273 14783 6307
rect 19073 6273 19107 6307
rect 32965 6273 32999 6307
rect 33149 6273 33183 6307
rect 34069 6273 34103 6307
rect 35909 6273 35943 6307
rect 37841 6273 37875 6307
rect 2697 6205 2731 6239
rect 2881 6205 2915 6239
rect 3249 6205 3283 6239
rect 5457 6205 5491 6239
rect 12725 6205 12759 6239
rect 14933 6205 14967 6239
rect 22293 6205 22327 6239
rect 33977 6205 34011 6239
rect 14105 6137 14139 6171
rect 27353 6137 27387 6171
rect 33701 6137 33735 6171
rect 5181 6069 5215 6103
rect 5365 6069 5399 6103
rect 8585 6069 8619 6103
rect 15485 6069 15519 6103
rect 19165 6069 19199 6103
rect 22845 6069 22879 6103
rect 33885 6069 33919 6103
rect 34529 6069 34563 6103
rect 38025 6069 38059 6103
rect 2697 5865 2731 5899
rect 3801 5865 3835 5899
rect 4813 5865 4847 5899
rect 14197 5865 14231 5899
rect 34713 5865 34747 5899
rect 17693 5797 17727 5831
rect 30205 5797 30239 5831
rect 33149 5797 33183 5831
rect 4905 5729 4939 5763
rect 9137 5729 9171 5763
rect 13093 5729 13127 5763
rect 13553 5729 13587 5763
rect 16773 5729 16807 5763
rect 22937 5729 22971 5763
rect 23121 5729 23155 5763
rect 33057 5729 33091 5763
rect 3985 5661 4019 5695
rect 4721 5661 4755 5695
rect 8953 5661 8987 5695
rect 15945 5661 15979 5695
rect 16313 5661 16347 5695
rect 16957 5661 16991 5695
rect 20085 5661 20119 5695
rect 20177 5661 20211 5695
rect 20453 5661 20487 5695
rect 23213 5661 23247 5695
rect 30113 5661 30147 5695
rect 32965 5661 32999 5695
rect 33241 5661 33275 5695
rect 4997 5593 5031 5627
rect 10793 5593 10827 5627
rect 13369 5593 13403 5627
rect 16037 5593 16071 5627
rect 16129 5593 16163 5627
rect 20269 5593 20303 5627
rect 4537 5525 4571 5559
rect 15761 5525 15795 5559
rect 17141 5525 17175 5559
rect 19901 5525 19935 5559
rect 21097 5525 21131 5559
rect 23581 5525 23615 5559
rect 32781 5525 32815 5559
rect 33793 5525 33827 5559
rect 1593 5321 1627 5355
rect 3709 5321 3743 5355
rect 15301 5321 15335 5355
rect 16681 5321 16715 5355
rect 22109 5321 22143 5355
rect 22477 5321 22511 5355
rect 22569 5321 22603 5355
rect 24685 5321 24719 5355
rect 25145 5321 25179 5355
rect 27445 5321 27479 5355
rect 29193 5321 29227 5355
rect 30297 5321 30331 5355
rect 32873 5321 32907 5355
rect 34253 5321 34287 5355
rect 4169 5253 4203 5287
rect 10333 5253 10367 5287
rect 13461 5253 13495 5287
rect 17049 5253 17083 5287
rect 20821 5253 20855 5287
rect 23489 5253 23523 5287
rect 27353 5253 27387 5287
rect 33609 5253 33643 5287
rect 1409 5185 1443 5219
rect 2053 5185 2087 5219
rect 3249 5185 3283 5219
rect 3893 5185 3927 5219
rect 5457 5185 5491 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 12081 5185 12115 5219
rect 13277 5185 13311 5219
rect 13369 5185 13403 5219
rect 13645 5185 13679 5219
rect 14197 5185 14231 5219
rect 15945 5185 15979 5219
rect 16865 5185 16899 5219
rect 16957 5185 16991 5219
rect 17233 5185 17267 5219
rect 17693 5185 17727 5219
rect 18981 5185 19015 5219
rect 19625 5185 19659 5219
rect 20545 5185 20579 5219
rect 20729 5185 20763 5219
rect 20949 5185 20983 5219
rect 23305 5185 23339 5219
rect 23581 5185 23615 5219
rect 23673 5185 23707 5219
rect 25053 5185 25087 5219
rect 25973 5185 26007 5219
rect 29190 5185 29224 5219
rect 30294 5185 30328 5219
rect 32781 5185 32815 5219
rect 32965 5185 32999 5219
rect 33425 5185 33459 5219
rect 33701 5185 33735 5219
rect 34161 5185 34195 5219
rect 4077 5117 4111 5151
rect 10057 5117 10091 5151
rect 10517 5117 10551 5151
rect 16129 5117 16163 5151
rect 19809 5117 19843 5151
rect 22753 5117 22787 5151
rect 25329 5117 25363 5151
rect 27537 5117 27571 5151
rect 29653 5117 29687 5151
rect 30757 5117 30791 5151
rect 12633 5049 12667 5083
rect 26985 5049 27019 5083
rect 29561 5049 29595 5083
rect 30665 5049 30699 5083
rect 3065 4981 3099 5015
rect 4169 4981 4203 5015
rect 4629 4981 4663 5015
rect 5273 4981 5307 5015
rect 11529 4981 11563 5015
rect 13093 4981 13127 5015
rect 15761 4981 15795 5015
rect 19441 4981 19475 5015
rect 20545 4981 20579 5015
rect 23857 4981 23891 5015
rect 29009 4981 29043 5015
rect 30113 4981 30147 5015
rect 33425 4981 33459 5015
rect 16773 4777 16807 4811
rect 20637 4777 20671 4811
rect 23489 4777 23523 4811
rect 25329 4777 25363 4811
rect 26893 4777 26927 4811
rect 28917 4777 28951 4811
rect 34161 4777 34195 4811
rect 5089 4641 5123 4675
rect 6745 4641 6779 4675
rect 12541 4641 12575 4675
rect 22569 4641 22603 4675
rect 24777 4641 24811 4675
rect 27353 4641 27387 4675
rect 27537 4641 27571 4675
rect 30205 4641 30239 4675
rect 31493 4641 31527 4675
rect 2697 4573 2731 4607
rect 4261 4573 4295 4607
rect 4905 4573 4939 4607
rect 9689 4573 9723 4607
rect 9873 4573 9907 4607
rect 10517 4573 10551 4607
rect 10609 4573 10643 4607
rect 10885 4573 10919 4607
rect 11437 4573 11471 4607
rect 12357 4573 12391 4607
rect 15393 4573 15427 4607
rect 17417 4573 17451 4607
rect 19257 4573 19291 4607
rect 21281 4573 21315 4607
rect 21465 4573 21499 4607
rect 21925 4573 21959 4607
rect 22753 4573 22787 4607
rect 22937 4573 22971 4607
rect 23581 4573 23615 4607
rect 24593 4573 24627 4607
rect 27261 4573 27295 4607
rect 28273 4573 28307 4607
rect 28457 4573 28491 4607
rect 29561 4573 29595 4607
rect 29745 4573 29779 4607
rect 32045 4573 32079 4607
rect 32229 4573 32263 4607
rect 32781 4573 32815 4607
rect 33048 4573 33082 4607
rect 9045 4505 9079 4539
rect 10701 4505 10735 4539
rect 15660 4505 15694 4539
rect 19502 4505 19536 4539
rect 21373 4505 21407 4539
rect 4445 4437 4479 4471
rect 9505 4437 9539 4471
rect 10333 4437 10367 4471
rect 17233 4437 17267 4471
rect 17969 4437 18003 4471
rect 24409 4437 24443 4471
rect 28365 4437 28399 4471
rect 29653 4437 29687 4471
rect 32137 4437 32171 4471
rect 8309 4233 8343 4267
rect 15761 4233 15795 4267
rect 18245 4233 18279 4267
rect 19349 4233 19383 4267
rect 23213 4233 23247 4267
rect 27629 4233 27663 4267
rect 30849 4233 30883 4267
rect 32689 4233 32723 4267
rect 2881 4165 2915 4199
rect 17132 4165 17166 4199
rect 28742 4165 28776 4199
rect 1409 4097 1443 4131
rect 2053 4097 2087 4131
rect 2697 4097 2731 4131
rect 4997 4097 5031 4131
rect 9422 4097 9456 4131
rect 10333 4097 10367 4131
rect 12541 4097 12575 4131
rect 13001 4097 13035 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 13921 4097 13955 4131
rect 15945 4097 15979 4131
rect 19165 4097 19199 4131
rect 20729 4097 20763 4131
rect 21833 4097 21867 4131
rect 22100 4097 22134 4131
rect 24409 4097 24443 4131
rect 29736 4097 29770 4131
rect 3893 4029 3927 4063
rect 9689 4029 9723 4063
rect 10517 4029 10551 4063
rect 16865 4029 16899 4063
rect 23765 4029 23799 4063
rect 29009 4029 29043 4063
rect 29469 4029 29503 4063
rect 1593 3893 1627 3927
rect 10149 3893 10183 3927
rect 11621 3893 11655 3927
rect 12357 3893 12391 3927
rect 24593 3893 24627 3927
rect 2513 3689 2547 3723
rect 14105 3689 14139 3723
rect 18337 3689 18371 3723
rect 25973 3689 26007 3723
rect 29561 3689 29595 3723
rect 30113 3689 30147 3723
rect 31033 3689 31067 3723
rect 32965 3689 32999 3723
rect 2881 3621 2915 3655
rect 8401 3621 8435 3655
rect 10333 3621 10367 3655
rect 10885 3621 10919 3655
rect 13553 3621 13587 3655
rect 2605 3553 2639 3587
rect 4537 3553 4571 3587
rect 8953 3553 8987 3587
rect 12173 3553 12207 3587
rect 24593 3553 24627 3587
rect 31585 3553 31619 3587
rect 2513 3485 2547 3519
rect 8217 3485 8251 3519
rect 12440 3485 12474 3519
rect 24849 3485 24883 3519
rect 4721 3417 4755 3451
rect 6377 3417 6411 3451
rect 9198 3417 9232 3451
rect 31852 3417 31886 3451
rect 2789 3145 2823 3179
rect 9321 3145 9355 3179
rect 10517 3145 10551 3179
rect 24501 3145 24535 3179
rect 2881 3009 2915 3043
rect 9505 3009 9539 3043
rect 1409 2805 1443 2839
rect 2053 2805 2087 2839
rect 2513 2601 2547 2635
rect 3801 2601 3835 2635
rect 2053 2533 2087 2567
rect 2697 2397 2731 2431
rect 3157 2397 3191 2431
rect 3985 2397 4019 2431
rect 4445 2397 4479 2431
rect 37841 2397 37875 2431
rect 1869 2329 1903 2363
rect 38025 2261 38059 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 3418 37408 3424 37460
rect 3476 37448 3482 37460
rect 23934 37448 23940 37460
rect 3476 37420 23940 37448
rect 3476 37408 3482 37420
rect 23934 37408 23940 37420
rect 23992 37408 23998 37460
rect 38010 37448 38016 37460
rect 37971 37420 38016 37448
rect 38010 37408 38016 37420
rect 38068 37408 38074 37460
rect 3234 37340 3240 37392
rect 3292 37380 3298 37392
rect 13354 37380 13360 37392
rect 3292 37352 13360 37380
rect 3292 37340 3298 37352
rect 13354 37340 13360 37352
rect 13412 37340 13418 37392
rect 16758 37312 16764 37324
rect 16719 37284 16764 37312
rect 16758 37272 16764 37284
rect 16816 37272 16822 37324
rect 22186 37204 22192 37256
rect 22244 37244 22250 37256
rect 22281 37247 22339 37253
rect 22281 37244 22293 37247
rect 22244 37216 22293 37244
rect 22244 37204 22250 37216
rect 22281 37213 22293 37216
rect 22327 37213 22339 37247
rect 22281 37207 22339 37213
rect 29914 37204 29920 37256
rect 29972 37244 29978 37256
rect 30009 37247 30067 37253
rect 30009 37244 30021 37247
rect 29972 37216 30021 37244
rect 29972 37204 29978 37216
rect 30009 37213 30021 37216
rect 30055 37213 30067 37247
rect 37829 37247 37887 37253
rect 37829 37244 37841 37247
rect 30009 37207 30067 37213
rect 37660 37216 37841 37244
rect 37660 37120 37688 37216
rect 37829 37213 37841 37216
rect 37875 37213 37887 37247
rect 37829 37207 37887 37213
rect 29178 37068 29184 37120
rect 29236 37108 29242 37120
rect 30193 37111 30251 37117
rect 30193 37108 30205 37111
rect 29236 37080 30205 37108
rect 29236 37068 29242 37080
rect 30193 37077 30205 37080
rect 30239 37077 30251 37111
rect 30193 37071 30251 37077
rect 37369 37111 37427 37117
rect 37369 37077 37381 37111
rect 37415 37108 37427 37111
rect 37642 37108 37648 37120
rect 37415 37080 37648 37108
rect 37415 37077 37427 37080
rect 37369 37071 37427 37077
rect 37642 37068 37648 37080
rect 37700 37068 37706 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 29914 36904 29920 36916
rect 29875 36876 29920 36904
rect 29914 36864 29920 36876
rect 29972 36864 29978 36916
rect 13357 36839 13415 36845
rect 13357 36805 13369 36839
rect 13403 36836 13415 36839
rect 14366 36836 14372 36848
rect 13403 36808 14372 36836
rect 13403 36805 13415 36808
rect 13357 36799 13415 36805
rect 14366 36796 14372 36808
rect 14424 36796 14430 36848
rect 22186 36768 22192 36780
rect 22147 36740 22192 36768
rect 22186 36728 22192 36740
rect 22244 36728 22250 36780
rect 2314 36660 2320 36712
rect 2372 36700 2378 36712
rect 2685 36703 2743 36709
rect 2685 36700 2697 36703
rect 2372 36672 2697 36700
rect 2372 36660 2378 36672
rect 2685 36669 2697 36672
rect 2731 36669 2743 36703
rect 2866 36700 2872 36712
rect 2827 36672 2872 36700
rect 2685 36663 2743 36669
rect 2866 36660 2872 36672
rect 2924 36660 2930 36712
rect 4154 36700 4160 36712
rect 4115 36672 4160 36700
rect 4154 36660 4160 36672
rect 4212 36700 4218 36712
rect 4706 36700 4712 36712
rect 4212 36672 4712 36700
rect 4212 36660 4218 36672
rect 4706 36660 4712 36672
rect 4764 36660 4770 36712
rect 12894 36660 12900 36712
rect 12952 36700 12958 36712
rect 13173 36703 13231 36709
rect 13173 36700 13185 36703
rect 12952 36672 13185 36700
rect 12952 36660 12958 36672
rect 13173 36669 13185 36672
rect 13219 36669 13231 36703
rect 13814 36700 13820 36712
rect 13775 36672 13820 36700
rect 13173 36663 13231 36669
rect 13814 36660 13820 36672
rect 13872 36660 13878 36712
rect 22370 36700 22376 36712
rect 22331 36672 22376 36700
rect 22370 36660 22376 36672
rect 22428 36660 22434 36712
rect 22649 36703 22707 36709
rect 22649 36669 22661 36703
rect 22695 36669 22707 36703
rect 22649 36663 22707 36669
rect 22094 36592 22100 36644
rect 22152 36632 22158 36644
rect 22664 36632 22692 36663
rect 22152 36604 22692 36632
rect 22152 36592 22158 36604
rect 4614 36524 4620 36576
rect 4672 36564 4678 36576
rect 4985 36567 5043 36573
rect 4985 36564 4997 36567
rect 4672 36536 4997 36564
rect 4672 36524 4678 36536
rect 4985 36533 4997 36536
rect 5031 36533 5043 36567
rect 4985 36527 5043 36533
rect 8938 36524 8944 36576
rect 8996 36564 9002 36576
rect 9033 36567 9091 36573
rect 9033 36564 9045 36567
rect 8996 36536 9045 36564
rect 8996 36524 9002 36536
rect 9033 36533 9045 36536
rect 9079 36533 9091 36567
rect 9033 36527 9091 36533
rect 17405 36567 17463 36573
rect 17405 36533 17417 36567
rect 17451 36564 17463 36567
rect 18690 36564 18696 36576
rect 17451 36536 18696 36564
rect 17451 36533 17463 36536
rect 17405 36527 17463 36533
rect 18690 36524 18696 36536
rect 18748 36524 18754 36576
rect 25406 36524 25412 36576
rect 25464 36564 25470 36576
rect 25501 36567 25559 36573
rect 25501 36564 25513 36567
rect 25464 36536 25513 36564
rect 25464 36524 25470 36536
rect 25501 36533 25513 36536
rect 25547 36533 25559 36567
rect 25501 36527 25559 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 2314 36360 2320 36372
rect 2275 36332 2320 36360
rect 2314 36320 2320 36332
rect 2372 36320 2378 36372
rect 12894 36360 12900 36372
rect 12855 36332 12900 36360
rect 12894 36320 12900 36332
rect 12952 36320 12958 36372
rect 3970 36252 3976 36304
rect 4028 36292 4034 36304
rect 5534 36292 5540 36304
rect 4028 36264 5540 36292
rect 4028 36252 4034 36264
rect 5534 36252 5540 36264
rect 5592 36252 5598 36304
rect 4062 36184 4068 36236
rect 4120 36224 4126 36236
rect 5261 36227 5319 36233
rect 5261 36224 5273 36227
rect 4120 36196 5273 36224
rect 4120 36184 4126 36196
rect 5261 36193 5273 36196
rect 5307 36224 5319 36227
rect 6914 36224 6920 36236
rect 5307 36196 6920 36224
rect 5307 36193 5319 36196
rect 5261 36187 5319 36193
rect 6914 36184 6920 36196
rect 6972 36184 6978 36236
rect 9401 36227 9459 36233
rect 9401 36224 9413 36227
rect 8312 36196 9413 36224
rect 2774 36156 2780 36168
rect 2735 36128 2780 36156
rect 2774 36116 2780 36128
rect 2832 36116 2838 36168
rect 4341 36159 4399 36165
rect 4341 36125 4353 36159
rect 4387 36156 4399 36159
rect 4801 36159 4859 36165
rect 4801 36156 4813 36159
rect 4387 36128 4813 36156
rect 4387 36125 4399 36128
rect 4341 36119 4399 36125
rect 4801 36125 4813 36128
rect 4847 36125 4859 36159
rect 4801 36119 4859 36125
rect 4982 36088 4988 36100
rect 4943 36060 4988 36088
rect 4982 36048 4988 36060
rect 5040 36048 5046 36100
rect 8312 36088 8340 36196
rect 9401 36193 9413 36196
rect 9447 36224 9459 36227
rect 13541 36227 13599 36233
rect 9447 36196 11744 36224
rect 9447 36193 9459 36196
rect 9401 36187 9459 36193
rect 8389 36159 8447 36165
rect 8389 36125 8401 36159
rect 8435 36156 8447 36159
rect 8941 36159 8999 36165
rect 8941 36156 8953 36159
rect 8435 36128 8953 36156
rect 8435 36125 8447 36128
rect 8389 36119 8447 36125
rect 8941 36125 8953 36128
rect 8987 36125 8999 36159
rect 8941 36119 8999 36125
rect 6886 36060 8340 36088
rect 9125 36091 9183 36097
rect 5534 35980 5540 36032
rect 5592 36020 5598 36032
rect 6886 36020 6914 36060
rect 9125 36057 9137 36091
rect 9171 36088 9183 36091
rect 9582 36088 9588 36100
rect 9171 36060 9588 36088
rect 9171 36057 9183 36060
rect 9125 36051 9183 36057
rect 9582 36048 9588 36060
rect 9640 36048 9646 36100
rect 11716 36088 11744 36196
rect 13541 36193 13553 36227
rect 13587 36224 13599 36227
rect 15933 36227 15991 36233
rect 15933 36224 15945 36227
rect 13587 36196 15945 36224
rect 13587 36193 13599 36196
rect 13541 36187 13599 36193
rect 15933 36193 15945 36196
rect 15979 36193 15991 36227
rect 18690 36224 18696 36236
rect 18651 36196 18696 36224
rect 15933 36187 15991 36193
rect 18690 36184 18696 36196
rect 18748 36184 18754 36236
rect 22094 36224 22100 36236
rect 22055 36196 22100 36224
rect 22094 36184 22100 36196
rect 22152 36184 22158 36236
rect 23474 36184 23480 36236
rect 23532 36224 23538 36236
rect 24397 36227 24455 36233
rect 24397 36224 24409 36227
rect 23532 36196 24409 36224
rect 23532 36184 23538 36196
rect 24397 36193 24409 36196
rect 24443 36193 24455 36227
rect 25406 36224 25412 36236
rect 25367 36196 25412 36224
rect 24397 36187 24455 36193
rect 25406 36184 25412 36196
rect 25464 36184 25470 36236
rect 12069 36159 12127 36165
rect 12069 36125 12081 36159
rect 12115 36156 12127 36159
rect 13630 36156 13636 36168
rect 12115 36128 13636 36156
rect 12115 36125 12127 36128
rect 12069 36119 12127 36125
rect 13630 36116 13636 36128
rect 13688 36116 13694 36168
rect 21177 36159 21235 36165
rect 21177 36125 21189 36159
rect 21223 36156 21235 36159
rect 21637 36159 21695 36165
rect 21637 36156 21649 36159
rect 21223 36128 21649 36156
rect 21223 36125 21235 36128
rect 21177 36119 21235 36125
rect 21637 36125 21649 36128
rect 21683 36125 21695 36159
rect 30926 36156 30932 36168
rect 30887 36128 30932 36156
rect 21637 36119 21695 36125
rect 30926 36116 30932 36128
rect 30984 36116 30990 36168
rect 13814 36088 13820 36100
rect 11716 36060 13820 36088
rect 13814 36048 13820 36060
rect 13872 36088 13878 36100
rect 14093 36091 14151 36097
rect 14093 36088 14105 36091
rect 13872 36060 14105 36088
rect 13872 36048 13878 36060
rect 14093 36057 14105 36060
rect 14139 36057 14151 36091
rect 14093 36051 14151 36057
rect 15749 36091 15807 36097
rect 15749 36057 15761 36091
rect 15795 36057 15807 36091
rect 16850 36088 16856 36100
rect 16811 36060 16856 36088
rect 15749 36051 15807 36057
rect 5592 35992 6914 36020
rect 15764 36020 15792 36051
rect 16850 36048 16856 36060
rect 16908 36048 16914 36100
rect 18509 36091 18567 36097
rect 18509 36057 18521 36091
rect 18555 36088 18567 36091
rect 19334 36088 19340 36100
rect 18555 36060 19340 36088
rect 18555 36057 18567 36060
rect 18509 36051 18567 36057
rect 19334 36048 19340 36060
rect 19392 36048 19398 36100
rect 21818 36088 21824 36100
rect 21779 36060 21824 36088
rect 21818 36048 21824 36060
rect 21876 36048 21882 36100
rect 25590 36088 25596 36100
rect 25551 36060 25596 36088
rect 25590 36048 25596 36060
rect 25648 36048 25654 36100
rect 27246 36088 27252 36100
rect 27207 36060 27252 36088
rect 27246 36048 27252 36060
rect 27304 36048 27310 36100
rect 30374 36048 30380 36100
rect 30432 36088 30438 36100
rect 30662 36091 30720 36097
rect 30662 36088 30674 36091
rect 30432 36060 30674 36088
rect 30432 36048 30438 36060
rect 30662 36057 30674 36060
rect 30708 36057 30720 36091
rect 30662 36051 30720 36057
rect 18414 36020 18420 36032
rect 15764 35992 18420 36020
rect 5592 35980 5598 35992
rect 18414 35980 18420 35992
rect 18472 35980 18478 36032
rect 29546 36020 29552 36032
rect 29507 35992 29552 36020
rect 29546 35980 29552 35992
rect 29604 35980 29610 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 2774 35816 2780 35828
rect 2700 35788 2780 35816
rect 2700 35689 2728 35788
rect 2774 35776 2780 35788
rect 2832 35776 2838 35828
rect 4982 35816 4988 35828
rect 4943 35788 4988 35816
rect 4982 35776 4988 35788
rect 5040 35776 5046 35828
rect 21818 35816 21824 35828
rect 21779 35788 21824 35816
rect 21818 35776 21824 35788
rect 21876 35776 21882 35828
rect 29733 35819 29791 35825
rect 29733 35785 29745 35819
rect 29779 35816 29791 35819
rect 30374 35816 30380 35828
rect 29779 35788 30380 35816
rect 29779 35785 29791 35788
rect 29733 35779 29791 35785
rect 30374 35776 30380 35788
rect 30432 35776 30438 35828
rect 4706 35708 4712 35760
rect 4764 35748 4770 35760
rect 22094 35748 22100 35760
rect 4764 35720 16620 35748
rect 4764 35708 4770 35720
rect 2685 35683 2743 35689
rect 2685 35649 2697 35683
rect 2731 35649 2743 35683
rect 5166 35680 5172 35692
rect 5127 35652 5172 35680
rect 2685 35643 2743 35649
rect 5166 35640 5172 35652
rect 5224 35640 5230 35692
rect 13630 35640 13636 35692
rect 13688 35680 13694 35692
rect 13688 35652 13733 35680
rect 13688 35640 13694 35652
rect 2869 35615 2927 35621
rect 2869 35581 2881 35615
rect 2915 35612 2927 35615
rect 2958 35612 2964 35624
rect 2915 35584 2964 35612
rect 2915 35581 2927 35584
rect 2869 35575 2927 35581
rect 2958 35572 2964 35584
rect 3016 35572 3022 35624
rect 3142 35612 3148 35624
rect 3103 35584 3148 35612
rect 3142 35572 3148 35584
rect 3200 35612 3206 35624
rect 7282 35612 7288 35624
rect 3200 35584 6914 35612
rect 7243 35584 7288 35612
rect 3200 35572 3206 35584
rect 6886 35544 6914 35584
rect 7282 35572 7288 35584
rect 7340 35572 7346 35624
rect 7469 35615 7527 35621
rect 7469 35581 7481 35615
rect 7515 35612 7527 35615
rect 7558 35612 7564 35624
rect 7515 35584 7564 35612
rect 7515 35581 7527 35584
rect 7469 35575 7527 35581
rect 7558 35572 7564 35584
rect 7616 35572 7622 35624
rect 9125 35615 9183 35621
rect 9125 35581 9137 35615
rect 9171 35612 9183 35615
rect 11790 35612 11796 35624
rect 9171 35584 11796 35612
rect 9171 35581 9183 35584
rect 9125 35575 9183 35581
rect 9140 35544 9168 35575
rect 11790 35572 11796 35584
rect 11848 35572 11854 35624
rect 13446 35612 13452 35624
rect 13407 35584 13452 35612
rect 13446 35572 13452 35584
rect 13504 35572 13510 35624
rect 6886 35516 9168 35544
rect 16592 35544 16620 35720
rect 18156 35720 22100 35748
rect 16758 35680 16764 35692
rect 16719 35652 16764 35680
rect 16758 35640 16764 35652
rect 16816 35640 16822 35692
rect 16945 35615 17003 35621
rect 16945 35581 16957 35615
rect 16991 35612 17003 35615
rect 17126 35612 17132 35624
rect 16991 35584 17132 35612
rect 16991 35581 17003 35584
rect 16945 35575 17003 35581
rect 17126 35572 17132 35584
rect 17184 35572 17190 35624
rect 17221 35615 17279 35621
rect 17221 35581 17233 35615
rect 17267 35612 17279 35615
rect 18156 35612 18184 35720
rect 22094 35708 22100 35720
rect 22152 35708 22158 35760
rect 19334 35680 19340 35692
rect 19295 35652 19340 35680
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 21726 35640 21732 35692
rect 21784 35680 21790 35692
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 21784 35652 22017 35680
rect 21784 35640 21790 35652
rect 22005 35649 22017 35652
rect 22051 35649 22063 35683
rect 22462 35680 22468 35692
rect 22423 35652 22468 35680
rect 22005 35643 22063 35649
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 23474 35680 23480 35692
rect 23435 35652 23480 35680
rect 23474 35640 23480 35652
rect 23532 35640 23538 35692
rect 28442 35640 28448 35692
rect 28500 35680 28506 35692
rect 28822 35683 28880 35689
rect 28822 35680 28834 35683
rect 28500 35652 28834 35680
rect 28500 35640 28506 35652
rect 28822 35649 28834 35652
rect 28868 35649 28880 35683
rect 28822 35643 28880 35649
rect 29549 35683 29607 35689
rect 29549 35649 29561 35683
rect 29595 35680 29607 35683
rect 29638 35680 29644 35692
rect 29595 35652 29644 35680
rect 29595 35649 29607 35652
rect 29549 35643 29607 35649
rect 29638 35640 29644 35652
rect 29696 35640 29702 35692
rect 19058 35612 19064 35624
rect 17267 35584 18184 35612
rect 19019 35584 19064 35612
rect 17267 35581 17279 35584
rect 17221 35575 17279 35581
rect 17236 35544 17264 35575
rect 19058 35572 19064 35584
rect 19116 35572 19122 35624
rect 23661 35615 23719 35621
rect 23661 35612 23673 35615
rect 22664 35584 23673 35612
rect 22664 35553 22692 35584
rect 23661 35581 23673 35584
rect 23707 35581 23719 35615
rect 23661 35575 23719 35581
rect 23842 35572 23848 35624
rect 23900 35612 23906 35624
rect 23937 35615 23995 35621
rect 23937 35612 23949 35615
rect 23900 35584 23949 35612
rect 23900 35572 23906 35584
rect 23937 35581 23949 35584
rect 23983 35581 23995 35615
rect 23937 35575 23995 35581
rect 29089 35615 29147 35621
rect 29089 35581 29101 35615
rect 29135 35612 29147 35615
rect 30926 35612 30932 35624
rect 29135 35584 30932 35612
rect 29135 35581 29147 35584
rect 29089 35575 29147 35581
rect 30926 35572 30932 35584
rect 30984 35612 30990 35624
rect 32582 35612 32588 35624
rect 30984 35584 32588 35612
rect 30984 35572 30990 35584
rect 32582 35572 32588 35584
rect 32640 35572 32646 35624
rect 16592 35516 17264 35544
rect 22649 35547 22707 35553
rect 22649 35513 22661 35547
rect 22695 35513 22707 35547
rect 22649 35507 22707 35513
rect 10965 35479 11023 35485
rect 10965 35445 10977 35479
rect 11011 35476 11023 35479
rect 13538 35476 13544 35488
rect 11011 35448 13544 35476
rect 11011 35445 11023 35448
rect 10965 35439 11023 35445
rect 13538 35436 13544 35448
rect 13596 35436 13602 35488
rect 15470 35476 15476 35488
rect 15431 35448 15476 35476
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 25961 35479 26019 35485
rect 25961 35445 25973 35479
rect 26007 35476 26019 35479
rect 26234 35476 26240 35488
rect 26007 35448 26240 35476
rect 26007 35445 26019 35448
rect 25961 35439 26019 35445
rect 26234 35436 26240 35448
rect 26292 35436 26298 35488
rect 27706 35476 27712 35488
rect 27667 35448 27712 35476
rect 27706 35436 27712 35448
rect 27764 35436 27770 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 7282 35232 7288 35284
rect 7340 35272 7346 35284
rect 7377 35275 7435 35281
rect 7377 35272 7389 35275
rect 7340 35244 7389 35272
rect 7340 35232 7346 35244
rect 7377 35241 7389 35244
rect 7423 35241 7435 35275
rect 7377 35235 7435 35241
rect 19058 35232 19064 35284
rect 19116 35272 19122 35284
rect 19429 35275 19487 35281
rect 19429 35272 19441 35275
rect 19116 35244 19441 35272
rect 19116 35232 19122 35244
rect 19429 35241 19441 35244
rect 19475 35241 19487 35275
rect 19429 35235 19487 35241
rect 19518 35232 19524 35284
rect 19576 35272 19582 35284
rect 19613 35275 19671 35281
rect 19613 35272 19625 35275
rect 19576 35244 19625 35272
rect 19576 35232 19582 35244
rect 19613 35241 19625 35244
rect 19659 35272 19671 35275
rect 20533 35275 20591 35281
rect 20533 35272 20545 35275
rect 19659 35244 20545 35272
rect 19659 35241 19671 35244
rect 19613 35235 19671 35241
rect 20533 35241 20545 35244
rect 20579 35272 20591 35275
rect 21269 35275 21327 35281
rect 21269 35272 21281 35275
rect 20579 35244 21281 35272
rect 20579 35241 20591 35244
rect 20533 35235 20591 35241
rect 21269 35241 21281 35244
rect 21315 35241 21327 35275
rect 21726 35272 21732 35284
rect 21687 35244 21732 35272
rect 21269 35235 21327 35241
rect 21726 35232 21732 35244
rect 21784 35232 21790 35284
rect 22370 35272 22376 35284
rect 22331 35244 22376 35272
rect 22370 35232 22376 35244
rect 22428 35232 22434 35284
rect 28442 35272 28448 35284
rect 28403 35244 28448 35272
rect 28442 35232 28448 35244
rect 28500 35232 28506 35284
rect 6914 35164 6920 35216
rect 6972 35204 6978 35216
rect 20349 35207 20407 35213
rect 20349 35204 20361 35207
rect 6972 35176 16896 35204
rect 6972 35164 6978 35176
rect 2866 35096 2872 35148
rect 2924 35136 2930 35148
rect 2961 35139 3019 35145
rect 2961 35136 2973 35139
rect 2924 35108 2973 35136
rect 2924 35096 2930 35108
rect 2961 35105 2973 35108
rect 3007 35105 3019 35139
rect 4614 35136 4620 35148
rect 4575 35108 4620 35136
rect 2961 35099 3019 35105
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 5534 35136 5540 35148
rect 5495 35108 5540 35136
rect 5534 35096 5540 35108
rect 5592 35096 5598 35148
rect 8938 35136 8944 35148
rect 8899 35108 8944 35136
rect 8938 35096 8944 35108
rect 8996 35096 9002 35148
rect 9416 35145 9444 35176
rect 16868 35148 16896 35176
rect 18708 35176 20361 35204
rect 9401 35139 9459 35145
rect 9401 35105 9413 35139
rect 9447 35105 9459 35139
rect 11790 35136 11796 35148
rect 11751 35108 11796 35136
rect 9401 35099 9459 35105
rect 11790 35096 11796 35108
rect 11848 35096 11854 35148
rect 13538 35136 13544 35148
rect 13499 35108 13544 35136
rect 13538 35096 13544 35108
rect 13596 35096 13602 35148
rect 14366 35136 14372 35148
rect 14327 35108 14372 35136
rect 14366 35096 14372 35108
rect 14424 35096 14430 35148
rect 15470 35136 15476 35148
rect 15431 35108 15476 35136
rect 15470 35096 15476 35108
rect 15528 35096 15534 35148
rect 16850 35136 16856 35148
rect 16811 35108 16856 35136
rect 16850 35096 16856 35108
rect 16908 35096 16914 35148
rect 18414 35136 18420 35148
rect 18375 35108 18420 35136
rect 18414 35096 18420 35108
rect 18472 35096 18478 35148
rect 18708 35145 18736 35176
rect 20349 35173 20361 35176
rect 20395 35173 20407 35207
rect 20806 35204 20812 35216
rect 20349 35167 20407 35173
rect 20640 35176 20812 35204
rect 20640 35145 20668 35176
rect 20806 35164 20812 35176
rect 20864 35204 20870 35216
rect 20864 35176 21404 35204
rect 20864 35164 20870 35176
rect 21376 35145 21404 35176
rect 18693 35139 18751 35145
rect 18693 35105 18705 35139
rect 18739 35105 18751 35139
rect 18693 35099 18751 35105
rect 19797 35139 19855 35145
rect 19797 35105 19809 35139
rect 19843 35136 19855 35139
rect 20625 35139 20683 35145
rect 20625 35136 20637 35139
rect 19843 35108 20637 35136
rect 19843 35105 19855 35108
rect 19797 35099 19855 35105
rect 20625 35105 20637 35108
rect 20671 35105 20683 35139
rect 20625 35099 20683 35105
rect 21361 35139 21419 35145
rect 21361 35105 21373 35139
rect 21407 35105 21419 35139
rect 21361 35099 21419 35105
rect 26234 35096 26240 35148
rect 26292 35136 26298 35148
rect 26292 35108 26337 35136
rect 26292 35096 26298 35108
rect 3237 35071 3295 35077
rect 3237 35037 3249 35071
rect 3283 35037 3295 35071
rect 3970 35068 3976 35080
rect 3931 35040 3976 35068
rect 3237 35031 3295 35037
rect 3252 35000 3280 35031
rect 3970 35028 3976 35040
rect 4028 35028 4034 35080
rect 14093 35071 14151 35077
rect 14093 35037 14105 35071
rect 14139 35068 14151 35071
rect 14182 35068 14188 35080
rect 14139 35040 14188 35068
rect 14139 35037 14151 35040
rect 14093 35031 14151 35037
rect 14182 35028 14188 35040
rect 14240 35028 14246 35080
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35068 19671 35071
rect 19978 35068 19984 35080
rect 19659 35040 19984 35068
rect 19659 35037 19671 35040
rect 19613 35031 19671 35037
rect 19978 35028 19984 35040
rect 20036 35068 20042 35080
rect 20533 35071 20591 35077
rect 20533 35068 20545 35071
rect 20036 35040 20545 35068
rect 20036 35028 20042 35040
rect 20533 35037 20545 35040
rect 20579 35068 20591 35071
rect 21545 35071 21603 35077
rect 21545 35068 21557 35071
rect 20579 35040 21557 35068
rect 20579 35037 20591 35040
rect 20533 35031 20591 35037
rect 21545 35037 21557 35040
rect 21591 35037 21603 35071
rect 22186 35068 22192 35080
rect 22147 35040 22192 35068
rect 21545 35031 21603 35037
rect 22186 35028 22192 35040
rect 22244 35028 22250 35080
rect 28261 35071 28319 35077
rect 28261 35037 28273 35071
rect 28307 35068 28319 35071
rect 28350 35068 28356 35080
rect 28307 35040 28356 35068
rect 28307 35037 28319 35040
rect 28261 35031 28319 35037
rect 28350 35028 28356 35040
rect 28408 35028 28414 35080
rect 4614 35000 4620 35012
rect 3252 34972 4620 35000
rect 4614 34960 4620 34972
rect 4672 34960 4678 35012
rect 4801 35003 4859 35009
rect 4801 34969 4813 35003
rect 4847 34969 4859 35003
rect 4801 34963 4859 34969
rect 4157 34935 4215 34941
rect 4157 34901 4169 34935
rect 4203 34932 4215 34935
rect 4816 34932 4844 34963
rect 8570 34960 8576 35012
rect 8628 35000 8634 35012
rect 9125 35003 9183 35009
rect 9125 35000 9137 35003
rect 8628 34972 9137 35000
rect 8628 34960 8634 34972
rect 9125 34969 9137 34972
rect 9171 34969 9183 35003
rect 9125 34963 9183 34969
rect 13262 34960 13268 35012
rect 13320 35000 13326 35012
rect 13357 35003 13415 35009
rect 13357 35000 13369 35003
rect 13320 34972 13369 35000
rect 13320 34960 13326 34972
rect 13357 34969 13369 34972
rect 13403 34969 13415 35003
rect 15654 35000 15660 35012
rect 15615 34972 15660 35000
rect 13357 34963 13415 34969
rect 15654 34960 15660 34972
rect 15712 34960 15718 35012
rect 19889 35003 19947 35009
rect 19889 34969 19901 35003
rect 19935 34969 19947 35003
rect 19889 34963 19947 34969
rect 4203 34904 4844 34932
rect 19904 34932 19932 34963
rect 20714 34960 20720 35012
rect 20772 35000 20778 35012
rect 20809 35003 20867 35009
rect 20809 35000 20821 35003
rect 20772 34972 20821 35000
rect 20772 34960 20778 34972
rect 20809 34969 20821 34972
rect 20855 35000 20867 35003
rect 21269 35003 21327 35009
rect 21269 35000 21281 35003
rect 20855 34972 21281 35000
rect 20855 34969 20867 34972
rect 20809 34963 20867 34969
rect 21269 34969 21281 34972
rect 21315 34969 21327 35003
rect 21269 34963 21327 34969
rect 23842 34960 23848 35012
rect 23900 35000 23906 35012
rect 24397 35003 24455 35009
rect 24397 35000 24409 35003
rect 23900 34972 24409 35000
rect 23900 34960 23906 34972
rect 24397 34969 24409 34972
rect 24443 34969 24455 35003
rect 24397 34963 24455 34969
rect 25038 34960 25044 35012
rect 25096 35000 25102 35012
rect 26053 35003 26111 35009
rect 26053 35000 26065 35003
rect 25096 34972 26065 35000
rect 25096 34960 25102 34972
rect 26053 34969 26065 34972
rect 26099 34969 26111 35003
rect 26053 34963 26111 34969
rect 20732 34932 20760 34960
rect 19904 34904 20760 34932
rect 4203 34901 4215 34904
rect 4157 34895 4215 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 3970 34688 3976 34740
rect 4028 34728 4034 34740
rect 4709 34731 4767 34737
rect 4709 34728 4721 34731
rect 4028 34700 4721 34728
rect 4028 34688 4034 34700
rect 4709 34697 4721 34700
rect 4755 34697 4767 34731
rect 7558 34728 7564 34740
rect 7519 34700 7564 34728
rect 4709 34691 4767 34697
rect 7558 34688 7564 34700
rect 7616 34688 7622 34740
rect 8570 34728 8576 34740
rect 8531 34700 8576 34728
rect 8570 34688 8576 34700
rect 8628 34688 8634 34740
rect 15565 34731 15623 34737
rect 15565 34697 15577 34731
rect 15611 34728 15623 34731
rect 15654 34728 15660 34740
rect 15611 34700 15660 34728
rect 15611 34697 15623 34700
rect 15565 34691 15623 34697
rect 15654 34688 15660 34700
rect 15712 34688 15718 34740
rect 17589 34731 17647 34737
rect 17589 34697 17601 34731
rect 17635 34697 17647 34731
rect 17589 34691 17647 34697
rect 21177 34731 21235 34737
rect 21177 34697 21189 34731
rect 21223 34728 21235 34731
rect 22462 34728 22468 34740
rect 21223 34700 22468 34728
rect 21223 34697 21235 34700
rect 21177 34691 21235 34697
rect 3418 34620 3424 34672
rect 3476 34660 3482 34672
rect 10873 34663 10931 34669
rect 10873 34660 10885 34663
rect 3476 34632 10885 34660
rect 3476 34620 3482 34632
rect 10873 34629 10885 34632
rect 10919 34660 10931 34663
rect 17604 34660 17632 34691
rect 22462 34688 22468 34700
rect 22520 34688 22526 34740
rect 28350 34728 28356 34740
rect 28311 34700 28356 34728
rect 28350 34688 28356 34700
rect 28408 34688 28414 34740
rect 29638 34728 29644 34740
rect 29599 34700 29644 34728
rect 29638 34688 29644 34700
rect 29696 34688 29702 34740
rect 18233 34663 18291 34669
rect 18233 34660 18245 34663
rect 10919 34632 17264 34660
rect 17604 34632 18245 34660
rect 10919 34629 10931 34632
rect 10873 34623 10931 34629
rect 2958 34552 2964 34604
rect 3016 34592 3022 34604
rect 3973 34595 4031 34601
rect 3973 34592 3985 34595
rect 3016 34564 3985 34592
rect 3016 34552 3022 34564
rect 3973 34561 3985 34564
rect 4019 34561 4031 34595
rect 4890 34592 4896 34604
rect 4851 34564 4896 34592
rect 3973 34555 4031 34561
rect 4890 34552 4896 34564
rect 4948 34552 4954 34604
rect 5169 34595 5227 34601
rect 5169 34561 5181 34595
rect 5215 34592 5227 34595
rect 5718 34592 5724 34604
rect 5215 34564 5724 34592
rect 5215 34561 5227 34564
rect 5169 34555 5227 34561
rect 5718 34552 5724 34564
rect 5776 34552 5782 34604
rect 7374 34592 7380 34604
rect 7335 34564 7380 34592
rect 7374 34552 7380 34564
rect 7432 34552 7438 34604
rect 8386 34592 8392 34604
rect 8347 34564 8392 34592
rect 8386 34552 8392 34564
rect 8444 34552 8450 34604
rect 13262 34592 13268 34604
rect 13223 34564 13268 34592
rect 13262 34552 13268 34564
rect 13320 34552 13326 34604
rect 13446 34552 13452 34604
rect 13504 34592 13510 34604
rect 14553 34595 14611 34601
rect 14553 34592 14565 34595
rect 13504 34564 14565 34592
rect 13504 34552 13510 34564
rect 14553 34561 14565 34564
rect 14599 34561 14611 34595
rect 15194 34592 15200 34604
rect 14553 34555 14611 34561
rect 14752 34564 15200 34592
rect 4062 34484 4068 34536
rect 4120 34524 4126 34536
rect 4249 34527 4307 34533
rect 4249 34524 4261 34527
rect 4120 34496 4261 34524
rect 4120 34484 4126 34496
rect 4249 34493 4261 34496
rect 4295 34493 4307 34527
rect 4982 34524 4988 34536
rect 4943 34496 4988 34524
rect 4249 34487 4307 34493
rect 4982 34484 4988 34496
rect 5040 34484 5046 34536
rect 9030 34524 9036 34536
rect 8991 34496 9036 34524
rect 9030 34484 9036 34496
rect 9088 34484 9094 34536
rect 9214 34524 9220 34536
rect 9175 34496 9220 34524
rect 9214 34484 9220 34496
rect 9272 34484 9278 34536
rect 13541 34527 13599 34533
rect 13541 34493 13553 34527
rect 13587 34524 13599 34527
rect 14752 34524 14780 34564
rect 15194 34552 15200 34564
rect 15252 34552 15258 34604
rect 15378 34592 15384 34604
rect 15339 34564 15384 34592
rect 15378 34552 15384 34564
rect 15436 34552 15442 34604
rect 13587 34496 14780 34524
rect 14829 34527 14887 34533
rect 13587 34493 13599 34496
rect 13541 34487 13599 34493
rect 14829 34493 14841 34527
rect 14875 34524 14887 34527
rect 15654 34524 15660 34536
rect 14875 34496 15660 34524
rect 14875 34493 14887 34496
rect 14829 34487 14887 34493
rect 15654 34484 15660 34496
rect 15712 34484 15718 34536
rect 17236 34524 17264 34632
rect 18233 34629 18245 34632
rect 18279 34629 18291 34663
rect 18233 34623 18291 34629
rect 19978 34620 19984 34672
rect 20036 34660 20042 34672
rect 20036 34632 21036 34660
rect 20036 34620 20042 34632
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34592 17463 34595
rect 17954 34592 17960 34604
rect 17451 34564 17960 34592
rect 17451 34561 17463 34564
rect 17405 34555 17463 34561
rect 17954 34552 17960 34564
rect 18012 34552 18018 34604
rect 20714 34592 20720 34604
rect 20675 34564 20720 34592
rect 20714 34552 20720 34564
rect 20772 34552 20778 34604
rect 21008 34601 21036 34632
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34561 21051 34595
rect 20993 34555 21051 34561
rect 23845 34595 23903 34601
rect 23845 34561 23857 34595
rect 23891 34592 23903 34595
rect 25038 34592 25044 34604
rect 23891 34564 25044 34592
rect 23891 34561 23903 34564
rect 23845 34555 23903 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25133 34595 25191 34601
rect 25133 34561 25145 34595
rect 25179 34592 25191 34595
rect 25590 34592 25596 34604
rect 25179 34564 25596 34592
rect 25179 34561 25191 34564
rect 25133 34555 25191 34561
rect 25590 34552 25596 34564
rect 25648 34552 25654 34604
rect 28534 34592 28540 34604
rect 28495 34564 28540 34592
rect 28534 34552 28540 34564
rect 28592 34552 28598 34604
rect 29454 34592 29460 34604
rect 29415 34564 29460 34592
rect 29454 34552 29460 34564
rect 29512 34552 29518 34604
rect 31294 34592 31300 34604
rect 31255 34564 31300 34592
rect 31294 34552 31300 34564
rect 31352 34552 31358 34604
rect 31481 34595 31539 34601
rect 31481 34561 31493 34595
rect 31527 34592 31539 34595
rect 32125 34595 32183 34601
rect 32125 34592 32137 34595
rect 31527 34564 32137 34592
rect 31527 34561 31539 34564
rect 31481 34555 31539 34561
rect 32125 34561 32137 34564
rect 32171 34561 32183 34595
rect 32125 34555 32183 34561
rect 18046 34524 18052 34536
rect 17236 34496 17908 34524
rect 18007 34496 18052 34524
rect 17880 34456 17908 34496
rect 18046 34484 18052 34496
rect 18104 34484 18110 34536
rect 18509 34527 18567 34533
rect 18509 34524 18521 34527
rect 18156 34496 18521 34524
rect 18156 34456 18184 34496
rect 18509 34493 18521 34496
rect 18555 34524 18567 34527
rect 19242 34524 19248 34536
rect 18555 34496 19248 34524
rect 18555 34493 18567 34496
rect 18509 34487 18567 34493
rect 19242 34484 19248 34496
rect 19300 34484 19306 34536
rect 20806 34524 20812 34536
rect 20767 34496 20812 34524
rect 20806 34484 20812 34496
rect 20864 34484 20870 34536
rect 23014 34484 23020 34536
rect 23072 34524 23078 34536
rect 23569 34527 23627 34533
rect 23569 34524 23581 34527
rect 23072 34496 23581 34524
rect 23072 34484 23078 34496
rect 23569 34493 23581 34496
rect 23615 34493 23627 34527
rect 23569 34487 23627 34493
rect 24026 34484 24032 34536
rect 24084 34524 24090 34536
rect 24857 34527 24915 34533
rect 24857 34524 24869 34527
rect 24084 34496 24869 34524
rect 24084 34484 24090 34496
rect 24857 34493 24869 34496
rect 24903 34493 24915 34527
rect 24857 34487 24915 34493
rect 28721 34527 28779 34533
rect 28721 34493 28733 34527
rect 28767 34524 28779 34527
rect 29273 34527 29331 34533
rect 29273 34524 29285 34527
rect 28767 34496 29285 34524
rect 28767 34493 28779 34496
rect 28721 34487 28779 34493
rect 29273 34493 29285 34496
rect 29319 34524 29331 34527
rect 31113 34527 31171 34533
rect 31113 34524 31125 34527
rect 29319 34496 31125 34524
rect 29319 34493 29331 34496
rect 29273 34487 29331 34493
rect 31113 34493 31125 34496
rect 31159 34524 31171 34527
rect 32030 34524 32036 34536
rect 31159 34496 32036 34524
rect 31159 34493 31171 34496
rect 31113 34487 31171 34493
rect 32030 34484 32036 34496
rect 32088 34484 32094 34536
rect 17880 34428 18184 34456
rect 4706 34348 4712 34400
rect 4764 34388 4770 34400
rect 4893 34391 4951 34397
rect 4893 34388 4905 34391
rect 4764 34360 4905 34388
rect 4764 34348 4770 34360
rect 4893 34357 4905 34360
rect 4939 34388 4951 34391
rect 5534 34388 5540 34400
rect 4939 34360 5540 34388
rect 4939 34357 4951 34360
rect 4893 34351 4951 34357
rect 5534 34348 5540 34360
rect 5592 34348 5598 34400
rect 5718 34388 5724 34400
rect 5679 34360 5724 34388
rect 5718 34348 5724 34360
rect 5776 34348 5782 34400
rect 19334 34348 19340 34400
rect 19392 34388 19398 34400
rect 20346 34388 20352 34400
rect 19392 34360 20352 34388
rect 19392 34348 19398 34360
rect 20346 34348 20352 34360
rect 20404 34388 20410 34400
rect 20717 34391 20775 34397
rect 20717 34388 20729 34391
rect 20404 34360 20729 34388
rect 20404 34348 20410 34360
rect 20717 34357 20729 34360
rect 20763 34357 20775 34391
rect 32306 34388 32312 34400
rect 32267 34360 32312 34388
rect 20717 34351 20775 34357
rect 32306 34348 32312 34360
rect 32364 34348 32370 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 4706 34184 4712 34196
rect 4667 34156 4712 34184
rect 4706 34144 4712 34156
rect 4764 34144 4770 34196
rect 4893 34187 4951 34193
rect 4893 34153 4905 34187
rect 4939 34184 4951 34187
rect 5166 34184 5172 34196
rect 4939 34156 5172 34184
rect 4939 34153 4951 34156
rect 4893 34147 4951 34153
rect 5166 34144 5172 34156
rect 5224 34144 5230 34196
rect 5534 34184 5540 34196
rect 5495 34156 5540 34184
rect 5534 34144 5540 34156
rect 5592 34144 5598 34196
rect 9125 34187 9183 34193
rect 9125 34153 9137 34187
rect 9171 34184 9183 34187
rect 9214 34184 9220 34196
rect 9171 34156 9220 34184
rect 9171 34153 9183 34156
rect 9125 34147 9183 34153
rect 9214 34144 9220 34156
rect 9272 34144 9278 34196
rect 9582 34184 9588 34196
rect 9543 34156 9588 34184
rect 9582 34144 9588 34156
rect 9640 34144 9646 34196
rect 15654 34184 15660 34196
rect 15615 34156 15660 34184
rect 15654 34144 15660 34156
rect 15712 34144 15718 34196
rect 16117 34187 16175 34193
rect 16117 34153 16129 34187
rect 16163 34184 16175 34187
rect 16390 34184 16396 34196
rect 16163 34156 16396 34184
rect 16163 34153 16175 34156
rect 16117 34147 16175 34153
rect 16390 34144 16396 34156
rect 16448 34144 16454 34196
rect 18417 34187 18475 34193
rect 18417 34153 18429 34187
rect 18463 34184 18475 34187
rect 19334 34184 19340 34196
rect 18463 34156 19340 34184
rect 18463 34153 18475 34156
rect 18417 34147 18475 34153
rect 19334 34144 19340 34156
rect 19392 34144 19398 34196
rect 4614 34076 4620 34128
rect 4672 34116 4678 34128
rect 5353 34119 5411 34125
rect 5353 34116 5365 34119
rect 4672 34088 5365 34116
rect 4672 34076 4678 34088
rect 5353 34085 5365 34088
rect 5399 34085 5411 34119
rect 5353 34079 5411 34085
rect 17954 34076 17960 34128
rect 18012 34116 18018 34128
rect 18601 34119 18659 34125
rect 18601 34116 18613 34119
rect 18012 34088 18613 34116
rect 18012 34076 18018 34088
rect 18601 34085 18613 34088
rect 18647 34085 18659 34119
rect 18601 34079 18659 34085
rect 4982 34048 4988 34060
rect 4632 34020 4988 34048
rect 4632 33992 4660 34020
rect 4982 34008 4988 34020
rect 5040 34048 5046 34060
rect 5629 34051 5687 34057
rect 5629 34048 5641 34051
rect 5040 34020 5641 34048
rect 5040 34008 5046 34020
rect 5629 34017 5641 34020
rect 5675 34017 5687 34051
rect 16022 34048 16028 34060
rect 15983 34020 16028 34048
rect 5629 34011 5687 34017
rect 16022 34008 16028 34020
rect 16080 34008 16086 34060
rect 26326 34048 26332 34060
rect 26287 34020 26332 34048
rect 26326 34008 26332 34020
rect 26384 34048 26390 34060
rect 27246 34048 27252 34060
rect 26384 34020 27252 34048
rect 26384 34008 26390 34020
rect 27246 34008 27252 34020
rect 27304 34008 27310 34060
rect 32582 34048 32588 34060
rect 32543 34020 32588 34048
rect 32582 34008 32588 34020
rect 32640 34008 32646 34060
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 2406 33940 2412 33992
rect 2464 33980 2470 33992
rect 2501 33983 2559 33989
rect 2501 33980 2513 33983
rect 2464 33952 2513 33980
rect 2464 33940 2470 33952
rect 2501 33949 2513 33952
rect 2547 33949 2559 33983
rect 3970 33980 3976 33992
rect 3931 33952 3976 33980
rect 2501 33943 2559 33949
rect 3970 33940 3976 33952
rect 4028 33940 4034 33992
rect 4614 33980 4620 33992
rect 4575 33952 4620 33980
rect 4614 33940 4620 33952
rect 4672 33940 4678 33992
rect 4709 33983 4767 33989
rect 4709 33949 4721 33983
rect 4755 33980 4767 33983
rect 4890 33980 4896 33992
rect 4755 33952 4896 33980
rect 4755 33949 4767 33952
rect 4709 33943 4767 33949
rect 4890 33940 4896 33952
rect 4948 33980 4954 33992
rect 5537 33983 5595 33989
rect 5537 33980 5549 33983
rect 4948 33952 5549 33980
rect 4948 33940 4954 33952
rect 5537 33949 5549 33952
rect 5583 33949 5595 33983
rect 8938 33980 8944 33992
rect 8899 33952 8944 33980
rect 5537 33943 5595 33949
rect 8938 33940 8944 33952
rect 8996 33940 9002 33992
rect 9766 33980 9772 33992
rect 9727 33952 9772 33980
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 12713 33983 12771 33989
rect 12713 33949 12725 33983
rect 12759 33980 12771 33983
rect 14274 33980 14280 33992
rect 12759 33952 14280 33980
rect 12759 33949 12771 33952
rect 12713 33943 12771 33949
rect 14274 33940 14280 33952
rect 14332 33940 14338 33992
rect 15838 33980 15844 33992
rect 15799 33952 15844 33980
rect 15838 33940 15844 33952
rect 15896 33940 15902 33992
rect 18322 33980 18328 33992
rect 18283 33952 18328 33980
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 18417 33983 18475 33989
rect 18417 33949 18429 33983
rect 18463 33980 18475 33983
rect 19978 33980 19984 33992
rect 18463 33952 19984 33980
rect 18463 33949 18475 33952
rect 18417 33943 18475 33949
rect 19978 33940 19984 33952
rect 20036 33940 20042 33992
rect 25406 33980 25412 33992
rect 25367 33952 25412 33980
rect 25406 33940 25412 33952
rect 25464 33940 25470 33992
rect 32306 33940 32312 33992
rect 32364 33989 32370 33992
rect 32364 33980 32376 33989
rect 37461 33983 37519 33989
rect 32364 33952 32409 33980
rect 32364 33943 32376 33952
rect 37461 33949 37473 33983
rect 37507 33980 37519 33983
rect 38102 33980 38108 33992
rect 37507 33952 38108 33980
rect 37507 33949 37519 33952
rect 37461 33943 37519 33949
rect 32364 33940 32370 33943
rect 38102 33940 38108 33952
rect 38160 33940 38166 33992
rect 4433 33915 4491 33921
rect 4433 33881 4445 33915
rect 4479 33912 4491 33915
rect 5813 33915 5871 33921
rect 5813 33912 5825 33915
rect 4479 33884 5825 33912
rect 4479 33881 4491 33884
rect 4433 33875 4491 33881
rect 5813 33881 5825 33884
rect 5859 33881 5871 33915
rect 16114 33912 16120 33924
rect 16027 33884 16120 33912
rect 5813 33875 5871 33881
rect 1581 33847 1639 33853
rect 1581 33813 1593 33847
rect 1627 33844 1639 33847
rect 2498 33844 2504 33856
rect 1627 33816 2504 33844
rect 1627 33813 1639 33816
rect 1581 33807 1639 33813
rect 2498 33804 2504 33816
rect 2556 33804 2562 33856
rect 2590 33804 2596 33856
rect 2648 33844 2654 33856
rect 3789 33847 3847 33853
rect 3789 33844 3801 33847
rect 2648 33816 3801 33844
rect 2648 33804 2654 33816
rect 3789 33813 3801 33816
rect 3835 33813 3847 33847
rect 3789 33807 3847 33813
rect 5718 33804 5724 33856
rect 5776 33844 5782 33856
rect 5828 33844 5856 33875
rect 16114 33872 16120 33884
rect 16172 33912 16178 33924
rect 18141 33915 18199 33921
rect 18141 33912 18153 33915
rect 16172 33884 18153 33912
rect 16172 33872 16178 33884
rect 18141 33881 18153 33884
rect 18187 33881 18199 33915
rect 25590 33912 25596 33924
rect 25551 33884 25596 33912
rect 18141 33875 18199 33881
rect 25590 33872 25596 33884
rect 25648 33872 25654 33924
rect 28626 33872 28632 33924
rect 28684 33912 28690 33924
rect 28997 33915 29055 33921
rect 28997 33912 29009 33915
rect 28684 33884 29009 33912
rect 28684 33872 28690 33884
rect 28997 33881 29009 33884
rect 29043 33912 29055 33915
rect 29043 33884 30512 33912
rect 29043 33881 29055 33884
rect 28997 33875 29055 33881
rect 6365 33847 6423 33853
rect 6365 33844 6377 33847
rect 5776 33816 6377 33844
rect 5776 33804 5782 33816
rect 6365 33813 6377 33816
rect 6411 33844 6423 33847
rect 8754 33844 8760 33856
rect 6411 33816 8760 33844
rect 6411 33813 6423 33816
rect 6365 33807 6423 33813
rect 8754 33804 8760 33816
rect 8812 33804 8818 33856
rect 29641 33847 29699 33853
rect 29641 33813 29653 33847
rect 29687 33844 29699 33847
rect 29730 33844 29736 33856
rect 29687 33816 29736 33844
rect 29687 33813 29699 33816
rect 29641 33807 29699 33813
rect 29730 33804 29736 33816
rect 29788 33804 29794 33856
rect 30484 33853 30512 33884
rect 35342 33872 35348 33924
rect 35400 33912 35406 33924
rect 35400 33884 37964 33912
rect 35400 33872 35406 33884
rect 30469 33847 30527 33853
rect 30469 33813 30481 33847
rect 30515 33844 30527 33847
rect 30926 33844 30932 33856
rect 30515 33816 30932 33844
rect 30515 33813 30527 33816
rect 30469 33807 30527 33813
rect 30926 33804 30932 33816
rect 30984 33804 30990 33856
rect 31202 33844 31208 33856
rect 31163 33816 31208 33844
rect 31202 33804 31208 33816
rect 31260 33804 31266 33856
rect 37936 33853 37964 33884
rect 37921 33847 37979 33853
rect 37921 33813 37933 33847
rect 37967 33813 37979 33847
rect 37921 33807 37979 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 3970 33600 3976 33652
rect 4028 33640 4034 33652
rect 4709 33643 4767 33649
rect 4709 33640 4721 33643
rect 4028 33612 4721 33640
rect 4028 33600 4034 33612
rect 4709 33609 4721 33612
rect 4755 33609 4767 33643
rect 5718 33640 5724 33652
rect 5679 33612 5724 33640
rect 4709 33603 4767 33609
rect 5718 33600 5724 33612
rect 5776 33600 5782 33652
rect 23109 33643 23167 33649
rect 23109 33609 23121 33643
rect 23155 33640 23167 33643
rect 24026 33640 24032 33652
rect 23155 33612 24032 33640
rect 23155 33609 23167 33612
rect 23109 33603 23167 33609
rect 24026 33600 24032 33612
rect 24084 33600 24090 33652
rect 28261 33643 28319 33649
rect 28261 33609 28273 33643
rect 28307 33640 28319 33643
rect 28534 33640 28540 33652
rect 28307 33612 28540 33640
rect 28307 33609 28319 33612
rect 28261 33603 28319 33609
rect 28534 33600 28540 33612
rect 28592 33600 28598 33652
rect 29273 33643 29331 33649
rect 29273 33609 29285 33643
rect 29319 33640 29331 33643
rect 29454 33640 29460 33652
rect 29319 33612 29460 33640
rect 29319 33609 29331 33612
rect 29273 33603 29331 33609
rect 29454 33600 29460 33612
rect 29512 33600 29518 33652
rect 31110 33640 31116 33652
rect 31036 33612 31116 33640
rect 1394 33572 1400 33584
rect 1355 33544 1400 33572
rect 1394 33532 1400 33544
rect 1452 33532 1458 33584
rect 2590 33572 2596 33584
rect 2551 33544 2596 33572
rect 2590 33532 2596 33544
rect 2648 33532 2654 33584
rect 14093 33575 14151 33581
rect 14093 33541 14105 33575
rect 14139 33572 14151 33575
rect 14139 33544 15332 33572
rect 14139 33541 14151 33544
rect 14093 33535 14151 33541
rect 2406 33504 2412 33516
rect 2367 33476 2412 33504
rect 2406 33464 2412 33476
rect 2464 33464 2470 33516
rect 4893 33507 4951 33513
rect 4893 33473 4905 33507
rect 4939 33504 4951 33507
rect 4982 33504 4988 33516
rect 4939 33476 4988 33504
rect 4939 33473 4951 33476
rect 4893 33467 4951 33473
rect 4982 33464 4988 33476
rect 5040 33464 5046 33516
rect 5169 33507 5227 33513
rect 5169 33473 5181 33507
rect 5215 33504 5227 33507
rect 5258 33504 5264 33516
rect 5215 33476 5264 33504
rect 5215 33473 5227 33476
rect 5169 33467 5227 33473
rect 5258 33464 5264 33476
rect 5316 33464 5322 33516
rect 9030 33504 9036 33516
rect 8991 33476 9036 33504
rect 9030 33464 9036 33476
rect 9088 33464 9094 33516
rect 14274 33464 14280 33516
rect 14332 33504 14338 33516
rect 15304 33513 15332 33544
rect 20714 33532 20720 33584
rect 20772 33572 20778 33584
rect 22649 33575 22707 33581
rect 22649 33572 22661 33575
rect 20772 33544 22661 33572
rect 20772 33532 20778 33544
rect 22649 33541 22661 33544
rect 22695 33541 22707 33575
rect 22649 33535 22707 33541
rect 27706 33532 27712 33584
rect 27764 33572 27770 33584
rect 27764 33544 28580 33572
rect 27764 33532 27770 33544
rect 15289 33507 15347 33513
rect 14332 33476 14377 33504
rect 14332 33464 14338 33476
rect 15289 33473 15301 33507
rect 15335 33473 15347 33507
rect 15289 33467 15347 33473
rect 18046 33464 18052 33516
rect 18104 33504 18110 33516
rect 18141 33507 18199 33513
rect 18141 33504 18153 33507
rect 18104 33476 18153 33504
rect 18104 33464 18110 33476
rect 18141 33473 18153 33476
rect 18187 33473 18199 33507
rect 20346 33504 20352 33516
rect 20307 33476 20352 33504
rect 18141 33467 18199 33473
rect 20346 33464 20352 33476
rect 20404 33464 20410 33516
rect 22922 33504 22928 33516
rect 22883 33476 22928 33504
rect 22922 33464 22928 33476
rect 22980 33464 22986 33516
rect 25406 33504 25412 33516
rect 25367 33476 25412 33504
rect 25406 33464 25412 33476
rect 25464 33464 25470 33516
rect 28552 33513 28580 33544
rect 28626 33532 28632 33584
rect 28684 33572 28690 33584
rect 29546 33572 29552 33584
rect 28684 33544 28729 33572
rect 29507 33544 29552 33572
rect 28684 33532 28690 33544
rect 29546 33532 29552 33544
rect 29604 33532 29610 33584
rect 29641 33575 29699 33581
rect 29641 33541 29653 33575
rect 29687 33572 29699 33575
rect 30926 33572 30932 33584
rect 29687 33544 30932 33572
rect 29687 33541 29699 33544
rect 29641 33535 29699 33541
rect 30926 33532 30932 33544
rect 30984 33532 30990 33584
rect 31036 33581 31064 33612
rect 31110 33600 31116 33612
rect 31168 33600 31174 33652
rect 31294 33640 31300 33652
rect 31255 33612 31300 33640
rect 31294 33600 31300 33612
rect 31352 33600 31358 33652
rect 31021 33575 31079 33581
rect 31021 33541 31033 33575
rect 31067 33541 31079 33575
rect 31021 33535 31079 33541
rect 28445 33507 28503 33513
rect 28445 33473 28457 33507
rect 28491 33473 28503 33507
rect 28445 33467 28503 33473
rect 28537 33507 28595 33513
rect 28537 33473 28549 33507
rect 28583 33473 28595 33507
rect 28810 33504 28816 33516
rect 28771 33476 28816 33504
rect 28537 33467 28595 33473
rect 2866 33436 2872 33448
rect 2827 33408 2872 33436
rect 2866 33396 2872 33408
rect 2924 33396 2930 33448
rect 4614 33396 4620 33448
rect 4672 33436 4678 33448
rect 5077 33439 5135 33445
rect 5077 33436 5089 33439
rect 4672 33408 5089 33436
rect 4672 33396 4678 33408
rect 5077 33405 5089 33408
rect 5123 33436 5135 33439
rect 5350 33436 5356 33448
rect 5123 33408 5356 33436
rect 5123 33405 5135 33408
rect 5077 33399 5135 33405
rect 5350 33396 5356 33408
rect 5408 33396 5414 33448
rect 12434 33396 12440 33448
rect 12492 33436 12498 33448
rect 15565 33439 15623 33445
rect 12492 33408 12537 33436
rect 12492 33396 12498 33408
rect 15565 33405 15577 33439
rect 15611 33436 15623 33439
rect 16574 33436 16580 33448
rect 15611 33408 16580 33436
rect 15611 33405 15623 33408
rect 15565 33399 15623 33405
rect 16574 33396 16580 33408
rect 16632 33396 16638 33448
rect 20625 33439 20683 33445
rect 20625 33405 20637 33439
rect 20671 33405 20683 33439
rect 20625 33399 20683 33405
rect 2884 33368 2912 33396
rect 6086 33368 6092 33380
rect 2884 33340 6092 33368
rect 6086 33328 6092 33340
rect 6144 33328 6150 33380
rect 20346 33328 20352 33380
rect 20404 33368 20410 33380
rect 20640 33368 20668 33399
rect 20806 33396 20812 33448
rect 20864 33436 20870 33448
rect 22741 33439 22799 33445
rect 22741 33436 22753 33439
rect 20864 33408 22753 33436
rect 20864 33396 20870 33408
rect 22741 33405 22753 33408
rect 22787 33405 22799 33439
rect 22741 33399 22799 33405
rect 20404 33340 20668 33368
rect 28460 33368 28488 33467
rect 28810 33464 28816 33476
rect 28868 33464 28874 33516
rect 29454 33504 29460 33516
rect 29415 33476 29460 33504
rect 29454 33464 29460 33476
rect 29512 33464 29518 33516
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33473 29883 33507
rect 30742 33504 30748 33516
rect 30703 33476 30748 33504
rect 29825 33467 29883 33473
rect 28994 33396 29000 33448
rect 29052 33436 29058 33448
rect 29730 33436 29736 33448
rect 29052 33408 29736 33436
rect 29052 33396 29058 33408
rect 29730 33396 29736 33408
rect 29788 33436 29794 33448
rect 29840 33436 29868 33467
rect 30742 33464 30748 33476
rect 30800 33464 30806 33516
rect 31113 33507 31171 33513
rect 31113 33473 31125 33507
rect 31159 33504 31171 33507
rect 31159 33476 31248 33504
rect 31159 33473 31171 33476
rect 31113 33467 31171 33473
rect 29788 33408 29868 33436
rect 29788 33396 29794 33408
rect 29454 33368 29460 33380
rect 28460 33340 29460 33368
rect 20404 33328 20410 33340
rect 29454 33328 29460 33340
rect 29512 33368 29518 33380
rect 31220 33368 31248 33476
rect 32490 33368 32496 33380
rect 29512 33340 32496 33368
rect 29512 33328 29518 33340
rect 32490 33328 32496 33340
rect 32548 33328 32554 33380
rect 5169 33303 5227 33309
rect 5169 33269 5181 33303
rect 5215 33300 5227 33303
rect 5534 33300 5540 33312
rect 5215 33272 5540 33300
rect 5215 33269 5227 33272
rect 5169 33263 5227 33269
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 22830 33300 22836 33312
rect 22791 33272 22836 33300
rect 22830 33260 22836 33272
rect 22888 33260 22894 33312
rect 27801 33303 27859 33309
rect 27801 33269 27813 33303
rect 27847 33300 27859 33303
rect 28350 33300 28356 33312
rect 27847 33272 28356 33300
rect 27847 33269 27859 33272
rect 27801 33263 27859 33269
rect 28350 33260 28356 33272
rect 28408 33300 28414 33312
rect 28810 33300 28816 33312
rect 28408 33272 28816 33300
rect 28408 33260 28414 33272
rect 28810 33260 28816 33272
rect 28868 33260 28874 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 4062 33096 4068 33108
rect 4023 33068 4068 33096
rect 4062 33056 4068 33068
rect 4120 33056 4126 33108
rect 4525 33099 4583 33105
rect 4525 33065 4537 33099
rect 4571 33096 4583 33099
rect 5534 33096 5540 33108
rect 4571 33068 5540 33096
rect 4571 33065 4583 33068
rect 4525 33059 4583 33065
rect 5534 33056 5540 33068
rect 5592 33056 5598 33108
rect 8113 33099 8171 33105
rect 8113 33065 8125 33099
rect 8159 33065 8171 33099
rect 8386 33096 8392 33108
rect 8347 33068 8392 33096
rect 8113 33059 8171 33065
rect 8128 33028 8156 33059
rect 8386 33056 8392 33068
rect 8444 33056 8450 33108
rect 8938 33096 8944 33108
rect 8899 33068 8944 33096
rect 8938 33056 8944 33068
rect 8996 33056 9002 33108
rect 9125 33099 9183 33105
rect 9125 33065 9137 33099
rect 9171 33065 9183 33099
rect 9125 33059 9183 33065
rect 16117 33099 16175 33105
rect 16117 33065 16129 33099
rect 16163 33096 16175 33099
rect 16574 33096 16580 33108
rect 16163 33068 16436 33096
rect 16535 33068 16580 33096
rect 16163 33065 16175 33068
rect 16117 33059 16175 33065
rect 8202 33028 8208 33040
rect 8115 33000 8208 33028
rect 8202 32988 8208 33000
rect 8260 33028 8266 33040
rect 9140 33028 9168 33059
rect 16408 33040 16436 33068
rect 16574 33056 16580 33068
rect 16632 33056 16638 33108
rect 16761 33099 16819 33105
rect 16761 33065 16773 33099
rect 16807 33065 16819 33099
rect 19978 33096 19984 33108
rect 19939 33068 19984 33096
rect 16761 33059 16819 33065
rect 15657 33031 15715 33037
rect 15657 33028 15669 33031
rect 8260 33000 9168 33028
rect 14936 33000 15669 33028
rect 8260 32988 8266 33000
rect 4433 32963 4491 32969
rect 4433 32929 4445 32963
rect 4479 32960 4491 32963
rect 5350 32960 5356 32972
rect 4479 32932 5356 32960
rect 4479 32929 4491 32932
rect 4433 32923 4491 32929
rect 5350 32920 5356 32932
rect 5408 32920 5414 32972
rect 8113 32963 8171 32969
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8386 32960 8392 32972
rect 8159 32932 8392 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 8386 32920 8392 32932
rect 8444 32960 8450 32972
rect 9309 32963 9367 32969
rect 9309 32960 9321 32963
rect 8444 32932 9321 32960
rect 8444 32920 8450 32932
rect 9309 32929 9321 32932
rect 9355 32960 9367 32963
rect 14826 32960 14832 32972
rect 9355 32932 14832 32960
rect 9355 32929 9367 32932
rect 9309 32923 9367 32929
rect 14826 32920 14832 32932
rect 14884 32920 14890 32972
rect 14936 32969 14964 33000
rect 15657 32997 15669 33000
rect 15703 32997 15715 33031
rect 15657 32991 15715 32997
rect 15838 32988 15844 33040
rect 15896 33028 15902 33040
rect 16298 33028 16304 33040
rect 15896 33000 16304 33028
rect 15896 32988 15902 33000
rect 16298 32988 16304 33000
rect 16356 32988 16362 33040
rect 16390 32988 16396 33040
rect 16448 33028 16454 33040
rect 16776 33028 16804 33059
rect 19978 33056 19984 33068
rect 20036 33056 20042 33108
rect 20625 33099 20683 33105
rect 20625 33065 20637 33099
rect 20671 33096 20683 33099
rect 20806 33096 20812 33108
rect 20671 33068 20812 33096
rect 20671 33065 20683 33068
rect 20625 33059 20683 33065
rect 20806 33056 20812 33068
rect 20864 33056 20870 33108
rect 21913 33099 21971 33105
rect 21913 33065 21925 33099
rect 21959 33065 21971 33099
rect 21913 33059 21971 33065
rect 22097 33099 22155 33105
rect 22097 33065 22109 33099
rect 22143 33096 22155 33099
rect 22186 33096 22192 33108
rect 22143 33068 22192 33096
rect 22143 33065 22155 33068
rect 22097 33059 22155 33065
rect 21928 33028 21956 33059
rect 22186 33056 22192 33068
rect 22244 33056 22250 33108
rect 22557 33099 22615 33105
rect 22557 33065 22569 33099
rect 22603 33065 22615 33099
rect 23014 33096 23020 33108
rect 22975 33068 23020 33096
rect 22557 33059 22615 33065
rect 22002 33028 22008 33040
rect 16448 33000 16804 33028
rect 21915 33000 22008 33028
rect 16448 32988 16454 33000
rect 22002 32988 22008 33000
rect 22060 33028 22066 33040
rect 22572 33028 22600 33059
rect 23014 33056 23020 33068
rect 23072 33056 23078 33108
rect 22060 33000 22600 33028
rect 22060 32988 22066 33000
rect 14921 32963 14979 32969
rect 14921 32929 14933 32963
rect 14967 32929 14979 32963
rect 14921 32923 14979 32929
rect 4249 32895 4307 32901
rect 4249 32861 4261 32895
rect 4295 32892 4307 32895
rect 4982 32892 4988 32904
rect 4295 32864 4988 32892
rect 4295 32861 4307 32864
rect 4249 32855 4307 32861
rect 4982 32852 4988 32864
rect 5040 32852 5046 32904
rect 5626 32892 5632 32904
rect 5587 32864 5632 32892
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 8205 32895 8263 32901
rect 8205 32861 8217 32895
rect 8251 32892 8263 32895
rect 8478 32892 8484 32904
rect 8251 32864 8484 32892
rect 8251 32861 8263 32864
rect 8205 32855 8263 32861
rect 8478 32852 8484 32864
rect 8536 32892 8542 32904
rect 9125 32895 9183 32901
rect 9125 32892 9137 32895
rect 8536 32864 9137 32892
rect 8536 32852 8542 32864
rect 9125 32861 9137 32864
rect 9171 32861 9183 32895
rect 9125 32855 9183 32861
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32861 12771 32895
rect 12713 32855 12771 32861
rect 4525 32827 4583 32833
rect 4525 32793 4537 32827
rect 4571 32824 4583 32827
rect 5258 32824 5264 32836
rect 4571 32796 5264 32824
rect 4571 32793 4583 32796
rect 4525 32787 4583 32793
rect 5258 32784 5264 32796
rect 5316 32784 5322 32836
rect 7929 32827 7987 32833
rect 7929 32793 7941 32827
rect 7975 32824 7987 32827
rect 8110 32824 8116 32836
rect 7975 32796 8116 32824
rect 7975 32793 7987 32796
rect 7929 32787 7987 32793
rect 8110 32784 8116 32796
rect 8168 32824 8174 32836
rect 9401 32827 9459 32833
rect 9401 32824 9413 32827
rect 8168 32796 9413 32824
rect 8168 32784 8174 32796
rect 9401 32793 9413 32796
rect 9447 32793 9459 32827
rect 12728 32824 12756 32855
rect 14090 32852 14096 32904
rect 14148 32892 14154 32904
rect 15856 32901 15884 32988
rect 16022 32960 16028 32972
rect 15935 32932 16028 32960
rect 16022 32920 16028 32932
rect 16080 32960 16086 32972
rect 16945 32963 17003 32969
rect 16945 32960 16957 32963
rect 16080 32932 16957 32960
rect 16080 32920 16086 32932
rect 16945 32929 16957 32932
rect 16991 32960 17003 32963
rect 18322 32960 18328 32972
rect 16991 32932 18328 32960
rect 16991 32929 17003 32932
rect 16945 32923 17003 32929
rect 18322 32920 18328 32932
rect 18380 32920 18386 32972
rect 21726 32960 21732 32972
rect 19812 32932 20576 32960
rect 21687 32932 21732 32960
rect 14645 32895 14703 32901
rect 14645 32892 14657 32895
rect 14148 32864 14657 32892
rect 14148 32852 14154 32864
rect 14645 32861 14657 32864
rect 14691 32861 14703 32895
rect 14645 32855 14703 32861
rect 15841 32895 15899 32901
rect 15841 32861 15853 32895
rect 15887 32861 15899 32895
rect 16114 32892 16120 32904
rect 16075 32864 16120 32892
rect 15841 32855 15899 32861
rect 16114 32852 16120 32864
rect 16172 32852 16178 32904
rect 16298 32852 16304 32904
rect 16356 32892 16362 32904
rect 16761 32895 16819 32901
rect 16761 32892 16773 32895
rect 16356 32864 16773 32892
rect 16356 32852 16362 32864
rect 16761 32861 16773 32864
rect 16807 32892 16819 32895
rect 18966 32892 18972 32904
rect 16807 32864 18972 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 18966 32852 18972 32864
rect 19024 32852 19030 32904
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 19812 32901 19840 32932
rect 19797 32895 19855 32901
rect 19797 32892 19809 32895
rect 19208 32864 19809 32892
rect 19208 32852 19214 32864
rect 19797 32861 19809 32864
rect 19843 32861 19855 32895
rect 20438 32892 20444 32904
rect 20399 32864 20444 32892
rect 19797 32855 19855 32861
rect 20438 32852 20444 32864
rect 20496 32852 20502 32904
rect 20548 32892 20576 32932
rect 21726 32920 21732 32932
rect 21784 32960 21790 32972
rect 22649 32963 22707 32969
rect 22649 32960 22661 32963
rect 21784 32932 22661 32960
rect 21784 32920 21790 32932
rect 22649 32929 22661 32932
rect 22695 32929 22707 32963
rect 22649 32923 22707 32929
rect 27157 32963 27215 32969
rect 27157 32929 27169 32963
rect 27203 32960 27215 32963
rect 27706 32960 27712 32972
rect 27203 32932 27712 32960
rect 27203 32929 27215 32932
rect 27157 32923 27215 32929
rect 27706 32920 27712 32932
rect 27764 32920 27770 32972
rect 28350 32960 28356 32972
rect 28311 32932 28356 32960
rect 28350 32920 28356 32932
rect 28408 32920 28414 32972
rect 21913 32895 21971 32901
rect 20548 32864 21772 32892
rect 14274 32824 14280 32836
rect 12728 32796 14280 32824
rect 9401 32787 9459 32793
rect 9416 32756 9444 32787
rect 14274 32784 14280 32796
rect 14332 32784 14338 32836
rect 16132 32824 16160 32852
rect 16482 32824 16488 32836
rect 16132 32796 16488 32824
rect 16482 32784 16488 32796
rect 16540 32824 16546 32836
rect 17037 32827 17095 32833
rect 17037 32824 17049 32827
rect 16540 32796 17049 32824
rect 16540 32784 16546 32796
rect 17037 32793 17049 32796
rect 17083 32793 17095 32827
rect 21637 32827 21695 32833
rect 21637 32824 21649 32827
rect 17037 32787 17095 32793
rect 17144 32796 21649 32824
rect 17144 32756 17172 32796
rect 21637 32793 21649 32796
rect 21683 32793 21695 32827
rect 21744 32824 21772 32864
rect 21913 32861 21925 32895
rect 21959 32892 21971 32895
rect 22833 32895 22891 32901
rect 22833 32892 22845 32895
rect 21959 32864 22845 32892
rect 21959 32861 21971 32864
rect 21913 32855 21971 32861
rect 22833 32861 22845 32864
rect 22879 32892 22891 32895
rect 23290 32892 23296 32904
rect 22879 32864 23296 32892
rect 22879 32861 22891 32864
rect 22833 32855 22891 32861
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 24854 32892 24860 32904
rect 24815 32864 24860 32892
rect 24854 32852 24860 32864
rect 24912 32852 24918 32904
rect 22370 32824 22376 32836
rect 21744 32796 22376 32824
rect 21637 32787 21695 32793
rect 22370 32784 22376 32796
rect 22428 32784 22434 32836
rect 22557 32827 22615 32833
rect 22557 32793 22569 32827
rect 22603 32824 22615 32827
rect 23106 32824 23112 32836
rect 22603 32796 23112 32824
rect 22603 32793 22615 32796
rect 22557 32787 22615 32793
rect 23106 32784 23112 32796
rect 23164 32784 23170 32836
rect 25041 32827 25099 32833
rect 25041 32793 25053 32827
rect 25087 32824 25099 32827
rect 25314 32824 25320 32836
rect 25087 32796 25320 32824
rect 25087 32793 25099 32796
rect 25041 32787 25099 32793
rect 25314 32784 25320 32796
rect 25372 32784 25378 32836
rect 26694 32824 26700 32836
rect 26655 32796 26700 32824
rect 26694 32784 26700 32796
rect 26752 32784 26758 32836
rect 27338 32824 27344 32836
rect 27299 32796 27344 32824
rect 27338 32784 27344 32796
rect 27396 32784 27402 32836
rect 30009 32827 30067 32833
rect 30009 32793 30021 32827
rect 30055 32824 30067 32827
rect 31018 32824 31024 32836
rect 30055 32796 31024 32824
rect 30055 32793 30067 32796
rect 30009 32787 30067 32793
rect 31018 32784 31024 32796
rect 31076 32784 31082 32836
rect 9416 32728 17172 32756
rect 30653 32759 30711 32765
rect 30653 32725 30665 32759
rect 30699 32756 30711 32759
rect 30742 32756 30748 32768
rect 30699 32728 30748 32756
rect 30699 32725 30711 32728
rect 30653 32719 30711 32725
rect 30742 32716 30748 32728
rect 30800 32756 30806 32768
rect 31570 32756 31576 32768
rect 30800 32728 31576 32756
rect 30800 32716 30806 32728
rect 31570 32716 31576 32728
rect 31628 32716 31634 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 5350 32552 5356 32564
rect 5311 32524 5356 32552
rect 5350 32512 5356 32524
rect 5408 32512 5414 32564
rect 7374 32552 7380 32564
rect 7335 32524 7380 32552
rect 7374 32512 7380 32524
rect 7432 32512 7438 32564
rect 8665 32555 8723 32561
rect 8665 32521 8677 32555
rect 8711 32552 8723 32555
rect 9766 32552 9772 32564
rect 8711 32524 9772 32552
rect 8711 32521 8723 32524
rect 8665 32515 8723 32521
rect 9766 32512 9772 32524
rect 9824 32512 9830 32564
rect 16482 32512 16488 32564
rect 16540 32552 16546 32564
rect 17129 32555 17187 32561
rect 17129 32552 17141 32555
rect 16540 32524 17141 32552
rect 16540 32512 16546 32524
rect 17129 32521 17141 32524
rect 17175 32521 17187 32555
rect 18322 32552 18328 32564
rect 18283 32524 18328 32552
rect 17129 32515 17187 32521
rect 18322 32512 18328 32524
rect 18380 32512 18386 32564
rect 20714 32552 20720 32564
rect 20675 32524 20720 32552
rect 20714 32512 20720 32524
rect 20772 32512 20778 32564
rect 22002 32552 22008 32564
rect 21963 32524 22008 32552
rect 22002 32512 22008 32524
rect 22060 32512 22066 32564
rect 23477 32555 23535 32561
rect 23477 32521 23489 32555
rect 23523 32521 23535 32555
rect 25314 32552 25320 32564
rect 25275 32524 25320 32552
rect 23477 32515 23535 32521
rect 6917 32487 6975 32493
rect 6917 32453 6929 32487
rect 6963 32484 6975 32487
rect 7282 32484 7288 32496
rect 6963 32456 7288 32484
rect 6963 32453 6975 32456
rect 6917 32447 6975 32453
rect 7282 32444 7288 32456
rect 7340 32484 7346 32496
rect 8110 32484 8116 32496
rect 7340 32456 8116 32484
rect 7340 32444 7346 32456
rect 8110 32444 8116 32456
rect 8168 32484 8174 32496
rect 8205 32487 8263 32493
rect 8205 32484 8217 32487
rect 8168 32456 8217 32484
rect 8168 32444 8174 32456
rect 8205 32453 8217 32456
rect 8251 32453 8263 32487
rect 14090 32484 14096 32496
rect 14051 32456 14096 32484
rect 8205 32447 8263 32453
rect 14090 32444 14096 32456
rect 14148 32444 14154 32496
rect 14826 32444 14832 32496
rect 14884 32484 14890 32496
rect 21726 32484 21732 32496
rect 14884 32456 21732 32484
rect 14884 32444 14890 32456
rect 21726 32444 21732 32456
rect 21784 32444 21790 32496
rect 1394 32416 1400 32428
rect 1355 32388 1400 32416
rect 1394 32376 1400 32388
rect 1452 32416 1458 32428
rect 2041 32419 2099 32425
rect 2041 32416 2053 32419
rect 1452 32388 2053 32416
rect 1452 32376 1458 32388
rect 2041 32385 2053 32388
rect 2087 32385 2099 32419
rect 2041 32379 2099 32385
rect 4709 32419 4767 32425
rect 4709 32385 4721 32419
rect 4755 32416 4767 32419
rect 5166 32416 5172 32428
rect 4755 32388 5172 32416
rect 4755 32385 4767 32388
rect 4709 32379 4767 32385
rect 5166 32376 5172 32388
rect 5224 32376 5230 32428
rect 7193 32419 7251 32425
rect 7193 32385 7205 32419
rect 7239 32385 7251 32419
rect 8478 32416 8484 32428
rect 8391 32388 8484 32416
rect 7193 32379 7251 32385
rect 6270 32308 6276 32360
rect 6328 32348 6334 32360
rect 7009 32351 7067 32357
rect 7009 32348 7021 32351
rect 6328 32320 7021 32348
rect 6328 32308 6334 32320
rect 7009 32317 7021 32320
rect 7055 32317 7067 32351
rect 7009 32311 7067 32317
rect 6178 32240 6184 32292
rect 6236 32280 6242 32292
rect 7208 32280 7236 32379
rect 8478 32376 8484 32388
rect 8536 32376 8542 32428
rect 14274 32376 14280 32428
rect 14332 32416 14338 32428
rect 16945 32419 17003 32425
rect 14332 32388 14377 32416
rect 14332 32376 14338 32388
rect 16945 32385 16957 32419
rect 16991 32416 17003 32419
rect 17589 32419 17647 32425
rect 17589 32416 17601 32419
rect 16991 32388 17601 32416
rect 16991 32385 17003 32388
rect 16945 32379 17003 32385
rect 17589 32385 17601 32388
rect 17635 32416 17647 32419
rect 17770 32416 17776 32428
rect 17635 32388 17776 32416
rect 17635 32385 17647 32388
rect 17589 32379 17647 32385
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32385 18567 32419
rect 19150 32416 19156 32428
rect 19111 32388 19156 32416
rect 18509 32379 18567 32385
rect 8386 32348 8392 32360
rect 8347 32320 8392 32348
rect 8386 32308 8392 32320
rect 8444 32308 8450 32360
rect 8496 32280 8524 32376
rect 12710 32348 12716 32360
rect 12671 32320 12716 32348
rect 12710 32308 12716 32320
rect 12768 32308 12774 32360
rect 15286 32348 15292 32360
rect 15247 32320 15292 32348
rect 15286 32308 15292 32320
rect 15344 32308 15350 32360
rect 15565 32351 15623 32357
rect 15565 32317 15577 32351
rect 15611 32348 15623 32351
rect 15746 32348 15752 32360
rect 15611 32320 15752 32348
rect 15611 32317 15623 32320
rect 15565 32311 15623 32317
rect 15746 32308 15752 32320
rect 15804 32308 15810 32360
rect 18524 32348 18552 32379
rect 19150 32376 19156 32388
rect 19208 32376 19214 32428
rect 19797 32419 19855 32425
rect 19797 32385 19809 32419
rect 19843 32416 19855 32419
rect 20346 32416 20352 32428
rect 19843 32388 20352 32416
rect 19843 32385 19855 32388
rect 19797 32379 19855 32385
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 20530 32416 20536 32428
rect 20491 32388 20536 32416
rect 20530 32376 20536 32388
rect 20588 32416 20594 32428
rect 21177 32419 21235 32425
rect 21177 32416 21189 32419
rect 20588 32388 21189 32416
rect 20588 32376 20594 32388
rect 21177 32385 21189 32388
rect 21223 32385 21235 32419
rect 21177 32379 21235 32385
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32385 22247 32419
rect 22189 32379 22247 32385
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32416 23075 32419
rect 23106 32416 23112 32428
rect 23063 32388 23112 32416
rect 23063 32385 23075 32388
rect 23017 32379 23075 32385
rect 20438 32348 20444 32360
rect 18524 32320 20444 32348
rect 20438 32308 20444 32320
rect 20496 32308 20502 32360
rect 6236 32252 8524 32280
rect 6236 32240 6242 32252
rect 20346 32240 20352 32292
rect 20404 32280 20410 32292
rect 22204 32280 22232 32379
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 23290 32416 23296 32428
rect 23251 32388 23296 32416
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 23492 32416 23520 32515
rect 25314 32512 25320 32524
rect 25372 32512 25378 32564
rect 24854 32444 24860 32496
rect 24912 32484 24918 32496
rect 29546 32484 29552 32496
rect 24912 32456 26004 32484
rect 24912 32444 24918 32456
rect 24673 32419 24731 32425
rect 24673 32416 24685 32419
rect 23492 32388 24685 32416
rect 24673 32385 24685 32388
rect 24719 32385 24731 32419
rect 25498 32416 25504 32428
rect 25459 32388 25504 32416
rect 24673 32379 24731 32385
rect 25498 32376 25504 32388
rect 25556 32376 25562 32428
rect 25976 32425 26004 32456
rect 28460 32456 29552 32484
rect 28460 32425 28488 32456
rect 29546 32444 29552 32456
rect 29604 32444 29610 32496
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 28445 32419 28503 32425
rect 28445 32385 28457 32419
rect 28491 32385 28503 32419
rect 28445 32379 28503 32385
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 32398 32416 32404 32428
rect 32355 32388 32404 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 32582 32376 32588 32428
rect 32640 32416 32646 32428
rect 33318 32425 33324 32428
rect 33045 32419 33103 32425
rect 33045 32416 33057 32419
rect 32640 32388 33057 32416
rect 32640 32376 32646 32388
rect 33045 32385 33057 32388
rect 33091 32385 33103 32419
rect 33045 32379 33103 32385
rect 33312 32379 33324 32425
rect 33376 32416 33382 32428
rect 33376 32388 33412 32416
rect 33318 32376 33324 32379
rect 33376 32376 33382 32388
rect 23201 32351 23259 32357
rect 23201 32317 23213 32351
rect 23247 32348 23259 32351
rect 28626 32348 28632 32360
rect 23247 32320 23980 32348
rect 28587 32320 28632 32348
rect 23247 32317 23259 32320
rect 23201 32311 23259 32317
rect 22554 32280 22560 32292
rect 20404 32252 22560 32280
rect 20404 32240 20410 32252
rect 22554 32240 22560 32252
rect 22612 32240 22618 32292
rect 23952 32224 23980 32320
rect 28626 32308 28632 32320
rect 28684 32308 28690 32360
rect 28994 32348 29000 32360
rect 28955 32320 29000 32348
rect 28994 32308 29000 32320
rect 29052 32308 29058 32360
rect 32030 32308 32036 32360
rect 32088 32348 32094 32360
rect 32125 32351 32183 32357
rect 32125 32348 32137 32351
rect 32088 32320 32137 32348
rect 32088 32308 32094 32320
rect 32125 32317 32137 32320
rect 32171 32317 32183 32351
rect 32125 32311 32183 32317
rect 24857 32283 24915 32289
rect 24857 32249 24869 32283
rect 24903 32280 24915 32283
rect 25590 32280 25596 32292
rect 24903 32252 25596 32280
rect 24903 32249 24915 32252
rect 24857 32243 24915 32249
rect 25590 32240 25596 32252
rect 25648 32240 25654 32292
rect 1578 32212 1584 32224
rect 1539 32184 1584 32212
rect 1578 32172 1584 32184
rect 1636 32172 1642 32224
rect 7190 32212 7196 32224
rect 7103 32184 7196 32212
rect 7190 32172 7196 32184
rect 7248 32212 7254 32224
rect 8202 32212 8208 32224
rect 7248 32184 8208 32212
rect 7248 32172 7254 32184
rect 8202 32172 8208 32184
rect 8260 32172 8266 32224
rect 18966 32212 18972 32224
rect 18927 32184 18972 32212
rect 18966 32172 18972 32184
rect 19024 32172 19030 32224
rect 19610 32212 19616 32224
rect 19571 32184 19616 32212
rect 19610 32172 19616 32184
rect 19668 32172 19674 32224
rect 22002 32172 22008 32224
rect 22060 32212 22066 32224
rect 23293 32215 23351 32221
rect 23293 32212 23305 32215
rect 22060 32184 23305 32212
rect 22060 32172 22066 32184
rect 23293 32181 23305 32184
rect 23339 32212 23351 32215
rect 23382 32212 23388 32224
rect 23339 32184 23388 32212
rect 23339 32181 23351 32184
rect 23293 32175 23351 32181
rect 23382 32172 23388 32184
rect 23440 32172 23446 32224
rect 23934 32212 23940 32224
rect 23895 32184 23940 32212
rect 23934 32172 23940 32184
rect 23992 32172 23998 32224
rect 32493 32215 32551 32221
rect 32493 32181 32505 32215
rect 32539 32212 32551 32215
rect 33042 32212 33048 32224
rect 32539 32184 33048 32212
rect 32539 32181 32551 32184
rect 32493 32175 32551 32181
rect 33042 32172 33048 32184
rect 33100 32172 33106 32224
rect 34422 32212 34428 32224
rect 34383 32184 34428 32212
rect 34422 32172 34428 32184
rect 34480 32172 34486 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 4982 32008 4988 32020
rect 4943 31980 4988 32008
rect 4982 31968 4988 31980
rect 5040 31968 5046 32020
rect 15746 32008 15752 32020
rect 15707 31980 15752 32008
rect 15746 31968 15752 31980
rect 15804 31968 15810 32020
rect 16209 32011 16267 32017
rect 16209 31977 16221 32011
rect 16255 32008 16267 32011
rect 16390 32008 16396 32020
rect 16255 31980 16396 32008
rect 16255 31977 16267 31980
rect 16209 31971 16267 31977
rect 16390 31968 16396 31980
rect 16448 32008 16454 32020
rect 19610 32008 19616 32020
rect 16448 31980 19616 32008
rect 16448 31968 16454 31980
rect 19610 31968 19616 31980
rect 19668 31968 19674 32020
rect 21910 31968 21916 32020
rect 21968 32008 21974 32020
rect 22097 32011 22155 32017
rect 22097 32008 22109 32011
rect 21968 31980 22109 32008
rect 21968 31968 21974 31980
rect 22097 31977 22109 31980
rect 22143 32008 22155 32011
rect 23290 32008 23296 32020
rect 22143 31980 23296 32008
rect 22143 31977 22155 31980
rect 22097 31971 22155 31977
rect 23290 31968 23296 31980
rect 23348 31968 23354 32020
rect 33229 32011 33287 32017
rect 33229 31977 33241 32011
rect 33275 32008 33287 32011
rect 33318 32008 33324 32020
rect 33275 31980 33324 32008
rect 33275 31977 33287 31980
rect 33229 31971 33287 31977
rect 33318 31968 33324 31980
rect 33376 31968 33382 32020
rect 8294 31940 8300 31952
rect 5184 31912 8300 31940
rect 5184 31813 5212 31912
rect 8294 31900 8300 31912
rect 8352 31900 8358 31952
rect 17770 31900 17776 31952
rect 17828 31940 17834 31952
rect 20530 31940 20536 31952
rect 17828 31912 20536 31940
rect 17828 31900 17834 31912
rect 20530 31900 20536 31912
rect 20588 31940 20594 31952
rect 20993 31943 21051 31949
rect 20993 31940 21005 31943
rect 20588 31912 21005 31940
rect 20588 31900 20594 31912
rect 20993 31909 21005 31912
rect 21039 31909 21051 31943
rect 31202 31940 31208 31952
rect 20993 31903 21051 31909
rect 30760 31912 31208 31940
rect 5626 31872 5632 31884
rect 5587 31844 5632 31872
rect 5626 31832 5632 31844
rect 5684 31832 5690 31884
rect 6086 31872 6092 31884
rect 6047 31844 6092 31872
rect 6086 31832 6092 31844
rect 6144 31872 6150 31884
rect 12434 31872 12440 31884
rect 6144 31844 12440 31872
rect 6144 31832 6150 31844
rect 12434 31832 12440 31844
rect 12492 31872 12498 31884
rect 12492 31844 12537 31872
rect 12492 31832 12498 31844
rect 13262 31832 13268 31884
rect 13320 31872 13326 31884
rect 13357 31875 13415 31881
rect 13357 31872 13369 31875
rect 13320 31844 13369 31872
rect 13320 31832 13326 31844
rect 13357 31841 13369 31844
rect 13403 31841 13415 31875
rect 16022 31872 16028 31884
rect 15983 31844 16028 31872
rect 13357 31835 13415 31841
rect 16022 31832 16028 31844
rect 16080 31832 16086 31884
rect 16298 31872 16304 31884
rect 16132 31844 16304 31872
rect 5169 31807 5227 31813
rect 5169 31773 5181 31807
rect 5215 31773 5227 31807
rect 5169 31767 5227 31773
rect 13538 31764 13544 31816
rect 13596 31804 13602 31816
rect 14277 31807 14335 31813
rect 13596 31776 13641 31804
rect 13596 31764 13602 31776
rect 14277 31773 14289 31807
rect 14323 31804 14335 31807
rect 14918 31804 14924 31816
rect 14323 31776 14924 31804
rect 14323 31773 14335 31776
rect 14277 31767 14335 31773
rect 14918 31764 14924 31776
rect 14976 31764 14982 31816
rect 15933 31807 15991 31813
rect 15933 31773 15945 31807
rect 15979 31804 15991 31807
rect 16132 31804 16160 31844
rect 16298 31832 16304 31844
rect 16356 31832 16362 31884
rect 19613 31875 19671 31881
rect 19613 31841 19625 31875
rect 19659 31872 19671 31875
rect 19978 31872 19984 31884
rect 19659 31844 19984 31872
rect 19659 31841 19671 31844
rect 19613 31835 19671 31841
rect 19978 31832 19984 31844
rect 20036 31832 20042 31884
rect 15979 31776 16160 31804
rect 16209 31807 16267 31813
rect 15979 31773 15991 31776
rect 15933 31767 15991 31773
rect 16209 31773 16221 31807
rect 16255 31804 16267 31807
rect 16482 31804 16488 31816
rect 16255 31776 16488 31804
rect 16255 31773 16267 31776
rect 16209 31767 16267 31773
rect 16482 31764 16488 31776
rect 16540 31764 16546 31816
rect 18966 31764 18972 31816
rect 19024 31804 19030 31816
rect 20548 31813 20576 31900
rect 21008 31872 21036 31903
rect 22646 31872 22652 31884
rect 21008 31844 22652 31872
rect 22646 31832 22652 31844
rect 22704 31832 22710 31884
rect 30760 31881 30788 31912
rect 31202 31900 31208 31912
rect 31260 31900 31266 31952
rect 30745 31875 30803 31881
rect 30745 31841 30757 31875
rect 30791 31841 30803 31875
rect 30926 31872 30932 31884
rect 30887 31844 30932 31872
rect 30745 31835 30803 31841
rect 30926 31832 30932 31844
rect 30984 31832 30990 31884
rect 31570 31872 31576 31884
rect 31531 31844 31576 31872
rect 31570 31832 31576 31844
rect 31628 31832 31634 31884
rect 19429 31807 19487 31813
rect 19429 31804 19441 31807
rect 19024 31776 19441 31804
rect 19024 31764 19030 31776
rect 19429 31773 19441 31776
rect 19475 31773 19487 31807
rect 19429 31767 19487 31773
rect 19705 31807 19763 31813
rect 19705 31773 19717 31807
rect 19751 31804 19763 31807
rect 20533 31807 20591 31813
rect 19751 31776 20392 31804
rect 19751 31773 19763 31776
rect 19705 31767 19763 31773
rect 5810 31736 5816 31748
rect 5771 31708 5816 31736
rect 5810 31696 5816 31708
rect 5868 31696 5874 31748
rect 18690 31628 18696 31680
rect 18748 31668 18754 31680
rect 20364 31677 20392 31776
rect 20533 31773 20545 31807
rect 20579 31773 20591 31807
rect 20533 31767 20591 31773
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31804 22339 31807
rect 22370 31804 22376 31816
rect 22327 31776 22376 31804
rect 22327 31773 22339 31776
rect 22281 31767 22339 31773
rect 22370 31764 22376 31776
rect 22428 31804 22434 31816
rect 22741 31807 22799 31813
rect 22741 31804 22753 31807
rect 22428 31776 22753 31804
rect 22428 31764 22434 31776
rect 22741 31773 22753 31776
rect 22787 31773 22799 31807
rect 23014 31804 23020 31816
rect 22975 31776 23020 31804
rect 22741 31767 22799 31773
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 33042 31804 33048 31816
rect 33003 31776 33048 31804
rect 33042 31764 33048 31776
rect 33100 31764 33106 31816
rect 19245 31671 19303 31677
rect 19245 31668 19257 31671
rect 18748 31640 19257 31668
rect 18748 31628 18754 31640
rect 19245 31637 19257 31640
rect 19291 31637 19303 31671
rect 19245 31631 19303 31637
rect 20349 31671 20407 31677
rect 20349 31637 20361 31671
rect 20395 31668 20407 31671
rect 22186 31668 22192 31680
rect 20395 31640 22192 31668
rect 20395 31637 20407 31640
rect 20349 31631 20407 31637
rect 22186 31628 22192 31640
rect 22244 31668 22250 31680
rect 23106 31668 23112 31680
rect 22244 31640 23112 31668
rect 22244 31628 22250 31640
rect 23106 31628 23112 31640
rect 23164 31628 23170 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 5534 31464 5540 31476
rect 5495 31436 5540 31464
rect 5534 31424 5540 31436
rect 5592 31424 5598 31476
rect 5810 31424 5816 31476
rect 5868 31464 5874 31476
rect 6365 31467 6423 31473
rect 6365 31464 6377 31467
rect 5868 31436 6377 31464
rect 5868 31424 5874 31436
rect 6365 31433 6377 31436
rect 6411 31433 6423 31467
rect 6365 31427 6423 31433
rect 19889 31467 19947 31473
rect 19889 31433 19901 31467
rect 19935 31464 19947 31467
rect 19978 31464 19984 31476
rect 19935 31436 19984 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 19978 31424 19984 31436
rect 20036 31424 20042 31476
rect 24305 31467 24363 31473
rect 24305 31433 24317 31467
rect 24351 31464 24363 31467
rect 25498 31464 25504 31476
rect 24351 31436 25504 31464
rect 24351 31433 24363 31436
rect 24305 31427 24363 31433
rect 25498 31424 25504 31436
rect 25556 31424 25562 31476
rect 32398 31424 32404 31476
rect 32456 31464 32462 31476
rect 32677 31467 32735 31473
rect 32677 31464 32689 31467
rect 32456 31436 32689 31464
rect 32456 31424 32462 31436
rect 32677 31433 32689 31436
rect 32723 31433 32735 31467
rect 32677 31427 32735 31433
rect 35069 31467 35127 31473
rect 35069 31433 35081 31467
rect 35115 31464 35127 31467
rect 35342 31464 35348 31476
rect 35115 31436 35348 31464
rect 35115 31433 35127 31436
rect 35069 31427 35127 31433
rect 35342 31424 35348 31436
rect 35400 31424 35406 31476
rect 1578 31356 1584 31408
rect 1636 31396 1642 31408
rect 2501 31399 2559 31405
rect 2501 31396 2513 31399
rect 1636 31368 2513 31396
rect 1636 31356 1642 31368
rect 2501 31365 2513 31368
rect 2547 31365 2559 31399
rect 7282 31396 7288 31408
rect 7243 31368 7288 31396
rect 2501 31359 2559 31365
rect 7282 31356 7288 31368
rect 7340 31356 7346 31408
rect 14737 31399 14795 31405
rect 14737 31365 14749 31399
rect 14783 31396 14795 31399
rect 15286 31396 15292 31408
rect 14783 31368 15292 31396
rect 14783 31365 14795 31368
rect 14737 31359 14795 31365
rect 15286 31356 15292 31368
rect 15344 31356 15350 31408
rect 21726 31356 21732 31408
rect 21784 31396 21790 31408
rect 21821 31399 21879 31405
rect 21821 31396 21833 31399
rect 21784 31368 21833 31396
rect 21784 31356 21790 31368
rect 21821 31365 21833 31368
rect 21867 31365 21879 31399
rect 21821 31359 21879 31365
rect 23290 31356 23296 31408
rect 23348 31396 23354 31408
rect 23348 31368 24164 31396
rect 23348 31356 23354 31368
rect 1394 31328 1400 31340
rect 1355 31300 1400 31328
rect 1394 31288 1400 31300
rect 1452 31288 1458 31340
rect 2777 31331 2835 31337
rect 2777 31297 2789 31331
rect 2823 31297 2835 31331
rect 2777 31291 2835 31297
rect 5721 31331 5779 31337
rect 5721 31297 5733 31331
rect 5767 31297 5779 31331
rect 5721 31291 5779 31297
rect 2498 31220 2504 31272
rect 2556 31260 2562 31272
rect 2593 31263 2651 31269
rect 2593 31260 2605 31263
rect 2556 31232 2605 31260
rect 2556 31220 2562 31232
rect 2593 31229 2605 31232
rect 2639 31229 2651 31263
rect 2593 31223 2651 31229
rect 1581 31195 1639 31201
rect 1581 31161 1593 31195
rect 1627 31192 1639 31195
rect 2792 31192 2820 31291
rect 5736 31260 5764 31291
rect 6362 31288 6368 31340
rect 6420 31328 6426 31340
rect 6549 31331 6607 31337
rect 6549 31328 6561 31331
rect 6420 31300 6561 31328
rect 6420 31288 6426 31300
rect 6549 31297 6561 31300
rect 6595 31297 6607 31331
rect 7466 31328 7472 31340
rect 7427 31300 7472 31328
rect 6549 31291 6607 31297
rect 7466 31288 7472 31300
rect 7524 31328 7530 31340
rect 8021 31331 8079 31337
rect 8021 31328 8033 31331
rect 7524 31300 8033 31328
rect 7524 31288 7530 31300
rect 8021 31297 8033 31300
rect 8067 31297 8079 31331
rect 8021 31291 8079 31297
rect 12345 31331 12403 31337
rect 12345 31297 12357 31331
rect 12391 31328 12403 31331
rect 13538 31328 13544 31340
rect 12391 31300 13544 31328
rect 12391 31297 12403 31300
rect 12345 31291 12403 31297
rect 13538 31288 13544 31300
rect 13596 31288 13602 31340
rect 14918 31288 14924 31340
rect 14976 31328 14982 31340
rect 14976 31300 15021 31328
rect 14976 31288 14982 31300
rect 21450 31288 21456 31340
rect 21508 31328 21514 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21508 31300 22017 31328
rect 21508 31288 21514 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22554 31328 22560 31340
rect 22515 31300 22560 31328
rect 22005 31291 22063 31297
rect 22554 31288 22560 31300
rect 22612 31288 22618 31340
rect 22830 31328 22836 31340
rect 22791 31300 22836 31328
rect 22830 31288 22836 31300
rect 22888 31288 22894 31340
rect 23106 31288 23112 31340
rect 23164 31328 23170 31340
rect 24136 31337 24164 31368
rect 31018 31356 31024 31408
rect 31076 31396 31082 31408
rect 31478 31396 31484 31408
rect 31076 31368 31484 31396
rect 31076 31356 31082 31368
rect 31478 31356 31484 31368
rect 31536 31396 31542 31408
rect 32309 31399 32367 31405
rect 32309 31396 32321 31399
rect 31536 31368 32321 31396
rect 31536 31356 31542 31368
rect 32309 31365 32321 31368
rect 32355 31365 32367 31399
rect 34422 31396 34428 31408
rect 32309 31359 32367 31365
rect 32416 31368 34428 31396
rect 32416 31340 32444 31368
rect 34422 31356 34428 31368
rect 34480 31396 34486 31408
rect 35161 31399 35219 31405
rect 35161 31396 35173 31399
rect 34480 31368 35173 31396
rect 34480 31356 34486 31368
rect 35161 31365 35173 31368
rect 35207 31365 35219 31399
rect 35161 31359 35219 31365
rect 23845 31331 23903 31337
rect 23845 31328 23857 31331
rect 23164 31300 23857 31328
rect 23164 31288 23170 31300
rect 23845 31297 23857 31300
rect 23891 31297 23903 31331
rect 23845 31291 23903 31297
rect 24121 31331 24179 31337
rect 24121 31297 24133 31331
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31328 27307 31331
rect 27338 31328 27344 31340
rect 27295 31300 27344 31328
rect 27295 31297 27307 31300
rect 27249 31291 27307 31297
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 30101 31331 30159 31337
rect 30101 31297 30113 31331
rect 30147 31328 30159 31331
rect 30926 31328 30932 31340
rect 30147 31300 30932 31328
rect 30147 31297 30159 31300
rect 30101 31291 30159 31297
rect 30926 31288 30932 31300
rect 30984 31288 30990 31340
rect 32122 31328 32128 31340
rect 32083 31300 32128 31328
rect 32122 31288 32128 31300
rect 32180 31288 32186 31340
rect 32398 31328 32404 31340
rect 32359 31300 32404 31328
rect 32398 31288 32404 31300
rect 32456 31288 32462 31340
rect 32490 31288 32496 31340
rect 32548 31328 32554 31340
rect 32548 31300 32593 31328
rect 32548 31288 32554 31300
rect 7098 31260 7104 31272
rect 5736 31232 7104 31260
rect 7098 31220 7104 31232
rect 7156 31220 7162 31272
rect 13078 31260 13084 31272
rect 13039 31232 13084 31260
rect 13078 31220 13084 31232
rect 13136 31220 13142 31272
rect 22848 31260 22876 31288
rect 23750 31260 23756 31272
rect 22848 31232 23756 31260
rect 23750 31220 23756 31232
rect 23808 31220 23814 31272
rect 23934 31220 23940 31272
rect 23992 31260 23998 31272
rect 24029 31263 24087 31269
rect 24029 31260 24041 31263
rect 23992 31232 24041 31260
rect 23992 31220 23998 31232
rect 24029 31229 24041 31232
rect 24075 31260 24087 31263
rect 24075 31232 24624 31260
rect 24075 31229 24087 31232
rect 24029 31223 24087 31229
rect 1627 31164 2820 31192
rect 1627 31161 1639 31164
rect 1581 31155 1639 31161
rect 24596 31136 24624 31232
rect 26234 31220 26240 31272
rect 26292 31260 26298 31272
rect 26973 31263 27031 31269
rect 26973 31260 26985 31263
rect 26292 31232 26985 31260
rect 26292 31220 26298 31232
rect 26973 31229 26985 31232
rect 27019 31229 27031 31263
rect 26973 31223 27031 31229
rect 27614 31220 27620 31272
rect 27672 31260 27678 31272
rect 29825 31263 29883 31269
rect 29825 31260 29837 31263
rect 27672 31232 29837 31260
rect 27672 31220 27678 31232
rect 29825 31229 29837 31232
rect 29871 31229 29883 31263
rect 29825 31223 29883 31229
rect 34885 31263 34943 31269
rect 34885 31229 34897 31263
rect 34931 31229 34943 31263
rect 34885 31223 34943 31229
rect 31386 31152 31392 31204
rect 31444 31192 31450 31204
rect 34241 31195 34299 31201
rect 34241 31192 34253 31195
rect 31444 31164 34253 31192
rect 31444 31152 31450 31164
rect 34241 31161 34253 31164
rect 34287 31192 34299 31195
rect 34900 31192 34928 31223
rect 34287 31164 34928 31192
rect 34287 31161 34299 31164
rect 34241 31155 34299 31161
rect 2498 31124 2504 31136
rect 2459 31096 2504 31124
rect 2498 31084 2504 31096
rect 2556 31084 2562 31136
rect 2866 31084 2872 31136
rect 2924 31124 2930 31136
rect 2961 31127 3019 31133
rect 2961 31124 2973 31127
rect 2924 31096 2973 31124
rect 2924 31084 2930 31096
rect 2961 31093 2973 31096
rect 3007 31093 3019 31127
rect 8938 31124 8944 31136
rect 8899 31096 8944 31124
rect 2961 31087 3019 31093
rect 8938 31084 8944 31096
rect 8996 31084 9002 31136
rect 21269 31127 21327 31133
rect 21269 31093 21281 31127
rect 21315 31124 21327 31127
rect 21450 31124 21456 31136
rect 21315 31096 21456 31124
rect 21315 31093 21327 31096
rect 21269 31087 21327 31093
rect 21450 31084 21456 31096
rect 21508 31084 21514 31136
rect 23382 31084 23388 31136
rect 23440 31124 23446 31136
rect 23845 31127 23903 31133
rect 23845 31124 23857 31127
rect 23440 31096 23857 31124
rect 23440 31084 23446 31096
rect 23845 31093 23857 31096
rect 23891 31093 23903 31127
rect 23845 31087 23903 31093
rect 24578 31084 24584 31136
rect 24636 31124 24642 31136
rect 24765 31127 24823 31133
rect 24765 31124 24777 31127
rect 24636 31096 24777 31124
rect 24636 31084 24642 31096
rect 24765 31093 24777 31096
rect 24811 31093 24823 31127
rect 31478 31124 31484 31136
rect 31439 31096 31484 31124
rect 24765 31087 24823 31093
rect 31478 31084 31484 31096
rect 31536 31084 31542 31136
rect 35434 31084 35440 31136
rect 35492 31124 35498 31136
rect 35529 31127 35587 31133
rect 35529 31124 35541 31127
rect 35492 31096 35541 31124
rect 35492 31084 35498 31096
rect 35529 31093 35541 31096
rect 35575 31093 35587 31127
rect 35529 31087 35587 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 6181 30923 6239 30929
rect 6181 30889 6193 30923
rect 6227 30889 6239 30923
rect 6362 30920 6368 30932
rect 6323 30892 6368 30920
rect 6181 30883 6239 30889
rect 1394 30852 1400 30864
rect 1355 30824 1400 30852
rect 1394 30812 1400 30824
rect 1452 30812 1458 30864
rect 6196 30852 6224 30883
rect 6362 30880 6368 30892
rect 6420 30880 6426 30932
rect 19978 30880 19984 30932
rect 20036 30920 20042 30932
rect 20806 30920 20812 30932
rect 20036 30892 20812 30920
rect 20036 30880 20042 30892
rect 20806 30880 20812 30892
rect 20864 30920 20870 30932
rect 21085 30923 21143 30929
rect 21085 30920 21097 30923
rect 20864 30892 21097 30920
rect 20864 30880 20870 30892
rect 21085 30889 21097 30892
rect 21131 30889 21143 30923
rect 21085 30883 21143 30889
rect 21913 30923 21971 30929
rect 21913 30889 21925 30923
rect 21959 30920 21971 30923
rect 22002 30920 22008 30932
rect 21959 30892 22008 30920
rect 21959 30889 21971 30892
rect 21913 30883 21971 30889
rect 7006 30852 7012 30864
rect 6196 30824 7012 30852
rect 7006 30812 7012 30824
rect 7064 30852 7070 30864
rect 7190 30852 7196 30864
rect 7064 30824 7196 30852
rect 7064 30812 7070 30824
rect 7190 30812 7196 30824
rect 7248 30812 7254 30864
rect 5534 30744 5540 30796
rect 5592 30784 5598 30796
rect 6089 30787 6147 30793
rect 6089 30784 6101 30787
rect 5592 30756 6101 30784
rect 5592 30744 5598 30756
rect 6089 30753 6101 30756
rect 6135 30784 6147 30787
rect 6270 30784 6276 30796
rect 6135 30756 6276 30784
rect 6135 30753 6147 30756
rect 6089 30747 6147 30753
rect 6270 30744 6276 30756
rect 6328 30744 6334 30796
rect 8938 30784 8944 30796
rect 8899 30756 8944 30784
rect 8938 30744 8944 30756
rect 8996 30744 9002 30796
rect 21100 30784 21128 30883
rect 22002 30880 22008 30892
rect 22060 30880 22066 30932
rect 25498 30880 25504 30932
rect 25556 30920 25562 30932
rect 25593 30923 25651 30929
rect 25593 30920 25605 30923
rect 25556 30892 25605 30920
rect 25556 30880 25562 30892
rect 25593 30889 25605 30892
rect 25639 30889 25651 30923
rect 25593 30883 25651 30889
rect 32033 30923 32091 30929
rect 32033 30889 32045 30923
rect 32079 30920 32091 30923
rect 32122 30920 32128 30932
rect 32079 30892 32128 30920
rect 32079 30889 32091 30892
rect 32033 30883 32091 30889
rect 22094 30812 22100 30864
rect 22152 30852 22158 30864
rect 22833 30855 22891 30861
rect 22152 30824 22197 30852
rect 22152 30812 22158 30824
rect 22833 30821 22845 30855
rect 22879 30852 22891 30855
rect 23934 30852 23940 30864
rect 22879 30824 23940 30852
rect 22879 30821 22891 30824
rect 22833 30815 22891 30821
rect 23934 30812 23940 30824
rect 23992 30812 23998 30864
rect 26053 30855 26111 30861
rect 26053 30821 26065 30855
rect 26099 30852 26111 30855
rect 32048 30852 32076 30883
rect 32122 30880 32128 30892
rect 32180 30880 32186 30932
rect 26099 30824 27384 30852
rect 26099 30821 26111 30824
rect 26053 30815 26111 30821
rect 21729 30787 21787 30793
rect 21729 30784 21741 30787
rect 21100 30756 21741 30784
rect 21729 30753 21741 30756
rect 21775 30753 21787 30787
rect 21729 30747 21787 30753
rect 25406 30744 25412 30796
rect 25464 30784 25470 30796
rect 27356 30793 27384 30824
rect 29564 30824 32076 30852
rect 25685 30787 25743 30793
rect 25685 30784 25697 30787
rect 25464 30756 25697 30784
rect 25464 30744 25470 30756
rect 25685 30753 25697 30756
rect 25731 30753 25743 30787
rect 25685 30747 25743 30753
rect 27341 30787 27399 30793
rect 27341 30753 27353 30787
rect 27387 30753 27399 30787
rect 27341 30747 27399 30753
rect 27617 30787 27675 30793
rect 27617 30753 27629 30787
rect 27663 30784 27675 30787
rect 28626 30784 28632 30796
rect 27663 30756 28632 30784
rect 27663 30753 27675 30756
rect 27617 30747 27675 30753
rect 28626 30744 28632 30756
rect 28684 30744 28690 30796
rect 2774 30716 2780 30728
rect 2735 30688 2780 30716
rect 2774 30676 2780 30688
rect 2832 30676 2838 30728
rect 6178 30716 6184 30728
rect 6139 30688 6184 30716
rect 6178 30676 6184 30688
rect 6236 30676 6242 30728
rect 12897 30719 12955 30725
rect 12897 30685 12909 30719
rect 12943 30716 12955 30719
rect 14458 30716 14464 30728
rect 12943 30688 14464 30716
rect 12943 30685 12955 30688
rect 12897 30679 12955 30685
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 17586 30676 17592 30728
rect 17644 30716 17650 30728
rect 17681 30719 17739 30725
rect 17681 30716 17693 30719
rect 17644 30688 17693 30716
rect 17644 30676 17650 30688
rect 17681 30685 17693 30688
rect 17727 30685 17739 30719
rect 18690 30716 18696 30728
rect 18651 30688 18696 30716
rect 17681 30679 17739 30685
rect 18690 30676 18696 30688
rect 18748 30676 18754 30728
rect 21910 30716 21916 30728
rect 21871 30688 21916 30716
rect 21910 30676 21916 30688
rect 21968 30676 21974 30728
rect 22186 30716 22192 30728
rect 22020 30688 22192 30716
rect 5074 30608 5080 30660
rect 5132 30648 5138 30660
rect 5905 30651 5963 30657
rect 5905 30648 5917 30651
rect 5132 30620 5917 30648
rect 5132 30608 5138 30620
rect 5905 30617 5917 30620
rect 5951 30617 5963 30651
rect 9122 30648 9128 30660
rect 9083 30620 9128 30648
rect 5905 30611 5963 30617
rect 9122 30608 9128 30620
rect 9180 30608 9186 30660
rect 10781 30651 10839 30657
rect 10781 30617 10793 30651
rect 10827 30648 10839 30651
rect 13078 30648 13084 30660
rect 10827 30620 13084 30648
rect 10827 30617 10839 30620
rect 10781 30611 10839 30617
rect 3234 30540 3240 30592
rect 3292 30580 3298 30592
rect 10796 30580 10824 30611
rect 13078 30608 13084 30620
rect 13136 30608 13142 30660
rect 21637 30651 21695 30657
rect 21637 30617 21649 30651
rect 21683 30648 21695 30651
rect 22020 30648 22048 30688
rect 22186 30676 22192 30688
rect 22244 30676 22250 30728
rect 25774 30676 25780 30728
rect 25832 30716 25838 30728
rect 25869 30719 25927 30725
rect 25869 30716 25881 30719
rect 25832 30688 25881 30716
rect 25832 30676 25838 30688
rect 25869 30685 25881 30688
rect 25915 30685 25927 30719
rect 25869 30679 25927 30685
rect 21683 30620 22048 30648
rect 22649 30651 22707 30657
rect 21683 30617 21695 30620
rect 21637 30611 21695 30617
rect 22649 30617 22661 30651
rect 22695 30648 22707 30651
rect 23293 30651 23351 30657
rect 23293 30648 23305 30651
rect 22695 30620 23305 30648
rect 22695 30617 22707 30620
rect 22649 30611 22707 30617
rect 23293 30617 23305 30620
rect 23339 30617 23351 30651
rect 25590 30648 25596 30660
rect 25551 30620 25596 30648
rect 23293 30611 23351 30617
rect 18506 30580 18512 30592
rect 3292 30552 10824 30580
rect 18467 30552 18512 30580
rect 3292 30540 3298 30552
rect 18506 30540 18512 30552
rect 18564 30540 18570 30592
rect 21450 30540 21456 30592
rect 21508 30580 21514 30592
rect 22664 30580 22692 30611
rect 25590 30608 25596 30620
rect 25648 30608 25654 30660
rect 29362 30608 29368 30660
rect 29420 30648 29426 30660
rect 29564 30657 29592 30824
rect 31389 30787 31447 30793
rect 31389 30753 31401 30787
rect 31435 30784 31447 30787
rect 32398 30784 32404 30796
rect 31435 30756 32404 30784
rect 31435 30753 31447 30756
rect 31389 30747 31447 30753
rect 32398 30744 32404 30756
rect 32456 30744 32462 30796
rect 29549 30651 29607 30657
rect 29549 30648 29561 30651
rect 29420 30620 29561 30648
rect 29420 30608 29426 30620
rect 29549 30617 29561 30620
rect 29595 30617 29607 30651
rect 29549 30611 29607 30617
rect 29638 30608 29644 30660
rect 29696 30648 29702 30660
rect 31205 30651 31263 30657
rect 31205 30648 31217 30651
rect 29696 30620 31217 30648
rect 29696 30608 29702 30620
rect 31205 30617 31217 30620
rect 31251 30617 31263 30651
rect 31205 30611 31263 30617
rect 21508 30552 22692 30580
rect 21508 30540 21514 30552
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 5074 30376 5080 30388
rect 5035 30348 5080 30376
rect 5074 30336 5080 30348
rect 5132 30336 5138 30388
rect 17773 30311 17831 30317
rect 17773 30277 17785 30311
rect 17819 30308 17831 30311
rect 18506 30308 18512 30320
rect 17819 30280 18512 30308
rect 17819 30277 17831 30280
rect 17773 30271 17831 30277
rect 18506 30268 18512 30280
rect 18564 30268 18570 30320
rect 22094 30308 22100 30320
rect 22066 30268 22100 30308
rect 22152 30268 22158 30320
rect 25501 30311 25559 30317
rect 25501 30277 25513 30311
rect 25547 30308 25559 30311
rect 25590 30308 25596 30320
rect 25547 30280 25596 30308
rect 25547 30277 25559 30280
rect 25501 30271 25559 30277
rect 25590 30268 25596 30280
rect 25648 30308 25654 30320
rect 26973 30311 27031 30317
rect 26973 30308 26985 30311
rect 25648 30280 26985 30308
rect 25648 30268 25654 30280
rect 26973 30277 26985 30280
rect 27019 30277 27031 30311
rect 31386 30308 31392 30320
rect 31347 30280 31392 30308
rect 26973 30271 27031 30277
rect 31386 30268 31392 30280
rect 31444 30268 31450 30320
rect 34790 30308 34796 30320
rect 33796 30280 34796 30308
rect 2774 30240 2780 30252
rect 2735 30212 2780 30240
rect 2774 30200 2780 30212
rect 2832 30200 2838 30252
rect 5074 30200 5080 30252
rect 5132 30240 5138 30252
rect 5261 30243 5319 30249
rect 5261 30240 5273 30243
rect 5132 30212 5273 30240
rect 5132 30200 5138 30212
rect 5261 30209 5273 30212
rect 5307 30240 5319 30243
rect 5721 30243 5779 30249
rect 5721 30240 5733 30243
rect 5307 30212 5733 30240
rect 5307 30209 5319 30212
rect 5261 30203 5319 30209
rect 5721 30209 5733 30212
rect 5767 30240 5779 30243
rect 7466 30240 7472 30252
rect 5767 30212 7472 30240
rect 5767 30209 5779 30212
rect 5721 30203 5779 30209
rect 7466 30200 7472 30212
rect 7524 30200 7530 30252
rect 14458 30200 14464 30252
rect 14516 30240 14522 30252
rect 17586 30240 17592 30252
rect 14516 30212 14561 30240
rect 17547 30212 17592 30240
rect 14516 30200 14522 30212
rect 17586 30200 17592 30212
rect 17644 30200 17650 30252
rect 21821 30243 21879 30249
rect 21821 30209 21833 30243
rect 21867 30240 21879 30243
rect 22066 30240 22094 30268
rect 25774 30240 25780 30252
rect 21867 30212 22094 30240
rect 25735 30212 25780 30240
rect 21867 30209 21879 30212
rect 21821 30203 21879 30209
rect 25774 30200 25780 30212
rect 25832 30240 25838 30252
rect 27249 30243 27307 30249
rect 27249 30240 27261 30243
rect 25832 30212 27261 30240
rect 25832 30200 25838 30212
rect 27249 30209 27261 30212
rect 27295 30209 27307 30243
rect 27249 30203 27307 30209
rect 28537 30243 28595 30249
rect 28537 30209 28549 30243
rect 28583 30240 28595 30243
rect 29638 30240 29644 30252
rect 28583 30212 29644 30240
rect 28583 30209 28595 30212
rect 28537 30203 28595 30209
rect 29638 30200 29644 30212
rect 29696 30200 29702 30252
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30240 29791 30243
rect 30282 30240 30288 30252
rect 29779 30212 30288 30240
rect 29779 30209 29791 30212
rect 29733 30203 29791 30209
rect 30282 30200 30288 30212
rect 30340 30240 30346 30252
rect 32582 30240 32588 30252
rect 30340 30212 32588 30240
rect 30340 30200 30346 30212
rect 32582 30200 32588 30212
rect 32640 30240 32646 30252
rect 33796 30249 33824 30280
rect 34790 30268 34796 30280
rect 34848 30268 34854 30320
rect 34054 30249 34060 30252
rect 33781 30243 33839 30249
rect 33781 30240 33793 30243
rect 32640 30212 33793 30240
rect 32640 30200 32646 30212
rect 33781 30209 33793 30212
rect 33827 30209 33839 30243
rect 33781 30203 33839 30209
rect 34048 30203 34060 30249
rect 34112 30240 34118 30252
rect 34112 30212 34148 30240
rect 34054 30200 34060 30203
rect 34112 30200 34118 30212
rect 2958 30172 2964 30184
rect 2919 30144 2964 30172
rect 2958 30132 2964 30144
rect 3016 30132 3022 30184
rect 3234 30172 3240 30184
rect 3195 30144 3240 30172
rect 3234 30132 3240 30144
rect 3292 30132 3298 30184
rect 7006 30172 7012 30184
rect 6967 30144 7012 30172
rect 7006 30132 7012 30144
rect 7064 30132 7070 30184
rect 7282 30172 7288 30184
rect 7243 30144 7288 30172
rect 7282 30132 7288 30144
rect 7340 30172 7346 30184
rect 7745 30175 7803 30181
rect 7745 30172 7757 30175
rect 7340 30144 7757 30172
rect 7340 30132 7346 30144
rect 7745 30141 7757 30144
rect 7791 30141 7803 30175
rect 7745 30135 7803 30141
rect 8481 30175 8539 30181
rect 8481 30141 8493 30175
rect 8527 30172 8539 30175
rect 8941 30175 8999 30181
rect 8941 30172 8953 30175
rect 8527 30144 8953 30172
rect 8527 30141 8539 30144
rect 8481 30135 8539 30141
rect 8941 30141 8953 30144
rect 8987 30141 8999 30175
rect 8941 30135 8999 30141
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30141 9183 30175
rect 9398 30172 9404 30184
rect 9359 30144 9404 30172
rect 9125 30135 9183 30141
rect 8386 30064 8392 30116
rect 8444 30104 8450 30116
rect 9140 30104 9168 30135
rect 9398 30132 9404 30144
rect 9456 30132 9462 30184
rect 13078 30172 13084 30184
rect 13039 30144 13084 30172
rect 13078 30132 13084 30144
rect 13136 30132 13142 30184
rect 14274 30172 14280 30184
rect 14235 30144 14280 30172
rect 14274 30132 14280 30144
rect 14332 30132 14338 30184
rect 18230 30172 18236 30184
rect 18191 30144 18236 30172
rect 18230 30132 18236 30144
rect 18288 30132 18294 30184
rect 22097 30175 22155 30181
rect 22097 30141 22109 30175
rect 22143 30172 22155 30175
rect 22278 30172 22284 30184
rect 22143 30144 22284 30172
rect 22143 30141 22155 30144
rect 22097 30135 22155 30141
rect 22278 30132 22284 30144
rect 22336 30132 22342 30184
rect 25406 30132 25412 30184
rect 25464 30172 25470 30184
rect 25593 30175 25651 30181
rect 25593 30172 25605 30175
rect 25464 30144 25605 30172
rect 25464 30132 25470 30144
rect 25593 30141 25605 30144
rect 25639 30172 25651 30175
rect 27065 30175 27123 30181
rect 27065 30172 27077 30175
rect 25639 30144 27077 30172
rect 25639 30141 25651 30144
rect 25593 30135 25651 30141
rect 27065 30141 27077 30144
rect 27111 30141 27123 30175
rect 28258 30172 28264 30184
rect 28219 30144 28264 30172
rect 27065 30135 27123 30141
rect 28258 30132 28264 30144
rect 28316 30132 28322 30184
rect 29270 30132 29276 30184
rect 29328 30172 29334 30184
rect 30009 30175 30067 30181
rect 30009 30172 30021 30175
rect 29328 30144 30021 30172
rect 29328 30132 29334 30144
rect 30009 30141 30021 30144
rect 30055 30141 30067 30175
rect 30009 30135 30067 30141
rect 8444 30076 9168 30104
rect 25961 30107 26019 30113
rect 8444 30064 8450 30076
rect 25961 30073 25973 30107
rect 26007 30104 26019 30107
rect 26234 30104 26240 30116
rect 26007 30076 26240 30104
rect 26007 30073 26019 30076
rect 25961 30067 26019 30073
rect 26234 30064 26240 30076
rect 26292 30064 26298 30116
rect 27433 30107 27491 30113
rect 27433 30073 27445 30107
rect 27479 30104 27491 30107
rect 27614 30104 27620 30116
rect 27479 30076 27620 30104
rect 27479 30073 27491 30076
rect 27433 30067 27491 30073
rect 27614 30064 27620 30076
rect 27672 30064 27678 30116
rect 2317 30039 2375 30045
rect 2317 30005 2329 30039
rect 2363 30036 2375 30039
rect 3786 30036 3792 30048
rect 2363 30008 3792 30036
rect 2363 30005 2375 30008
rect 2317 29999 2375 30005
rect 3786 29996 3792 30008
rect 3844 29996 3850 30048
rect 16666 30036 16672 30048
rect 16627 30008 16672 30036
rect 16666 29996 16672 30008
rect 16724 29996 16730 30048
rect 20901 30039 20959 30045
rect 20901 30005 20913 30039
rect 20947 30036 20959 30039
rect 22462 30036 22468 30048
rect 20947 30008 22468 30036
rect 20947 30005 20959 30008
rect 20901 29999 20959 30005
rect 22462 29996 22468 30008
rect 22520 29996 22526 30048
rect 25041 30039 25099 30045
rect 25041 30005 25053 30039
rect 25087 30036 25099 30039
rect 25222 30036 25228 30048
rect 25087 30008 25228 30036
rect 25087 30005 25099 30008
rect 25041 29999 25099 30005
rect 25222 29996 25228 30008
rect 25280 29996 25286 30048
rect 25498 30036 25504 30048
rect 25459 30008 25504 30036
rect 25498 29996 25504 30008
rect 25556 30036 25562 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 25556 30008 26985 30036
rect 25556 29996 25562 30008
rect 26973 30005 26985 30008
rect 27019 30005 27031 30039
rect 26973 29999 27031 30005
rect 35161 30039 35219 30045
rect 35161 30005 35173 30039
rect 35207 30036 35219 30039
rect 35342 30036 35348 30048
rect 35207 30008 35348 30036
rect 35207 30005 35219 30008
rect 35161 29999 35219 30005
rect 35342 29996 35348 30008
rect 35400 29996 35406 30048
rect 38102 30036 38108 30048
rect 38063 30008 38108 30036
rect 38102 29996 38108 30008
rect 38160 29996 38166 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1581 29835 1639 29841
rect 1581 29801 1593 29835
rect 1627 29832 1639 29835
rect 2498 29832 2504 29844
rect 1627 29804 2504 29832
rect 1627 29801 1639 29804
rect 1581 29795 1639 29801
rect 2498 29792 2504 29804
rect 2556 29792 2562 29844
rect 6178 29792 6184 29844
rect 6236 29832 6242 29844
rect 6825 29835 6883 29841
rect 6825 29832 6837 29835
rect 6236 29804 6837 29832
rect 6236 29792 6242 29804
rect 6825 29801 6837 29804
rect 6871 29801 6883 29835
rect 9122 29832 9128 29844
rect 9083 29804 9128 29832
rect 6825 29795 6883 29801
rect 9122 29792 9128 29804
rect 9180 29792 9186 29844
rect 14182 29792 14188 29844
rect 14240 29832 14246 29844
rect 14461 29835 14519 29841
rect 14461 29832 14473 29835
rect 14240 29804 14473 29832
rect 14240 29792 14246 29804
rect 14461 29801 14473 29804
rect 14507 29801 14519 29835
rect 14461 29795 14519 29801
rect 14921 29835 14979 29841
rect 14921 29801 14933 29835
rect 14967 29832 14979 29835
rect 15102 29832 15108 29844
rect 14967 29804 15108 29832
rect 14967 29801 14979 29804
rect 14921 29795 14979 29801
rect 15102 29792 15108 29804
rect 15160 29792 15166 29844
rect 3786 29696 3792 29708
rect 3747 29668 3792 29696
rect 3786 29656 3792 29668
rect 3844 29656 3850 29708
rect 4614 29696 4620 29708
rect 4575 29668 4620 29696
rect 4614 29656 4620 29668
rect 4672 29656 4678 29708
rect 13262 29696 13268 29708
rect 13223 29668 13268 29696
rect 13262 29656 13268 29668
rect 13320 29656 13326 29708
rect 14829 29699 14887 29705
rect 14829 29665 14841 29699
rect 14875 29696 14887 29699
rect 15010 29696 15016 29708
rect 14875 29668 15016 29696
rect 14875 29665 14887 29668
rect 14829 29659 14887 29665
rect 15010 29656 15016 29668
rect 15068 29656 15074 29708
rect 16666 29696 16672 29708
rect 16627 29668 16672 29696
rect 16666 29656 16672 29668
rect 16724 29656 16730 29708
rect 18509 29699 18567 29705
rect 18509 29665 18521 29699
rect 18555 29696 18567 29699
rect 19334 29696 19340 29708
rect 18555 29668 19340 29696
rect 18555 29665 18567 29668
rect 18509 29659 18567 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 20714 29696 20720 29708
rect 20675 29668 20720 29696
rect 20714 29656 20720 29668
rect 20772 29656 20778 29708
rect 22278 29696 22284 29708
rect 22239 29668 22284 29696
rect 22278 29656 22284 29668
rect 22336 29656 22342 29708
rect 22462 29696 22468 29708
rect 22423 29668 22468 29696
rect 22462 29656 22468 29668
rect 22520 29656 22526 29708
rect 25222 29696 25228 29708
rect 25183 29668 25228 29696
rect 25222 29656 25228 29668
rect 25280 29656 25286 29708
rect 26694 29696 26700 29708
rect 26655 29668 26700 29696
rect 26694 29656 26700 29668
rect 26752 29656 26758 29708
rect 34790 29656 34796 29708
rect 34848 29696 34854 29708
rect 36357 29699 36415 29705
rect 36357 29696 36369 29699
rect 34848 29668 36369 29696
rect 34848 29656 34854 29668
rect 36357 29665 36369 29668
rect 36403 29665 36415 29699
rect 36357 29659 36415 29665
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29628 1458 29640
rect 2041 29631 2099 29637
rect 2041 29628 2053 29631
rect 1452 29600 2053 29628
rect 1452 29588 1458 29600
rect 2041 29597 2053 29600
rect 2087 29597 2099 29631
rect 2041 29591 2099 29597
rect 3053 29631 3111 29637
rect 3053 29597 3065 29631
rect 3099 29628 3111 29631
rect 3694 29628 3700 29640
rect 3099 29600 3700 29628
rect 3099 29597 3111 29600
rect 3053 29591 3111 29597
rect 3694 29588 3700 29600
rect 3752 29588 3758 29640
rect 6638 29628 6644 29640
rect 6551 29600 6644 29628
rect 6638 29588 6644 29600
rect 6696 29628 6702 29640
rect 7285 29631 7343 29637
rect 7285 29628 7297 29631
rect 6696 29600 7297 29628
rect 6696 29588 6702 29600
rect 7285 29597 7297 29600
rect 7331 29597 7343 29631
rect 7285 29591 7343 29597
rect 8478 29588 8484 29640
rect 8536 29628 8542 29640
rect 8941 29631 8999 29637
rect 8941 29628 8953 29631
rect 8536 29600 8953 29628
rect 8536 29588 8542 29600
rect 8941 29597 8953 29600
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 9585 29631 9643 29637
rect 9585 29597 9597 29631
rect 9631 29597 9643 29631
rect 12250 29628 12256 29640
rect 12211 29600 12256 29628
rect 9585 29591 9643 29597
rect 3973 29563 4031 29569
rect 3973 29529 3985 29563
rect 4019 29529 4031 29563
rect 3973 29523 4031 29529
rect 3237 29495 3295 29501
rect 3237 29461 3249 29495
rect 3283 29492 3295 29495
rect 3988 29492 4016 29523
rect 8846 29520 8852 29572
rect 8904 29560 8910 29572
rect 9600 29560 9628 29591
rect 12250 29588 12256 29600
rect 12308 29588 12314 29640
rect 13541 29631 13599 29637
rect 13541 29597 13553 29631
rect 13587 29628 13599 29631
rect 13722 29628 13728 29640
rect 13587 29600 13728 29628
rect 13587 29597 13599 29600
rect 13541 29591 13599 29597
rect 13722 29588 13728 29600
rect 13780 29588 13786 29640
rect 14642 29628 14648 29640
rect 14603 29600 14648 29628
rect 14642 29588 14648 29600
rect 14700 29588 14706 29640
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 20530 29628 20536 29640
rect 19475 29600 20536 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 20530 29588 20536 29600
rect 20588 29588 20594 29640
rect 22646 29588 22652 29640
rect 22704 29628 22710 29640
rect 23109 29631 23167 29637
rect 23109 29628 23121 29631
rect 22704 29600 23121 29628
rect 22704 29588 22710 29600
rect 23109 29597 23121 29600
rect 23155 29628 23167 29631
rect 23569 29631 23627 29637
rect 23569 29628 23581 29631
rect 23155 29600 23581 29628
rect 23155 29597 23167 29600
rect 23109 29591 23167 29597
rect 23569 29597 23581 29600
rect 23615 29597 23627 29631
rect 23569 29591 23627 29597
rect 24486 29588 24492 29640
rect 24544 29628 24550 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 24544 29600 24593 29628
rect 24544 29588 24550 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 14918 29560 14924 29572
rect 8904 29532 9628 29560
rect 14879 29532 14924 29560
rect 8904 29520 8910 29532
rect 14918 29520 14924 29532
rect 14976 29520 14982 29572
rect 16850 29560 16856 29572
rect 16811 29532 16856 29560
rect 16850 29520 16856 29532
rect 16908 29520 16914 29572
rect 25409 29563 25467 29569
rect 25409 29529 25421 29563
rect 25455 29529 25467 29563
rect 25409 29523 25467 29529
rect 3283 29464 4016 29492
rect 3283 29461 3295 29464
rect 3237 29455 3295 29461
rect 4614 29452 4620 29504
rect 4672 29492 4678 29504
rect 9398 29492 9404 29504
rect 4672 29464 9404 29492
rect 4672 29452 4678 29464
rect 9398 29452 9404 29464
rect 9456 29492 9462 29504
rect 12710 29492 12716 29504
rect 9456 29464 12716 29492
rect 9456 29452 9462 29464
rect 12710 29452 12716 29464
rect 12768 29452 12774 29504
rect 22830 29452 22836 29504
rect 22888 29492 22894 29504
rect 22925 29495 22983 29501
rect 22925 29492 22937 29495
rect 22888 29464 22937 29492
rect 22888 29452 22894 29464
rect 22925 29461 22937 29464
rect 22971 29461 22983 29495
rect 22925 29455 22983 29461
rect 24765 29495 24823 29501
rect 24765 29461 24777 29495
rect 24811 29492 24823 29495
rect 25424 29492 25452 29523
rect 36446 29520 36452 29572
rect 36504 29560 36510 29572
rect 36602 29563 36660 29569
rect 36602 29560 36614 29563
rect 36504 29532 36614 29560
rect 36504 29520 36510 29532
rect 36602 29529 36614 29532
rect 36648 29529 36660 29563
rect 36602 29523 36660 29529
rect 24811 29464 25452 29492
rect 35713 29495 35771 29501
rect 24811 29461 24823 29464
rect 24765 29455 24823 29461
rect 35713 29461 35725 29495
rect 35759 29492 35771 29495
rect 35802 29492 35808 29504
rect 35759 29464 35808 29492
rect 35759 29461 35771 29464
rect 35713 29455 35771 29461
rect 35802 29452 35808 29464
rect 35860 29452 35866 29504
rect 37366 29452 37372 29504
rect 37424 29492 37430 29504
rect 37737 29495 37795 29501
rect 37737 29492 37749 29495
rect 37424 29464 37749 29492
rect 37424 29452 37430 29464
rect 37737 29461 37749 29464
rect 37783 29461 37795 29495
rect 37737 29455 37795 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 2869 29291 2927 29297
rect 2869 29257 2881 29291
rect 2915 29288 2927 29291
rect 2958 29288 2964 29300
rect 2915 29260 2964 29288
rect 2915 29257 2927 29260
rect 2869 29251 2927 29257
rect 2958 29248 2964 29260
rect 3016 29248 3022 29300
rect 8386 29288 8392 29300
rect 8347 29260 8392 29288
rect 8386 29248 8392 29260
rect 8444 29248 8450 29300
rect 15378 29288 15384 29300
rect 15339 29260 15384 29288
rect 15378 29248 15384 29260
rect 15436 29248 15442 29300
rect 16850 29288 16856 29300
rect 16811 29260 16856 29288
rect 16850 29248 16856 29260
rect 16908 29248 16914 29300
rect 22925 29291 22983 29297
rect 22925 29257 22937 29291
rect 22971 29257 22983 29291
rect 22925 29251 22983 29257
rect 14918 29220 14924 29232
rect 14831 29192 14924 29220
rect 14918 29180 14924 29192
rect 14976 29220 14982 29232
rect 16574 29220 16580 29232
rect 14976 29192 16580 29220
rect 14976 29180 14982 29192
rect 16574 29180 16580 29192
rect 16632 29180 16638 29232
rect 22465 29223 22523 29229
rect 22465 29189 22477 29223
rect 22511 29220 22523 29223
rect 22830 29220 22836 29232
rect 22511 29192 22836 29220
rect 22511 29189 22523 29192
rect 22465 29183 22523 29189
rect 22830 29180 22836 29192
rect 22888 29180 22894 29232
rect 22940 29220 22968 29251
rect 23014 29248 23020 29300
rect 23072 29288 23078 29300
rect 23658 29288 23664 29300
rect 23072 29260 23664 29288
rect 23072 29248 23078 29260
rect 23658 29248 23664 29260
rect 23716 29288 23722 29300
rect 24302 29288 24308 29300
rect 23716 29260 24308 29288
rect 23716 29248 23722 29260
rect 24302 29248 24308 29260
rect 24360 29248 24366 29300
rect 24486 29288 24492 29300
rect 24447 29260 24492 29288
rect 24486 29248 24492 29260
rect 24544 29248 24550 29300
rect 29270 29288 29276 29300
rect 29231 29260 29276 29288
rect 29270 29248 29276 29260
rect 29328 29248 29334 29300
rect 35161 29291 35219 29297
rect 35161 29257 35173 29291
rect 35207 29288 35219 29291
rect 36446 29288 36452 29300
rect 35207 29260 36124 29288
rect 36407 29260 36452 29288
rect 35207 29257 35219 29260
rect 35161 29251 35219 29257
rect 28258 29220 28264 29232
rect 22940 29192 28264 29220
rect 28258 29180 28264 29192
rect 28316 29180 28322 29232
rect 35342 29220 35348 29232
rect 34992 29192 35348 29220
rect 2685 29155 2743 29161
rect 2685 29121 2697 29155
rect 2731 29152 2743 29155
rect 3234 29152 3240 29164
rect 2731 29124 3240 29152
rect 2731 29121 2743 29124
rect 2685 29115 2743 29121
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 8205 29155 8263 29161
rect 8205 29121 8217 29155
rect 8251 29152 8263 29155
rect 8386 29152 8392 29164
rect 8251 29124 8392 29152
rect 8251 29121 8263 29124
rect 8205 29115 8263 29121
rect 8386 29112 8392 29124
rect 8444 29112 8450 29164
rect 8846 29152 8852 29164
rect 8807 29124 8852 29152
rect 8846 29112 8852 29124
rect 8904 29112 8910 29164
rect 12250 29152 12256 29164
rect 12211 29124 12256 29152
rect 12250 29112 12256 29124
rect 12308 29112 12314 29164
rect 14642 29112 14648 29164
rect 14700 29152 14706 29164
rect 15194 29152 15200 29164
rect 14700 29124 15200 29152
rect 14700 29112 14706 29124
rect 15194 29112 15200 29124
rect 15252 29112 15258 29164
rect 16666 29152 16672 29164
rect 16627 29124 16672 29152
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 20530 29112 20536 29164
rect 20588 29152 20594 29164
rect 21821 29155 21879 29161
rect 20588 29124 20633 29152
rect 20588 29112 20594 29124
rect 21821 29121 21833 29155
rect 21867 29121 21879 29155
rect 22738 29152 22744 29164
rect 22699 29124 22744 29152
rect 21821 29115 21879 29121
rect 2225 29087 2283 29093
rect 2225 29053 2237 29087
rect 2271 29084 2283 29087
rect 3329 29087 3387 29093
rect 3329 29084 3341 29087
rect 2271 29056 3341 29084
rect 2271 29053 2283 29056
rect 2225 29047 2283 29053
rect 3329 29053 3341 29056
rect 3375 29053 3387 29087
rect 3510 29084 3516 29096
rect 3471 29056 3516 29084
rect 3329 29047 3387 29053
rect 3510 29044 3516 29056
rect 3568 29044 3574 29096
rect 3878 29084 3884 29096
rect 3839 29056 3884 29084
rect 3878 29044 3884 29056
rect 3936 29084 3942 29096
rect 9030 29084 9036 29096
rect 3936 29056 6914 29084
rect 8991 29056 9036 29084
rect 3936 29044 3942 29056
rect 6886 29016 6914 29056
rect 9030 29044 9036 29056
rect 9088 29044 9094 29096
rect 10689 29087 10747 29093
rect 10689 29053 10701 29087
rect 10735 29053 10747 29087
rect 12434 29084 12440 29096
rect 12395 29056 12440 29084
rect 10689 29047 10747 29053
rect 10704 29016 10732 29047
rect 12434 29044 12440 29056
rect 12492 29044 12498 29096
rect 12710 29084 12716 29096
rect 12671 29056 12716 29084
rect 12710 29044 12716 29056
rect 12768 29044 12774 29096
rect 15010 29084 15016 29096
rect 14971 29056 15016 29084
rect 15010 29044 15016 29056
rect 15068 29044 15074 29096
rect 19153 29087 19211 29093
rect 19153 29053 19165 29087
rect 19199 29084 19211 29087
rect 19334 29084 19340 29096
rect 19199 29056 19340 29084
rect 19199 29053 19211 29056
rect 19153 29047 19211 29053
rect 19334 29044 19340 29056
rect 19392 29044 19398 29096
rect 20162 29044 20168 29096
rect 20220 29084 20226 29096
rect 20349 29087 20407 29093
rect 20349 29084 20361 29087
rect 20220 29056 20361 29084
rect 20220 29044 20226 29056
rect 20349 29053 20361 29056
rect 20395 29053 20407 29087
rect 20349 29047 20407 29053
rect 18230 29016 18236 29028
rect 6886 28988 18236 29016
rect 18230 28976 18236 28988
rect 18288 28976 18294 29028
rect 19978 28976 19984 29028
rect 20036 29016 20042 29028
rect 20438 29016 20444 29028
rect 20036 28988 20444 29016
rect 20036 28976 20042 28988
rect 20438 28976 20444 28988
rect 20496 29016 20502 29028
rect 21836 29016 21864 29115
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 22848 29152 22876 29180
rect 24029 29155 24087 29161
rect 24029 29152 24041 29155
rect 22848 29124 24041 29152
rect 24029 29121 24041 29124
rect 24075 29152 24087 29155
rect 24075 29124 24256 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 22557 29087 22615 29093
rect 22557 29053 22569 29087
rect 22603 29084 22615 29087
rect 24121 29087 24179 29093
rect 24121 29084 24133 29087
rect 22603 29056 24133 29084
rect 22603 29053 22615 29056
rect 22557 29047 22615 29053
rect 24121 29053 24133 29056
rect 24167 29053 24179 29087
rect 24228 29084 24256 29124
rect 24302 29112 24308 29164
rect 24360 29152 24366 29164
rect 29086 29152 29092 29164
rect 24360 29124 24405 29152
rect 29047 29124 29092 29152
rect 24360 29112 24366 29124
rect 29086 29112 29092 29124
rect 29144 29112 29150 29164
rect 34992 29161 35020 29192
rect 35342 29180 35348 29192
rect 35400 29180 35406 29232
rect 34977 29155 35035 29161
rect 34977 29121 34989 29155
rect 35023 29121 35035 29155
rect 35802 29152 35808 29164
rect 35763 29124 35808 29152
rect 34977 29115 35035 29121
rect 35802 29112 35808 29124
rect 35860 29112 35866 29164
rect 35986 29152 35992 29164
rect 35947 29124 35992 29152
rect 35986 29112 35992 29124
rect 36044 29112 36050 29164
rect 36096 29161 36124 29260
rect 36446 29248 36452 29260
rect 36504 29248 36510 29300
rect 36081 29155 36139 29161
rect 36081 29121 36093 29155
rect 36127 29121 36139 29155
rect 36081 29115 36139 29121
rect 36173 29155 36231 29161
rect 36173 29121 36185 29155
rect 36219 29152 36231 29155
rect 37366 29152 37372 29164
rect 36219 29124 37372 29152
rect 36219 29121 36231 29124
rect 36173 29115 36231 29121
rect 25590 29084 25596 29096
rect 24228 29056 25596 29084
rect 24121 29047 24179 29053
rect 20496 28988 21864 29016
rect 22005 29019 22063 29025
rect 20496 28976 20502 28988
rect 22005 28985 22017 29019
rect 22051 29016 22063 29019
rect 22572 29016 22600 29047
rect 22051 28988 22600 29016
rect 24136 29016 24164 29047
rect 25590 29044 25596 29056
rect 25648 29044 25654 29096
rect 35345 29087 35403 29093
rect 35345 29053 35357 29087
rect 35391 29084 35403 29087
rect 35894 29084 35900 29096
rect 35391 29056 35900 29084
rect 35391 29053 35403 29056
rect 35345 29047 35403 29053
rect 35894 29044 35900 29056
rect 35952 29044 35958 29096
rect 36096 29084 36124 29115
rect 37366 29112 37372 29124
rect 37424 29112 37430 29164
rect 36998 29084 37004 29096
rect 36096 29056 37004 29084
rect 36998 29044 37004 29056
rect 37056 29044 37062 29096
rect 25406 29016 25412 29028
rect 24136 28988 25412 29016
rect 22051 28985 22063 28988
rect 22005 28979 22063 28985
rect 25406 28976 25412 28988
rect 25464 28976 25470 29028
rect 15102 28908 15108 28960
rect 15160 28948 15166 28960
rect 15197 28951 15255 28957
rect 15197 28948 15209 28951
rect 15160 28920 15209 28948
rect 15160 28908 15166 28920
rect 15197 28917 15209 28920
rect 15243 28948 15255 28951
rect 15470 28948 15476 28960
rect 15243 28920 15476 28948
rect 15243 28917 15255 28920
rect 15197 28911 15255 28917
rect 15470 28908 15476 28920
rect 15528 28908 15534 28960
rect 22094 28908 22100 28960
rect 22152 28948 22158 28960
rect 22465 28951 22523 28957
rect 22465 28948 22477 28951
rect 22152 28920 22477 28948
rect 22152 28908 22158 28920
rect 22465 28917 22477 28920
rect 22511 28917 22523 28951
rect 22465 28911 22523 28917
rect 23750 28908 23756 28960
rect 23808 28948 23814 28960
rect 24029 28951 24087 28957
rect 24029 28948 24041 28951
rect 23808 28920 24041 28948
rect 23808 28908 23814 28920
rect 24029 28917 24041 28920
rect 24075 28917 24087 28951
rect 24029 28911 24087 28917
rect 34698 28908 34704 28960
rect 34756 28948 34762 28960
rect 34793 28951 34851 28957
rect 34793 28948 34805 28951
rect 34756 28920 34805 28948
rect 34756 28908 34762 28920
rect 34793 28917 34805 28920
rect 34839 28917 34851 28951
rect 34793 28911 34851 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 3237 28747 3295 28753
rect 3237 28713 3249 28747
rect 3283 28744 3295 28747
rect 3510 28744 3516 28756
rect 3283 28716 3516 28744
rect 3283 28713 3295 28716
rect 3237 28707 3295 28713
rect 3510 28704 3516 28716
rect 3568 28704 3574 28756
rect 3694 28704 3700 28756
rect 3752 28744 3758 28756
rect 3789 28747 3847 28753
rect 3789 28744 3801 28747
rect 3752 28716 3801 28744
rect 3752 28704 3758 28716
rect 3789 28713 3801 28716
rect 3835 28713 3847 28747
rect 3789 28707 3847 28713
rect 4249 28747 4307 28753
rect 4249 28713 4261 28747
rect 4295 28744 4307 28747
rect 4706 28744 4712 28756
rect 4295 28716 4712 28744
rect 4295 28713 4307 28716
rect 4249 28707 4307 28713
rect 4706 28704 4712 28716
rect 4764 28704 4770 28756
rect 7926 28744 7932 28756
rect 7887 28716 7932 28744
rect 7926 28704 7932 28716
rect 7984 28704 7990 28756
rect 8386 28744 8392 28756
rect 8347 28716 8392 28744
rect 8386 28704 8392 28716
rect 8444 28704 8450 28756
rect 9030 28704 9036 28756
rect 9088 28744 9094 28756
rect 9125 28747 9183 28753
rect 9125 28744 9137 28747
rect 9088 28716 9137 28744
rect 9088 28704 9094 28716
rect 9125 28713 9137 28716
rect 9171 28713 9183 28747
rect 15470 28744 15476 28756
rect 15431 28716 15476 28744
rect 9125 28707 9183 28713
rect 15470 28704 15476 28716
rect 15528 28704 15534 28756
rect 28445 28747 28503 28753
rect 28445 28713 28457 28747
rect 28491 28744 28503 28747
rect 29086 28744 29092 28756
rect 28491 28716 29092 28744
rect 28491 28713 28503 28716
rect 28445 28707 28503 28713
rect 29086 28704 29092 28716
rect 29144 28704 29150 28756
rect 35986 28704 35992 28756
rect 36044 28744 36050 28756
rect 37185 28747 37243 28753
rect 37185 28744 37197 28747
rect 36044 28716 37197 28744
rect 36044 28704 36050 28716
rect 37185 28713 37197 28716
rect 37231 28713 37243 28747
rect 37185 28707 37243 28713
rect 15286 28636 15292 28688
rect 15344 28676 15350 28688
rect 15841 28679 15899 28685
rect 15841 28676 15853 28679
rect 15344 28648 15853 28676
rect 15344 28636 15350 28648
rect 15841 28645 15853 28648
rect 15887 28645 15899 28679
rect 15841 28639 15899 28645
rect 4062 28608 4068 28620
rect 3975 28580 4068 28608
rect 4062 28568 4068 28580
rect 4120 28608 4126 28620
rect 5534 28608 5540 28620
rect 4120 28580 5540 28608
rect 4120 28568 4126 28580
rect 5534 28568 5540 28580
rect 5592 28568 5598 28620
rect 8018 28608 8024 28620
rect 7979 28580 8024 28608
rect 8018 28568 8024 28580
rect 8076 28568 8082 28620
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 13265 28611 13323 28617
rect 13265 28608 13277 28611
rect 12492 28580 13277 28608
rect 12492 28568 12498 28580
rect 13265 28577 13277 28580
rect 13311 28577 13323 28611
rect 13265 28571 13323 28577
rect 14274 28568 14280 28620
rect 14332 28608 14338 28620
rect 14369 28611 14427 28617
rect 14369 28608 14381 28611
rect 14332 28580 14381 28608
rect 14332 28568 14338 28580
rect 14369 28577 14381 28580
rect 14415 28577 14427 28611
rect 14369 28571 14427 28577
rect 14458 28568 14464 28620
rect 14516 28608 14522 28620
rect 15473 28611 15531 28617
rect 15473 28608 15485 28611
rect 14516 28580 15485 28608
rect 14516 28568 14522 28580
rect 15473 28577 15485 28580
rect 15519 28577 15531 28611
rect 18230 28608 18236 28620
rect 18191 28580 18236 28608
rect 15473 28571 15531 28577
rect 18230 28568 18236 28580
rect 18288 28568 18294 28620
rect 20162 28608 20168 28620
rect 20123 28580 20168 28608
rect 20162 28568 20168 28580
rect 20220 28568 20226 28620
rect 34790 28568 34796 28620
rect 34848 28608 34854 28620
rect 35253 28611 35311 28617
rect 35253 28608 35265 28611
rect 34848 28580 35265 28608
rect 34848 28568 34854 28580
rect 35253 28577 35265 28580
rect 35299 28577 35311 28611
rect 35253 28571 35311 28577
rect 36998 28568 37004 28620
rect 37056 28608 37062 28620
rect 37093 28611 37151 28617
rect 37093 28608 37105 28611
rect 37056 28580 37105 28608
rect 37056 28568 37062 28580
rect 37093 28577 37105 28580
rect 37139 28577 37151 28611
rect 37093 28571 37151 28577
rect 1394 28540 1400 28552
rect 1355 28512 1400 28540
rect 1394 28500 1400 28512
rect 1452 28540 1458 28552
rect 2041 28543 2099 28549
rect 2041 28540 2053 28543
rect 1452 28512 2053 28540
rect 1452 28500 1458 28512
rect 2041 28509 2053 28512
rect 2087 28509 2099 28543
rect 2041 28503 2099 28509
rect 3053 28543 3111 28549
rect 3053 28509 3065 28543
rect 3099 28540 3111 28543
rect 3694 28540 3700 28552
rect 3099 28512 3700 28540
rect 3099 28509 3111 28512
rect 3053 28503 3111 28509
rect 3694 28500 3700 28512
rect 3752 28500 3758 28552
rect 3878 28500 3884 28552
rect 3936 28540 3942 28552
rect 3973 28543 4031 28549
rect 3973 28540 3985 28543
rect 3936 28512 3985 28540
rect 3936 28500 3942 28512
rect 3973 28509 3985 28512
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 4154 28500 4160 28552
rect 4212 28540 4218 28552
rect 4249 28543 4307 28549
rect 4249 28540 4261 28543
rect 4212 28512 4261 28540
rect 4212 28500 4218 28512
rect 4249 28509 4261 28512
rect 4295 28540 4307 28543
rect 4982 28540 4988 28552
rect 4295 28512 4988 28540
rect 4295 28509 4307 28512
rect 4249 28503 4307 28509
rect 4982 28500 4988 28512
rect 5040 28500 5046 28552
rect 5258 28500 5264 28552
rect 5316 28540 5322 28552
rect 7834 28540 7840 28552
rect 5316 28512 7840 28540
rect 5316 28500 5322 28512
rect 7834 28500 7840 28512
rect 7892 28540 7898 28552
rect 7929 28543 7987 28549
rect 7929 28540 7941 28543
rect 7892 28512 7941 28540
rect 7892 28500 7898 28512
rect 7929 28509 7941 28512
rect 7975 28509 7987 28543
rect 8202 28540 8208 28552
rect 8163 28512 8208 28540
rect 7929 28503 7987 28509
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 8938 28540 8944 28552
rect 8899 28512 8944 28540
rect 8938 28500 8944 28512
rect 8996 28500 9002 28552
rect 13538 28540 13544 28552
rect 13499 28512 13544 28540
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 14090 28540 14096 28552
rect 14051 28512 14096 28540
rect 14090 28500 14096 28512
rect 14148 28500 14154 28552
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 15657 28543 15715 28549
rect 15657 28540 15669 28543
rect 15160 28512 15669 28540
rect 15160 28500 15166 28512
rect 15657 28509 15669 28512
rect 15703 28509 15715 28543
rect 16850 28540 16856 28552
rect 16811 28512 16856 28540
rect 15657 28503 15715 28509
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 20070 28500 20076 28552
rect 20128 28540 20134 28552
rect 20441 28543 20499 28549
rect 20441 28540 20453 28543
rect 20128 28512 20453 28540
rect 20128 28500 20134 28512
rect 20441 28509 20453 28512
rect 20487 28509 20499 28543
rect 20441 28503 20499 28509
rect 36446 28500 36452 28552
rect 36504 28540 36510 28552
rect 37277 28543 37335 28549
rect 37277 28540 37289 28543
rect 36504 28512 37289 28540
rect 36504 28500 36510 28512
rect 37277 28509 37289 28512
rect 37323 28509 37335 28543
rect 37277 28503 37335 28509
rect 37366 28500 37372 28552
rect 37424 28540 37430 28552
rect 37424 28512 37469 28540
rect 37424 28500 37430 28512
rect 15378 28472 15384 28484
rect 15339 28444 15384 28472
rect 15378 28432 15384 28444
rect 15436 28432 15442 28484
rect 17034 28472 17040 28484
rect 16995 28444 17040 28472
rect 17034 28432 17040 28444
rect 17092 28432 17098 28484
rect 28074 28472 28080 28484
rect 28035 28444 28080 28472
rect 28074 28432 28080 28444
rect 28132 28432 28138 28484
rect 28261 28475 28319 28481
rect 28261 28441 28273 28475
rect 28307 28472 28319 28475
rect 35520 28475 35578 28481
rect 28307 28444 29040 28472
rect 28307 28441 28319 28444
rect 28261 28435 28319 28441
rect 1578 28404 1584 28416
rect 1539 28376 1584 28404
rect 1578 28364 1584 28376
rect 1636 28364 1642 28416
rect 29012 28413 29040 28444
rect 35520 28441 35532 28475
rect 35566 28472 35578 28475
rect 35618 28472 35624 28484
rect 35566 28444 35624 28472
rect 35566 28441 35578 28444
rect 35520 28435 35578 28441
rect 35618 28432 35624 28444
rect 35676 28432 35682 28484
rect 37384 28472 37412 28500
rect 35866 28444 37412 28472
rect 28997 28407 29055 28413
rect 28997 28373 29009 28407
rect 29043 28404 29055 28407
rect 29270 28404 29276 28416
rect 29043 28376 29276 28404
rect 29043 28373 29055 28376
rect 28997 28367 29055 28373
rect 29270 28364 29276 28376
rect 29328 28364 29334 28416
rect 32306 28364 32312 28416
rect 32364 28404 32370 28416
rect 35866 28404 35894 28444
rect 32364 28376 35894 28404
rect 32364 28364 32370 28376
rect 35986 28364 35992 28416
rect 36044 28404 36050 28416
rect 36633 28407 36691 28413
rect 36633 28404 36645 28407
rect 36044 28376 36645 28404
rect 36044 28364 36050 28376
rect 36633 28373 36645 28376
rect 36679 28373 36691 28407
rect 36633 28367 36691 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3694 28200 3700 28212
rect 3655 28172 3700 28200
rect 3694 28160 3700 28172
rect 3752 28160 3758 28212
rect 8389 28203 8447 28209
rect 8389 28169 8401 28203
rect 8435 28200 8447 28203
rect 8478 28200 8484 28212
rect 8435 28172 8484 28200
rect 8435 28169 8447 28172
rect 8389 28163 8447 28169
rect 8478 28160 8484 28172
rect 8536 28160 8542 28212
rect 13722 28200 13728 28212
rect 13683 28172 13728 28200
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 15289 28203 15347 28209
rect 15289 28169 15301 28203
rect 15335 28200 15347 28203
rect 16666 28200 16672 28212
rect 15335 28172 16672 28200
rect 15335 28169 15347 28172
rect 15289 28163 15347 28169
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 20625 28203 20683 28209
rect 20625 28169 20637 28203
rect 20671 28200 20683 28203
rect 20806 28200 20812 28212
rect 20671 28172 20812 28200
rect 20671 28169 20683 28172
rect 20625 28163 20683 28169
rect 20806 28160 20812 28172
rect 20864 28200 20870 28212
rect 21085 28203 21143 28209
rect 21085 28200 21097 28203
rect 20864 28172 21097 28200
rect 20864 28160 20870 28172
rect 21085 28169 21097 28172
rect 21131 28169 21143 28203
rect 34054 28200 34060 28212
rect 34015 28172 34060 28200
rect 21085 28163 21143 28169
rect 34054 28160 34060 28172
rect 34112 28160 34118 28212
rect 4154 28132 4160 28144
rect 4115 28104 4160 28132
rect 4154 28092 4160 28104
rect 4212 28092 4218 28144
rect 7834 28092 7840 28144
rect 7892 28132 7898 28144
rect 7929 28135 7987 28141
rect 7929 28132 7941 28135
rect 7892 28104 7941 28132
rect 7892 28092 7898 28104
rect 7929 28101 7941 28104
rect 7975 28101 7987 28135
rect 7929 28095 7987 28101
rect 8294 28092 8300 28144
rect 8352 28132 8358 28144
rect 9217 28135 9275 28141
rect 9217 28132 9229 28135
rect 8352 28104 9229 28132
rect 8352 28092 8358 28104
rect 9217 28101 9229 28104
rect 9263 28101 9275 28135
rect 9217 28095 9275 28101
rect 14185 28135 14243 28141
rect 14185 28101 14197 28135
rect 14231 28132 14243 28135
rect 14366 28132 14372 28144
rect 14231 28104 14372 28132
rect 14231 28101 14243 28104
rect 14185 28095 14243 28101
rect 14366 28092 14372 28104
rect 14424 28132 14430 28144
rect 14829 28135 14887 28141
rect 14829 28132 14841 28135
rect 14424 28104 14841 28132
rect 14424 28092 14430 28104
rect 14829 28101 14841 28104
rect 14875 28132 14887 28135
rect 15378 28132 15384 28144
rect 14875 28104 15384 28132
rect 14875 28101 14887 28104
rect 14829 28095 14887 28101
rect 15378 28092 15384 28104
rect 15436 28092 15442 28144
rect 30282 28132 30288 28144
rect 27632 28104 30288 28132
rect 3694 28024 3700 28076
rect 3752 28064 3758 28076
rect 3878 28064 3884 28076
rect 3752 28036 3884 28064
rect 3752 28024 3758 28036
rect 3878 28024 3884 28036
rect 3936 28024 3942 28076
rect 3973 28067 4031 28073
rect 3973 28033 3985 28067
rect 4019 28064 4031 28067
rect 4062 28064 4068 28076
rect 4019 28036 4068 28064
rect 4019 28033 4031 28036
rect 3973 28027 4031 28033
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 8202 28064 8208 28076
rect 8163 28036 8208 28064
rect 8202 28024 8208 28036
rect 8260 28024 8266 28076
rect 13909 28067 13967 28073
rect 13909 28033 13921 28067
rect 13955 28064 13967 28067
rect 15102 28064 15108 28076
rect 13955 28036 15108 28064
rect 13955 28033 13967 28036
rect 13909 28027 13967 28033
rect 15102 28024 15108 28036
rect 15160 28024 15166 28076
rect 16850 28024 16856 28076
rect 16908 28064 16914 28076
rect 27632 28073 27660 28104
rect 30282 28092 30288 28104
rect 30340 28092 30346 28144
rect 31573 28135 31631 28141
rect 31573 28101 31585 28135
rect 31619 28132 31631 28135
rect 34698 28132 34704 28144
rect 31619 28104 34704 28132
rect 31619 28101 31631 28104
rect 31573 28095 31631 28101
rect 34698 28092 34704 28104
rect 34756 28092 34762 28144
rect 16945 28067 17003 28073
rect 16945 28064 16957 28067
rect 16908 28036 16957 28064
rect 16908 28024 16914 28036
rect 16945 28033 16957 28036
rect 16991 28033 17003 28067
rect 16945 28027 17003 28033
rect 27617 28067 27675 28073
rect 27617 28033 27629 28067
rect 27663 28033 27675 28067
rect 27617 28027 27675 28033
rect 27884 28067 27942 28073
rect 27884 28033 27896 28067
rect 27930 28064 27942 28067
rect 28166 28064 28172 28076
rect 27930 28036 28172 28064
rect 27930 28033 27942 28036
rect 27884 28027 27942 28033
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 30466 28064 30472 28076
rect 30427 28036 30472 28064
rect 30466 28024 30472 28036
rect 30524 28024 30530 28076
rect 30926 28024 30932 28076
rect 30984 28064 30990 28076
rect 31021 28067 31079 28073
rect 31021 28064 31033 28067
rect 30984 28036 31033 28064
rect 30984 28024 30990 28036
rect 31021 28033 31033 28036
rect 31067 28033 31079 28067
rect 31021 28027 31079 28033
rect 31113 28067 31171 28073
rect 31113 28033 31125 28067
rect 31159 28033 31171 28067
rect 31113 28027 31171 28033
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28033 31355 28067
rect 31297 28027 31355 28033
rect 8018 27996 8024 28008
rect 7979 27968 8024 27996
rect 8018 27956 8024 27968
rect 8076 27956 8082 28008
rect 14093 27999 14151 28005
rect 14093 27965 14105 27999
rect 14139 27996 14151 27999
rect 14458 27996 14464 28008
rect 14139 27968 14464 27996
rect 14139 27965 14151 27968
rect 14093 27959 14151 27965
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 14608 27968 14933 27996
rect 14608 27956 14614 27968
rect 14921 27965 14933 27968
rect 14967 27996 14979 27999
rect 15010 27996 15016 28008
rect 14967 27968 15016 27996
rect 14967 27965 14979 27968
rect 14921 27959 14979 27965
rect 15010 27956 15016 27968
rect 15068 27956 15074 28008
rect 3786 27888 3792 27940
rect 3844 27928 3850 27940
rect 4798 27928 4804 27940
rect 3844 27900 4804 27928
rect 3844 27888 3850 27900
rect 4798 27888 4804 27900
rect 4856 27888 4862 27940
rect 9401 27931 9459 27937
rect 9401 27897 9413 27931
rect 9447 27928 9459 27931
rect 20254 27928 20260 27940
rect 9447 27900 20260 27928
rect 9447 27897 9459 27900
rect 9401 27891 9459 27897
rect 20254 27888 20260 27900
rect 20312 27888 20318 27940
rect 28626 27888 28632 27940
rect 28684 27928 28690 27940
rect 28997 27931 29055 27937
rect 28997 27928 29009 27931
rect 28684 27900 29009 27928
rect 28684 27888 28690 27900
rect 28997 27897 29009 27900
rect 29043 27928 29055 27931
rect 31128 27928 31156 28027
rect 31312 27996 31340 28027
rect 31386 28024 31392 28076
rect 31444 28064 31450 28076
rect 32122 28064 32128 28076
rect 31444 28036 31489 28064
rect 32083 28036 32128 28064
rect 31444 28024 31450 28036
rect 32122 28024 32128 28036
rect 32180 28024 32186 28076
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 34238 28064 34244 28076
rect 34199 28036 34244 28064
rect 34238 28024 34244 28036
rect 34296 28024 34302 28076
rect 34977 28067 35035 28073
rect 34977 28033 34989 28067
rect 35023 28064 35035 28067
rect 35342 28064 35348 28076
rect 35023 28036 35348 28064
rect 35023 28033 35035 28036
rect 34977 28027 35035 28033
rect 35342 28024 35348 28036
rect 35400 28024 35406 28076
rect 35526 28024 35532 28076
rect 35584 28064 35590 28076
rect 36446 28064 36452 28076
rect 35584 28036 36452 28064
rect 35584 28024 35590 28036
rect 36446 28024 36452 28036
rect 36504 28024 36510 28076
rect 32493 27999 32551 28005
rect 32493 27996 32505 27999
rect 31312 27968 32505 27996
rect 32493 27965 32505 27968
rect 32539 27965 32551 27999
rect 34514 27996 34520 28008
rect 34475 27968 34520 27996
rect 32493 27959 32551 27965
rect 34514 27956 34520 27968
rect 34572 27996 34578 28008
rect 35253 27999 35311 28005
rect 35253 27996 35265 27999
rect 34572 27968 35265 27996
rect 34572 27956 34578 27968
rect 35253 27965 35265 27968
rect 35299 27996 35311 27999
rect 36633 27999 36691 28005
rect 36633 27996 36645 27999
rect 35299 27968 36645 27996
rect 35299 27965 35311 27968
rect 35253 27959 35311 27965
rect 36633 27965 36645 27968
rect 36679 27965 36691 27999
rect 36633 27959 36691 27965
rect 29043 27900 31156 27928
rect 29043 27897 29055 27900
rect 28997 27891 29055 27897
rect 4157 27863 4215 27869
rect 4157 27829 4169 27863
rect 4203 27860 4215 27863
rect 4706 27860 4712 27872
rect 4203 27832 4712 27860
rect 4203 27829 4215 27832
rect 4157 27823 4215 27829
rect 4706 27820 4712 27832
rect 4764 27820 4770 27872
rect 7926 27860 7932 27872
rect 7887 27832 7932 27860
rect 7926 27820 7932 27832
rect 7984 27820 7990 27872
rect 14185 27863 14243 27869
rect 14185 27829 14197 27863
rect 14231 27860 14243 27863
rect 15105 27863 15163 27869
rect 15105 27860 15117 27863
rect 14231 27832 15117 27860
rect 14231 27829 14243 27832
rect 14185 27823 14243 27829
rect 15105 27829 15117 27832
rect 15151 27860 15163 27863
rect 15470 27860 15476 27872
rect 15151 27832 15476 27860
rect 15151 27829 15163 27832
rect 15105 27823 15163 27829
rect 15470 27820 15476 27832
rect 15528 27820 15534 27872
rect 21818 27860 21824 27872
rect 21779 27832 21824 27860
rect 21818 27820 21824 27832
rect 21876 27820 21882 27872
rect 34422 27860 34428 27872
rect 34383 27832 34428 27860
rect 34422 27820 34428 27832
rect 34480 27820 34486 27872
rect 36262 27860 36268 27872
rect 36223 27832 36268 27860
rect 36262 27820 36268 27832
rect 36320 27820 36326 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 4249 27659 4307 27665
rect 4249 27625 4261 27659
rect 4295 27656 4307 27659
rect 4706 27656 4712 27668
rect 4295 27628 4712 27656
rect 4295 27625 4307 27628
rect 4249 27619 4307 27625
rect 4706 27616 4712 27628
rect 4764 27616 4770 27668
rect 7469 27659 7527 27665
rect 7469 27625 7481 27659
rect 7515 27656 7527 27659
rect 7926 27656 7932 27668
rect 7515 27628 7932 27656
rect 7515 27625 7527 27628
rect 7469 27619 7527 27625
rect 7926 27616 7932 27628
rect 7984 27616 7990 27668
rect 8389 27659 8447 27665
rect 8389 27625 8401 27659
rect 8435 27656 8447 27659
rect 8938 27656 8944 27668
rect 8435 27628 8944 27656
rect 8435 27625 8447 27628
rect 8389 27619 8447 27625
rect 8938 27616 8944 27628
rect 8996 27616 9002 27668
rect 14090 27656 14096 27668
rect 14051 27628 14096 27656
rect 14090 27616 14096 27628
rect 14148 27616 14154 27668
rect 14182 27616 14188 27668
rect 14240 27656 14246 27668
rect 14277 27659 14335 27665
rect 14277 27656 14289 27659
rect 14240 27628 14289 27656
rect 14240 27616 14246 27628
rect 14277 27625 14289 27628
rect 14323 27625 14335 27659
rect 20070 27656 20076 27668
rect 20031 27628 20076 27656
rect 14277 27619 14335 27625
rect 20070 27616 20076 27628
rect 20128 27616 20134 27668
rect 20257 27659 20315 27665
rect 20257 27656 20269 27659
rect 20180 27628 20269 27656
rect 3234 27548 3240 27600
rect 3292 27588 3298 27600
rect 3789 27591 3847 27597
rect 3789 27588 3801 27591
rect 3292 27560 3801 27588
rect 3292 27548 3298 27560
rect 3789 27557 3801 27560
rect 3835 27557 3847 27591
rect 3789 27551 3847 27557
rect 3970 27548 3976 27600
rect 4028 27588 4034 27600
rect 4028 27560 4108 27588
rect 4028 27548 4034 27560
rect 4080 27529 4108 27560
rect 4065 27523 4123 27529
rect 4065 27489 4077 27523
rect 4111 27489 4123 27523
rect 8018 27520 8024 27532
rect 7979 27492 8024 27520
rect 4065 27483 4123 27489
rect 8018 27480 8024 27492
rect 8076 27480 8082 27532
rect 9585 27523 9643 27529
rect 9585 27489 9597 27523
rect 9631 27520 9643 27523
rect 16485 27523 16543 27529
rect 9631 27492 16344 27520
rect 9631 27489 9643 27492
rect 9585 27483 9643 27489
rect 3694 27412 3700 27464
rect 3752 27452 3758 27464
rect 3973 27455 4031 27461
rect 3973 27452 3985 27455
rect 3752 27424 3985 27452
rect 3752 27412 3758 27424
rect 3973 27421 3985 27424
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 4154 27412 4160 27464
rect 4212 27452 4218 27464
rect 4249 27455 4307 27461
rect 4249 27452 4261 27455
rect 4212 27424 4261 27452
rect 4212 27412 4218 27424
rect 4249 27421 4261 27424
rect 4295 27452 4307 27455
rect 4614 27452 4620 27464
rect 4295 27424 4620 27452
rect 4295 27421 4307 27424
rect 4249 27415 4307 27421
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27452 4951 27455
rect 4939 27424 5304 27452
rect 4939 27421 4951 27424
rect 4893 27415 4951 27421
rect 5276 27328 5304 27424
rect 7098 27412 7104 27464
rect 7156 27452 7162 27464
rect 7285 27455 7343 27461
rect 7285 27452 7297 27455
rect 7156 27424 7297 27452
rect 7156 27412 7162 27424
rect 7285 27421 7297 27424
rect 7331 27421 7343 27455
rect 7285 27415 7343 27421
rect 7300 27384 7328 27415
rect 7834 27412 7840 27464
rect 7892 27452 7898 27464
rect 7929 27455 7987 27461
rect 7929 27452 7941 27455
rect 7892 27424 7941 27452
rect 7892 27412 7898 27424
rect 7929 27421 7941 27424
rect 7975 27421 7987 27455
rect 8202 27452 8208 27464
rect 8163 27424 8208 27452
rect 7929 27415 7987 27421
rect 8202 27412 8208 27424
rect 8260 27412 8266 27464
rect 14274 27452 14280 27464
rect 14235 27424 14280 27452
rect 14274 27412 14280 27424
rect 14332 27412 14338 27464
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27452 14427 27455
rect 14458 27452 14464 27464
rect 14415 27424 14464 27452
rect 14415 27421 14427 27424
rect 14369 27415 14427 27421
rect 9401 27387 9459 27393
rect 9401 27384 9413 27387
rect 7300 27356 9413 27384
rect 9401 27353 9413 27356
rect 9447 27353 9459 27387
rect 9401 27347 9459 27353
rect 13998 27344 14004 27396
rect 14056 27384 14062 27396
rect 14384 27384 14412 27415
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 15344 27424 16221 27452
rect 15344 27412 15350 27424
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16316 27452 16344 27492
rect 16485 27489 16497 27523
rect 16531 27520 16543 27523
rect 17034 27520 17040 27532
rect 16531 27492 17040 27520
rect 16531 27489 16543 27492
rect 16485 27483 16543 27489
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 20180 27452 20208 27628
rect 20257 27625 20269 27628
rect 20303 27656 20315 27659
rect 20806 27656 20812 27668
rect 20303 27628 20812 27656
rect 20303 27625 20315 27628
rect 20257 27619 20315 27625
rect 20806 27616 20812 27628
rect 20864 27656 20870 27668
rect 21269 27659 21327 27665
rect 21269 27656 21281 27659
rect 20864 27628 21281 27656
rect 20864 27616 20870 27628
rect 21269 27625 21281 27628
rect 21315 27656 21327 27659
rect 22002 27656 22008 27668
rect 21315 27628 22008 27656
rect 21315 27625 21327 27628
rect 21269 27619 21327 27625
rect 22002 27616 22008 27628
rect 22060 27616 22066 27668
rect 28166 27656 28172 27668
rect 28127 27628 28172 27656
rect 28166 27616 28172 27628
rect 28224 27616 28230 27668
rect 31386 27616 31392 27668
rect 31444 27656 31450 27668
rect 31481 27659 31539 27665
rect 31481 27656 31493 27659
rect 31444 27628 31493 27656
rect 31444 27616 31450 27628
rect 31481 27625 31493 27628
rect 31527 27625 31539 27659
rect 31481 27619 31539 27625
rect 33873 27659 33931 27665
rect 33873 27625 33885 27659
rect 33919 27656 33931 27659
rect 34238 27656 34244 27668
rect 33919 27628 34244 27656
rect 33919 27625 33931 27628
rect 33873 27619 33931 27625
rect 34238 27616 34244 27628
rect 34296 27616 34302 27668
rect 35618 27656 35624 27668
rect 35579 27628 35624 27656
rect 35618 27616 35624 27628
rect 35676 27616 35682 27668
rect 21729 27591 21787 27597
rect 21729 27557 21741 27591
rect 21775 27588 21787 27591
rect 22094 27588 22100 27600
rect 21775 27560 22100 27588
rect 21775 27557 21787 27560
rect 21729 27551 21787 27557
rect 22094 27548 22100 27560
rect 22152 27548 22158 27600
rect 35253 27591 35311 27597
rect 35253 27557 35265 27591
rect 35299 27588 35311 27591
rect 36262 27588 36268 27600
rect 35299 27560 36268 27588
rect 35299 27557 35311 27560
rect 35253 27551 35311 27557
rect 36262 27548 36268 27560
rect 36320 27548 36326 27600
rect 20441 27523 20499 27529
rect 20441 27489 20453 27523
rect 20487 27520 20499 27523
rect 20990 27520 20996 27532
rect 20487 27492 20996 27520
rect 20487 27489 20499 27492
rect 20441 27483 20499 27489
rect 20990 27480 20996 27492
rect 21048 27520 21054 27532
rect 21361 27523 21419 27529
rect 21361 27520 21373 27523
rect 21048 27492 21373 27520
rect 21048 27480 21054 27492
rect 21361 27489 21373 27492
rect 21407 27489 21419 27523
rect 22738 27520 22744 27532
rect 21361 27483 21419 27489
rect 22066 27492 22744 27520
rect 16316 27424 20208 27452
rect 16209 27415 16267 27421
rect 20254 27412 20260 27464
rect 20312 27452 20318 27464
rect 20533 27455 20591 27461
rect 20312 27424 20357 27452
rect 20312 27412 20318 27424
rect 20533 27421 20545 27455
rect 20579 27452 20591 27455
rect 20898 27452 20904 27464
rect 20579 27424 20904 27452
rect 20579 27421 20591 27424
rect 20533 27415 20591 27421
rect 20898 27412 20904 27424
rect 20956 27452 20962 27464
rect 21082 27452 21088 27464
rect 20956 27424 21088 27452
rect 20956 27412 20962 27424
rect 21082 27412 21088 27424
rect 21140 27452 21146 27464
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 21140 27424 21281 27452
rect 21140 27412 21146 27424
rect 21269 27421 21281 27424
rect 21315 27421 21327 27455
rect 21269 27415 21327 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27452 21603 27455
rect 22066 27452 22094 27492
rect 22738 27480 22744 27492
rect 22796 27480 22802 27532
rect 26513 27523 26571 27529
rect 26513 27489 26525 27523
rect 26559 27520 26571 27523
rect 27062 27520 27068 27532
rect 26559 27492 27068 27520
rect 26559 27489 26571 27492
rect 26513 27483 26571 27489
rect 27062 27480 27068 27492
rect 27120 27520 27126 27532
rect 27525 27523 27583 27529
rect 27525 27520 27537 27523
rect 27120 27492 27537 27520
rect 27120 27480 27126 27492
rect 27525 27489 27537 27492
rect 27571 27489 27583 27523
rect 35526 27520 35532 27532
rect 27525 27483 27583 27489
rect 34164 27492 35532 27520
rect 22370 27452 22376 27464
rect 21591 27424 22094 27452
rect 22331 27424 22376 27452
rect 21591 27421 21603 27424
rect 21545 27415 21603 27421
rect 14056 27356 14412 27384
rect 14553 27387 14611 27393
rect 14056 27344 14062 27356
rect 14553 27353 14565 27387
rect 14599 27384 14611 27387
rect 15562 27384 15568 27396
rect 14599 27356 15568 27384
rect 14599 27353 14611 27356
rect 14553 27347 14611 27353
rect 4706 27316 4712 27328
rect 4667 27288 4712 27316
rect 4706 27276 4712 27288
rect 4764 27276 4770 27328
rect 5258 27276 5264 27328
rect 5316 27316 5322 27328
rect 5353 27319 5411 27325
rect 5353 27316 5365 27319
rect 5316 27288 5365 27316
rect 5316 27276 5322 27288
rect 5353 27285 5365 27288
rect 5399 27316 5411 27319
rect 7282 27316 7288 27328
rect 5399 27288 7288 27316
rect 5399 27285 5411 27288
rect 5353 27279 5411 27285
rect 7282 27276 7288 27288
rect 7340 27276 7346 27328
rect 14366 27276 14372 27328
rect 14424 27316 14430 27328
rect 14568 27316 14596 27347
rect 15562 27344 15568 27356
rect 15620 27344 15626 27396
rect 20272 27384 20300 27412
rect 20622 27384 20628 27396
rect 20272 27356 20628 27384
rect 20622 27344 20628 27356
rect 20680 27384 20686 27396
rect 21560 27384 21588 27415
rect 22370 27412 22376 27424
rect 22428 27412 22434 27464
rect 22830 27452 22836 27464
rect 22791 27424 22836 27452
rect 22830 27412 22836 27424
rect 22888 27412 22894 27464
rect 26050 27412 26056 27464
rect 26108 27452 26114 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 26108 27424 28365 27452
rect 26108 27412 26114 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 28353 27415 28411 27421
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27421 31447 27455
rect 31389 27415 31447 27421
rect 31573 27455 31631 27461
rect 31573 27421 31585 27455
rect 31619 27452 31631 27455
rect 32306 27452 32312 27464
rect 31619 27424 32312 27452
rect 31619 27421 31631 27424
rect 31573 27415 31631 27421
rect 20680 27356 21588 27384
rect 27433 27387 27491 27393
rect 20680 27344 20686 27356
rect 27433 27353 27445 27387
rect 27479 27384 27491 27387
rect 27614 27384 27620 27396
rect 27479 27356 27620 27384
rect 27479 27353 27491 27356
rect 27433 27347 27491 27353
rect 27614 27344 27620 27356
rect 27672 27384 27678 27396
rect 28626 27384 28632 27396
rect 27672 27356 28632 27384
rect 27672 27344 27678 27356
rect 28626 27344 28632 27356
rect 28684 27344 28690 27396
rect 31404 27384 31432 27415
rect 32306 27412 32312 27424
rect 32364 27412 32370 27464
rect 34164 27461 34192 27492
rect 35526 27480 35532 27492
rect 35584 27480 35590 27532
rect 34149 27455 34207 27461
rect 34149 27421 34161 27455
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 34330 27412 34336 27464
rect 34388 27452 34394 27464
rect 35161 27455 35219 27461
rect 35161 27452 35173 27455
rect 34388 27424 35173 27452
rect 34388 27412 34394 27424
rect 35161 27421 35173 27424
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 35437 27455 35495 27461
rect 35437 27421 35449 27455
rect 35483 27452 35495 27455
rect 35618 27452 35624 27464
rect 35483 27424 35624 27452
rect 35483 27421 35495 27424
rect 35437 27415 35495 27421
rect 32122 27384 32128 27396
rect 31404 27356 32128 27384
rect 32122 27344 32128 27356
rect 32180 27344 32186 27396
rect 33873 27387 33931 27393
rect 33873 27353 33885 27387
rect 33919 27353 33931 27387
rect 35176 27384 35204 27415
rect 35618 27412 35624 27424
rect 35676 27452 35682 27464
rect 35802 27452 35808 27464
rect 35676 27424 35808 27452
rect 35676 27412 35682 27424
rect 35802 27412 35808 27424
rect 35860 27452 35866 27464
rect 36081 27455 36139 27461
rect 36081 27452 36093 27455
rect 35860 27424 36093 27452
rect 35860 27412 35866 27424
rect 36081 27421 36093 27424
rect 36127 27421 36139 27455
rect 36081 27415 36139 27421
rect 36262 27384 36268 27396
rect 35176 27356 36268 27384
rect 33873 27347 33931 27353
rect 14424 27288 14596 27316
rect 14424 27276 14430 27288
rect 22002 27276 22008 27328
rect 22060 27316 22066 27328
rect 22189 27319 22247 27325
rect 22189 27316 22201 27319
rect 22060 27288 22201 27316
rect 22060 27276 22066 27288
rect 22189 27285 22201 27288
rect 22235 27285 22247 27319
rect 26970 27316 26976 27328
rect 26931 27288 26976 27316
rect 22189 27279 22247 27285
rect 26970 27276 26976 27288
rect 27028 27276 27034 27328
rect 27338 27316 27344 27328
rect 27299 27288 27344 27316
rect 27338 27276 27344 27288
rect 27396 27316 27402 27328
rect 28350 27316 28356 27328
rect 27396 27288 28356 27316
rect 27396 27276 27402 27288
rect 28350 27276 28356 27288
rect 28408 27316 28414 27328
rect 28813 27319 28871 27325
rect 28813 27316 28825 27319
rect 28408 27288 28825 27316
rect 28408 27276 28414 27288
rect 28813 27285 28825 27288
rect 28859 27285 28871 27319
rect 28813 27279 28871 27285
rect 29270 27276 29276 27328
rect 29328 27316 29334 27328
rect 29825 27319 29883 27325
rect 29825 27316 29837 27319
rect 29328 27288 29837 27316
rect 29328 27276 29334 27288
rect 29825 27285 29837 27288
rect 29871 27285 29883 27319
rect 33318 27316 33324 27328
rect 33279 27288 33324 27316
rect 29825 27279 29883 27285
rect 33318 27276 33324 27288
rect 33376 27316 33382 27328
rect 33888 27316 33916 27347
rect 36262 27344 36268 27356
rect 36320 27344 36326 27396
rect 33376 27288 33916 27316
rect 34057 27319 34115 27325
rect 33376 27276 33382 27288
rect 34057 27285 34069 27319
rect 34103 27316 34115 27319
rect 34514 27316 34520 27328
rect 34103 27288 34520 27316
rect 34103 27285 34115 27288
rect 34057 27279 34115 27285
rect 34514 27276 34520 27288
rect 34572 27276 34578 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 5169 27115 5227 27121
rect 5169 27081 5181 27115
rect 5215 27112 5227 27115
rect 5534 27112 5540 27124
rect 5215 27084 5540 27112
rect 5215 27081 5227 27084
rect 5169 27075 5227 27081
rect 1394 26976 1400 26988
rect 1355 26948 1400 26976
rect 1394 26936 1400 26948
rect 1452 26976 1458 26988
rect 2041 26979 2099 26985
rect 2041 26976 2053 26979
rect 1452 26948 2053 26976
rect 1452 26936 1458 26948
rect 2041 26945 2053 26948
rect 2087 26945 2099 26979
rect 2041 26939 2099 26945
rect 4617 26979 4675 26985
rect 4617 26945 4629 26979
rect 4663 26976 4675 26979
rect 5184 26976 5212 27075
rect 5534 27072 5540 27084
rect 5592 27112 5598 27124
rect 6638 27112 6644 27124
rect 5592 27084 6644 27112
rect 5592 27072 5598 27084
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 7377 27115 7435 27121
rect 7377 27081 7389 27115
rect 7423 27112 7435 27115
rect 8202 27112 8208 27124
rect 7423 27084 8208 27112
rect 7423 27081 7435 27084
rect 7377 27075 7435 27081
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 13538 27072 13544 27124
rect 13596 27112 13602 27124
rect 13725 27115 13783 27121
rect 13725 27112 13737 27115
rect 13596 27084 13737 27112
rect 13596 27072 13602 27084
rect 13725 27081 13737 27084
rect 13771 27081 13783 27115
rect 15013 27115 15071 27121
rect 13725 27075 13783 27081
rect 14108 27084 14964 27112
rect 7282 27044 7288 27056
rect 7195 27016 7288 27044
rect 7208 26985 7236 27016
rect 7282 27004 7288 27016
rect 7340 27044 7346 27056
rect 8294 27044 8300 27056
rect 7340 27016 8300 27044
rect 7340 27004 7346 27016
rect 8294 27004 8300 27016
rect 8352 27004 8358 27056
rect 8754 27004 8760 27056
rect 8812 27044 8818 27056
rect 9125 27047 9183 27053
rect 9125 27044 9137 27047
rect 8812 27016 9137 27044
rect 8812 27004 8818 27016
rect 9125 27013 9137 27016
rect 9171 27044 9183 27047
rect 14108 27044 14136 27084
rect 9171 27016 14136 27044
rect 14185 27047 14243 27053
rect 9171 27013 9183 27016
rect 9125 27007 9183 27013
rect 14185 27013 14197 27047
rect 14231 27044 14243 27047
rect 14366 27044 14372 27056
rect 14231 27016 14372 27044
rect 14231 27013 14243 27016
rect 14185 27007 14243 27013
rect 14366 27004 14372 27016
rect 14424 27004 14430 27056
rect 4663 26948 5212 26976
rect 7193 26979 7251 26985
rect 4663 26945 4675 26948
rect 4617 26939 4675 26945
rect 7193 26945 7205 26979
rect 7239 26945 7251 26979
rect 7193 26939 7251 26945
rect 7650 26936 7656 26988
rect 7708 26976 7714 26988
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 7708 26948 7849 26976
rect 7708 26936 7714 26948
rect 7837 26945 7849 26948
rect 7883 26976 7895 26979
rect 9309 26979 9367 26985
rect 9309 26976 9321 26979
rect 7883 26948 9321 26976
rect 7883 26945 7895 26948
rect 7837 26939 7895 26945
rect 9309 26945 9321 26948
rect 9355 26945 9367 26979
rect 10042 26976 10048 26988
rect 10003 26948 10048 26976
rect 9309 26939 9367 26945
rect 10042 26936 10048 26948
rect 10100 26936 10106 26988
rect 13909 26979 13967 26985
rect 13909 26945 13921 26979
rect 13955 26976 13967 26979
rect 13955 26948 14136 26976
rect 13955 26945 13967 26948
rect 13909 26939 13967 26945
rect 8113 26911 8171 26917
rect 8113 26908 8125 26911
rect 7852 26880 8125 26908
rect 7852 26852 7880 26880
rect 8113 26877 8125 26880
rect 8159 26877 8171 26911
rect 13998 26908 14004 26920
rect 13959 26880 14004 26908
rect 8113 26871 8171 26877
rect 13998 26868 14004 26880
rect 14056 26868 14062 26920
rect 14108 26908 14136 26948
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 14829 26979 14887 26985
rect 14829 26976 14841 26979
rect 14792 26948 14841 26976
rect 14792 26936 14798 26948
rect 14829 26945 14841 26948
rect 14875 26945 14887 26979
rect 14936 26976 14964 27084
rect 15013 27081 15025 27115
rect 15059 27112 15071 27115
rect 15102 27112 15108 27124
rect 15059 27084 15108 27112
rect 15059 27081 15071 27084
rect 15013 27075 15071 27081
rect 15102 27072 15108 27084
rect 15160 27072 15166 27124
rect 15470 27112 15476 27124
rect 15431 27084 15476 27112
rect 15470 27072 15476 27084
rect 15528 27072 15534 27124
rect 26050 27112 26056 27124
rect 26011 27084 26056 27112
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 29641 27115 29699 27121
rect 29641 27112 29653 27115
rect 26252 27084 29653 27112
rect 20622 27004 20628 27056
rect 20680 27044 20686 27056
rect 22002 27044 22008 27056
rect 20680 27016 21128 27044
rect 21963 27016 22008 27044
rect 20680 27004 20686 27016
rect 15654 26976 15660 26988
rect 14936 26948 15240 26976
rect 15615 26948 15660 26976
rect 14829 26939 14887 26945
rect 14274 26908 14280 26920
rect 14108 26880 14280 26908
rect 14274 26868 14280 26880
rect 14332 26908 14338 26920
rect 15010 26908 15016 26920
rect 14332 26880 15016 26908
rect 14332 26868 14338 26880
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 7834 26800 7840 26852
rect 7892 26800 7898 26852
rect 15102 26840 15108 26852
rect 14200 26812 15108 26840
rect 14200 26784 14228 26812
rect 15102 26800 15108 26812
rect 15160 26800 15166 26852
rect 15212 26840 15240 26948
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20272 26948 20821 26976
rect 20162 26840 20168 26852
rect 15212 26812 20168 26840
rect 20162 26800 20168 26812
rect 20220 26840 20226 26852
rect 20272 26849 20300 26948
rect 20809 26945 20821 26948
rect 20855 26945 20867 26979
rect 20990 26976 20996 26988
rect 20951 26948 20996 26976
rect 20809 26939 20867 26945
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 21100 26985 21128 27016
rect 22002 27004 22008 27016
rect 22060 27004 22066 27056
rect 26252 27053 26280 27084
rect 29641 27081 29653 27084
rect 29687 27112 29699 27115
rect 33318 27112 33324 27124
rect 29687 27084 33324 27112
rect 29687 27081 29699 27084
rect 29641 27075 29699 27081
rect 33318 27072 33324 27084
rect 33376 27072 33382 27124
rect 34149 27115 34207 27121
rect 34149 27081 34161 27115
rect 34195 27112 34207 27115
rect 34422 27112 34428 27124
rect 34195 27084 34428 27112
rect 34195 27081 34207 27084
rect 34149 27075 34207 27081
rect 34422 27072 34428 27084
rect 34480 27072 34486 27124
rect 25593 27047 25651 27053
rect 25593 27013 25605 27047
rect 25639 27044 25651 27047
rect 26237 27047 26295 27053
rect 26237 27044 26249 27047
rect 25639 27016 26249 27044
rect 25639 27013 25651 27016
rect 25593 27007 25651 27013
rect 26237 27013 26249 27016
rect 26283 27013 26295 27047
rect 26237 27007 26295 27013
rect 26421 27047 26479 27053
rect 26421 27013 26433 27047
rect 26467 27044 26479 27047
rect 26970 27044 26976 27056
rect 26467 27016 26976 27044
rect 26467 27013 26479 27016
rect 26421 27007 26479 27013
rect 26970 27004 26976 27016
rect 27028 27004 27034 27056
rect 30460 27047 30518 27053
rect 30460 27013 30472 27047
rect 30506 27044 30518 27047
rect 30558 27044 30564 27056
rect 30506 27016 30564 27044
rect 30506 27013 30518 27016
rect 30460 27007 30518 27013
rect 30558 27004 30564 27016
rect 30616 27004 30622 27056
rect 21085 26979 21143 26985
rect 21085 26945 21097 26979
rect 21131 26945 21143 26979
rect 21818 26976 21824 26988
rect 21779 26948 21824 26976
rect 21085 26939 21143 26945
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 23382 26936 23388 26988
rect 23440 26976 23446 26988
rect 23661 26979 23719 26985
rect 23661 26976 23673 26979
rect 23440 26948 23673 26976
rect 23440 26936 23446 26948
rect 23661 26945 23673 26948
rect 23707 26976 23719 26979
rect 26326 26976 26332 26988
rect 23707 26948 26332 26976
rect 23707 26945 23719 26948
rect 23661 26939 23719 26945
rect 26326 26936 26332 26948
rect 26384 26936 26390 26988
rect 29270 26936 29276 26988
rect 29328 26976 29334 26988
rect 29365 26979 29423 26985
rect 29365 26976 29377 26979
rect 29328 26948 29377 26976
rect 29328 26936 29334 26948
rect 29365 26945 29377 26948
rect 29411 26945 29423 26979
rect 29365 26939 29423 26945
rect 30193 26979 30251 26985
rect 30193 26945 30205 26979
rect 30239 26976 30251 26979
rect 30282 26976 30288 26988
rect 30239 26948 30288 26976
rect 30239 26945 30251 26948
rect 30193 26939 30251 26945
rect 30282 26936 30288 26948
rect 30340 26936 30346 26988
rect 33594 26936 33600 26988
rect 33652 26976 33658 26988
rect 34057 26979 34115 26985
rect 34057 26976 34069 26979
rect 33652 26948 34069 26976
rect 33652 26936 33658 26948
rect 34057 26945 34069 26948
rect 34103 26945 34115 26979
rect 34057 26939 34115 26945
rect 34241 26979 34299 26985
rect 34241 26945 34253 26979
rect 34287 26976 34299 26979
rect 34330 26976 34336 26988
rect 34287 26948 34336 26976
rect 34287 26945 34299 26948
rect 34241 26939 34299 26945
rect 34330 26936 34336 26948
rect 34388 26936 34394 26988
rect 34698 26976 34704 26988
rect 34659 26948 34704 26976
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 34793 26979 34851 26985
rect 34793 26945 34805 26979
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 34977 26979 35035 26985
rect 34977 26945 34989 26979
rect 35023 26976 35035 26979
rect 35713 26979 35771 26985
rect 35713 26976 35725 26979
rect 35023 26948 35725 26976
rect 35023 26945 35035 26948
rect 34977 26939 35035 26945
rect 35713 26945 35725 26948
rect 35759 26976 35771 26979
rect 35894 26976 35900 26988
rect 35759 26948 35900 26976
rect 35759 26945 35771 26948
rect 35713 26939 35771 26945
rect 26973 26911 27031 26917
rect 26973 26877 26985 26911
rect 27019 26877 27031 26911
rect 27154 26908 27160 26920
rect 27115 26880 27160 26908
rect 26973 26871 27031 26877
rect 20257 26843 20315 26849
rect 20257 26840 20269 26843
rect 20220 26812 20269 26840
rect 20220 26800 20226 26812
rect 20257 26809 20269 26812
rect 20303 26809 20315 26843
rect 26988 26840 27016 26871
rect 27154 26868 27160 26880
rect 27212 26868 27218 26920
rect 27338 26868 27344 26920
rect 27396 26908 27402 26920
rect 27433 26911 27491 26917
rect 27433 26908 27445 26911
rect 27396 26880 27445 26908
rect 27396 26868 27402 26880
rect 27433 26877 27445 26880
rect 27479 26877 27491 26911
rect 27433 26871 27491 26877
rect 34422 26868 34428 26920
rect 34480 26908 34486 26920
rect 34808 26908 34836 26939
rect 35894 26936 35900 26948
rect 35952 26936 35958 26988
rect 34480 26880 34836 26908
rect 35989 26911 36047 26917
rect 34480 26868 34486 26880
rect 35989 26877 36001 26911
rect 36035 26908 36047 26911
rect 36262 26908 36268 26920
rect 36035 26880 36268 26908
rect 36035 26877 36047 26880
rect 35989 26871 36047 26877
rect 36262 26868 36268 26880
rect 36320 26868 36326 26920
rect 27614 26840 27620 26852
rect 26988 26812 27620 26840
rect 20257 26803 20315 26809
rect 27614 26800 27620 26812
rect 27672 26800 27678 26852
rect 34977 26843 35035 26849
rect 34977 26809 34989 26843
rect 35023 26840 35035 26843
rect 35526 26840 35532 26852
rect 35023 26812 35532 26840
rect 35023 26809 35035 26812
rect 34977 26803 35035 26809
rect 35526 26800 35532 26812
rect 35584 26800 35590 26852
rect 1581 26775 1639 26781
rect 1581 26741 1593 26775
rect 1627 26772 1639 26775
rect 2774 26772 2780 26784
rect 1627 26744 2780 26772
rect 1627 26741 1639 26744
rect 1581 26735 1639 26741
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 3694 26732 3700 26784
rect 3752 26772 3758 26784
rect 4433 26775 4491 26781
rect 4433 26772 4445 26775
rect 3752 26744 4445 26772
rect 3752 26732 3758 26744
rect 4433 26741 4445 26744
rect 4479 26741 4491 26775
rect 4433 26735 4491 26741
rect 9861 26775 9919 26781
rect 9861 26741 9873 26775
rect 9907 26772 9919 26775
rect 10594 26772 10600 26784
rect 9907 26744 10600 26772
rect 9907 26741 9919 26744
rect 9861 26735 9919 26741
rect 10594 26732 10600 26744
rect 10652 26732 10658 26784
rect 10689 26775 10747 26781
rect 10689 26741 10701 26775
rect 10735 26772 10747 26775
rect 10778 26772 10784 26784
rect 10735 26744 10784 26772
rect 10735 26741 10747 26744
rect 10689 26735 10747 26741
rect 10778 26732 10784 26744
rect 10836 26732 10842 26784
rect 14182 26772 14188 26784
rect 14095 26744 14188 26772
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 20806 26772 20812 26784
rect 20767 26744 20812 26772
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 21269 26775 21327 26781
rect 21269 26741 21281 26775
rect 21315 26772 21327 26775
rect 21726 26772 21732 26784
rect 21315 26744 21732 26772
rect 21315 26741 21327 26744
rect 21269 26735 21327 26741
rect 21726 26732 21732 26744
rect 21784 26732 21790 26784
rect 30374 26732 30380 26784
rect 30432 26772 30438 26784
rect 30926 26772 30932 26784
rect 30432 26744 30932 26772
rect 30432 26732 30438 26744
rect 30926 26732 30932 26744
rect 30984 26772 30990 26784
rect 31573 26775 31631 26781
rect 31573 26772 31585 26775
rect 30984 26744 31585 26772
rect 30984 26732 30990 26744
rect 31573 26741 31585 26744
rect 31619 26741 31631 26775
rect 33594 26772 33600 26784
rect 33555 26744 33600 26772
rect 31573 26735 31631 26741
rect 33594 26732 33600 26744
rect 33652 26732 33658 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 7926 26568 7932 26580
rect 7887 26540 7932 26568
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 15102 26568 15108 26580
rect 10336 26540 14320 26568
rect 15063 26540 15108 26568
rect 3970 26432 3976 26444
rect 3931 26404 3976 26432
rect 3970 26392 3976 26404
rect 4028 26392 4034 26444
rect 4798 26432 4804 26444
rect 4759 26404 4804 26432
rect 4798 26392 4804 26404
rect 4856 26432 4862 26444
rect 10336 26441 10364 26540
rect 14182 26500 14188 26512
rect 14143 26472 14188 26500
rect 14182 26460 14188 26472
rect 14240 26460 14246 26512
rect 14292 26500 14320 26540
rect 15102 26528 15108 26540
rect 15160 26528 15166 26580
rect 15286 26568 15292 26580
rect 15247 26540 15292 26568
rect 15286 26528 15292 26540
rect 15344 26528 15350 26580
rect 20162 26568 20168 26580
rect 20123 26540 20168 26568
rect 20162 26528 20168 26540
rect 20220 26528 20226 26580
rect 20806 26568 20812 26580
rect 20767 26540 20812 26568
rect 20806 26528 20812 26540
rect 20864 26528 20870 26580
rect 21177 26571 21235 26577
rect 21177 26537 21189 26571
rect 21223 26568 21235 26571
rect 22370 26568 22376 26580
rect 21223 26540 22376 26568
rect 21223 26537 21235 26540
rect 21177 26531 21235 26537
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 30469 26571 30527 26577
rect 30469 26537 30481 26571
rect 30515 26568 30527 26571
rect 30558 26568 30564 26580
rect 30515 26540 30564 26568
rect 30515 26537 30527 26540
rect 30469 26531 30527 26537
rect 30558 26528 30564 26540
rect 30616 26528 30622 26580
rect 19426 26500 19432 26512
rect 14292 26472 19432 26500
rect 19426 26460 19432 26472
rect 19484 26460 19490 26512
rect 10321 26435 10379 26441
rect 10321 26432 10333 26435
rect 4856 26404 10333 26432
rect 4856 26392 4862 26404
rect 10321 26401 10333 26404
rect 10367 26401 10379 26435
rect 10594 26432 10600 26444
rect 10555 26404 10600 26432
rect 10321 26395 10379 26401
rect 10594 26392 10600 26404
rect 10652 26392 10658 26444
rect 10778 26432 10784 26444
rect 10739 26404 10784 26432
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 13998 26392 14004 26444
rect 14056 26432 14062 26444
rect 14918 26432 14924 26444
rect 14056 26404 14924 26432
rect 14056 26392 14062 26404
rect 14918 26392 14924 26404
rect 14976 26392 14982 26444
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26364 3295 26367
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 3283 26336 3801 26364
rect 3283 26333 3295 26336
rect 3237 26327 3295 26333
rect 3789 26333 3801 26336
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 5626 26324 5632 26376
rect 5684 26364 5690 26376
rect 6641 26367 6699 26373
rect 6641 26364 6653 26367
rect 5684 26336 6653 26364
rect 5684 26324 5690 26336
rect 6641 26333 6653 26336
rect 6687 26333 6699 26367
rect 6641 26327 6699 26333
rect 6914 26324 6920 26376
rect 6972 26364 6978 26376
rect 8018 26364 8024 26376
rect 6972 26336 7017 26364
rect 7979 26336 8024 26364
rect 6972 26324 6978 26336
rect 8018 26324 8024 26336
rect 8076 26324 8082 26376
rect 8113 26367 8171 26373
rect 8113 26333 8125 26367
rect 8159 26364 8171 26367
rect 8202 26364 8208 26376
rect 8159 26336 8208 26364
rect 8159 26333 8171 26336
rect 8113 26327 8171 26333
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 12066 26364 12072 26376
rect 12027 26336 12072 26364
rect 12066 26324 12072 26336
rect 12124 26324 12130 26376
rect 14369 26367 14427 26373
rect 14369 26333 14381 26367
rect 14415 26333 14427 26367
rect 14369 26327 14427 26333
rect 7837 26299 7895 26305
rect 7837 26265 7849 26299
rect 7883 26296 7895 26299
rect 7926 26296 7932 26308
rect 7883 26268 7932 26296
rect 7883 26265 7895 26268
rect 7837 26259 7895 26265
rect 7926 26256 7932 26268
rect 7984 26256 7990 26308
rect 14384 26296 14412 26327
rect 15010 26324 15016 26376
rect 15068 26364 15074 26376
rect 15105 26367 15163 26373
rect 15105 26364 15117 26367
rect 15068 26336 15117 26364
rect 15068 26324 15074 26336
rect 15105 26333 15117 26336
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 18012 26336 18061 26364
rect 18012 26324 18018 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 20180 26364 20208 26528
rect 20990 26500 20996 26512
rect 20916 26472 20996 26500
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 20916 26441 20944 26472
rect 20990 26460 20996 26472
rect 21048 26460 21054 26512
rect 29362 26500 29368 26512
rect 26988 26472 29368 26500
rect 26988 26444 27016 26472
rect 29362 26460 29368 26472
rect 29420 26460 29426 26512
rect 38010 26500 38016 26512
rect 37971 26472 38016 26500
rect 38010 26460 38016 26472
rect 38068 26460 38074 26512
rect 20901 26435 20959 26441
rect 20680 26404 20852 26432
rect 20680 26392 20686 26404
rect 20717 26367 20775 26373
rect 20717 26364 20729 26367
rect 20180 26336 20729 26364
rect 18049 26327 18107 26333
rect 20717 26333 20729 26336
rect 20763 26333 20775 26367
rect 20824 26364 20852 26404
rect 20901 26401 20913 26435
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 22005 26435 22063 26441
rect 22005 26401 22017 26435
rect 22051 26432 22063 26435
rect 22830 26432 22836 26444
rect 22051 26404 22836 26432
rect 22051 26401 22063 26404
rect 22005 26395 22063 26401
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 23842 26432 23848 26444
rect 23803 26404 23848 26432
rect 23842 26392 23848 26404
rect 23900 26392 23906 26444
rect 26970 26432 26976 26444
rect 26931 26404 26976 26432
rect 26970 26392 26976 26404
rect 27028 26392 27034 26444
rect 27985 26435 28043 26441
rect 27985 26401 27997 26435
rect 28031 26432 28043 26435
rect 30374 26432 30380 26444
rect 28031 26404 30380 26432
rect 28031 26401 28043 26404
rect 27985 26395 28043 26401
rect 30374 26392 30380 26404
rect 30432 26392 30438 26444
rect 20993 26367 21051 26373
rect 20993 26364 21005 26367
rect 20824 26336 21005 26364
rect 20717 26327 20775 26333
rect 20993 26333 21005 26336
rect 21039 26333 21051 26367
rect 24394 26364 24400 26376
rect 24355 26336 24400 26364
rect 20993 26327 21051 26333
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 30282 26364 30288 26376
rect 30243 26336 30288 26364
rect 30282 26324 30288 26336
rect 30340 26324 30346 26376
rect 37826 26364 37832 26376
rect 37787 26336 37832 26364
rect 37826 26324 37832 26336
rect 37884 26324 37890 26376
rect 14826 26296 14832 26308
rect 14384 26268 14688 26296
rect 14787 26268 14832 26296
rect 3050 26188 3056 26240
rect 3108 26228 3114 26240
rect 3970 26228 3976 26240
rect 3108 26200 3976 26228
rect 3108 26188 3114 26200
rect 3970 26188 3976 26200
rect 4028 26188 4034 26240
rect 8294 26228 8300 26240
rect 8255 26200 8300 26228
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 14660 26228 14688 26268
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 15654 26296 15660 26308
rect 14936 26268 15660 26296
rect 14936 26228 14964 26268
rect 15654 26256 15660 26268
rect 15712 26256 15718 26308
rect 19426 26256 19432 26308
rect 19484 26296 19490 26308
rect 20622 26296 20628 26308
rect 19484 26268 20628 26296
rect 19484 26256 19490 26268
rect 20622 26256 20628 26268
rect 20680 26256 20686 26308
rect 22186 26296 22192 26308
rect 22147 26268 22192 26296
rect 22186 26256 22192 26268
rect 22244 26256 22250 26308
rect 26234 26256 26240 26308
rect 26292 26296 26298 26308
rect 27801 26299 27859 26305
rect 27801 26296 27813 26299
rect 26292 26268 27813 26296
rect 26292 26256 26298 26268
rect 27801 26265 27813 26268
rect 27847 26265 27859 26299
rect 27801 26259 27859 26265
rect 14660 26200 14964 26228
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 3050 26024 3056 26036
rect 3011 25996 3056 26024
rect 3050 25984 3056 25996
rect 3108 25984 3114 26036
rect 3513 26027 3571 26033
rect 3513 25993 3525 26027
rect 3559 25993 3571 26027
rect 3513 25987 3571 25993
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25888 1458 25900
rect 2041 25891 2099 25897
rect 2041 25888 2053 25891
rect 1452 25860 2053 25888
rect 1452 25848 1458 25860
rect 2041 25857 2053 25860
rect 2087 25857 2099 25891
rect 2041 25851 2099 25857
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25888 2927 25891
rect 3528 25888 3556 25987
rect 3602 25984 3608 26036
rect 3660 26024 3666 26036
rect 24949 26027 25007 26033
rect 3660 25996 22094 26024
rect 3660 25984 3666 25996
rect 3973 25959 4031 25965
rect 3973 25925 3985 25959
rect 4019 25956 4031 25959
rect 4614 25956 4620 25968
rect 4019 25928 4620 25956
rect 4019 25925 4031 25928
rect 3973 25919 4031 25925
rect 4614 25916 4620 25928
rect 4672 25916 4678 25968
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 7009 25959 7067 25965
rect 7009 25956 7021 25959
rect 6972 25928 7021 25956
rect 6972 25916 6978 25928
rect 7009 25925 7021 25928
rect 7055 25925 7067 25959
rect 10778 25956 10784 25968
rect 10691 25928 10784 25956
rect 7009 25919 7067 25925
rect 10778 25916 10784 25928
rect 10836 25956 10842 25968
rect 18230 25956 18236 25968
rect 10836 25928 18236 25956
rect 10836 25916 10842 25928
rect 18230 25916 18236 25928
rect 18288 25916 18294 25968
rect 22066 25956 22094 25996
rect 24949 25993 24961 26027
rect 24995 26024 25007 26027
rect 26234 26024 26240 26036
rect 24995 25996 26240 26024
rect 24995 25993 25007 25996
rect 24949 25987 25007 25993
rect 26234 25984 26240 25996
rect 26292 25984 26298 26036
rect 27709 26027 27767 26033
rect 27709 25993 27721 26027
rect 27755 26024 27767 26027
rect 28074 26024 28080 26036
rect 27755 25996 28080 26024
rect 27755 25993 27767 25996
rect 27709 25987 27767 25993
rect 28074 25984 28080 25996
rect 28132 25984 28138 26036
rect 29362 26024 29368 26036
rect 29323 25996 29368 26024
rect 29362 25984 29368 25996
rect 29420 25984 29426 26036
rect 30374 26024 30380 26036
rect 30335 25996 30380 26024
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 22373 25959 22431 25965
rect 22373 25956 22385 25959
rect 22066 25928 22385 25956
rect 22373 25925 22385 25928
rect 22419 25956 22431 25959
rect 23934 25956 23940 25968
rect 22419 25928 23940 25956
rect 22419 25925 22431 25928
rect 22373 25919 22431 25925
rect 23934 25916 23940 25928
rect 23992 25956 23998 25968
rect 26694 25956 26700 25968
rect 23992 25928 26700 25956
rect 23992 25916 23998 25928
rect 26694 25916 26700 25928
rect 26752 25916 26758 25968
rect 26878 25916 26884 25968
rect 26936 25956 26942 25968
rect 27341 25959 27399 25965
rect 27341 25956 27353 25959
rect 26936 25928 27353 25956
rect 26936 25916 26942 25928
rect 27341 25925 27353 25928
rect 27387 25925 27399 25959
rect 27341 25919 27399 25925
rect 28261 25959 28319 25965
rect 28261 25925 28273 25959
rect 28307 25956 28319 25959
rect 30558 25956 30564 25968
rect 28307 25928 30564 25956
rect 28307 25925 28319 25928
rect 28261 25919 28319 25925
rect 2915 25860 3556 25888
rect 2915 25857 2927 25860
rect 2869 25851 2927 25857
rect 3694 25848 3700 25900
rect 3752 25888 3758 25900
rect 4062 25888 4068 25900
rect 3752 25860 4068 25888
rect 3752 25848 3758 25860
rect 4062 25848 4068 25860
rect 4120 25848 4126 25900
rect 7742 25848 7748 25900
rect 7800 25888 7806 25900
rect 7837 25891 7895 25897
rect 7837 25888 7849 25891
rect 7800 25860 7849 25888
rect 7800 25848 7806 25860
rect 7837 25857 7849 25860
rect 7883 25888 7895 25891
rect 7926 25888 7932 25900
rect 7883 25860 7932 25888
rect 7883 25857 7895 25860
rect 7837 25851 7895 25857
rect 7926 25848 7932 25860
rect 7984 25848 7990 25900
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25888 8171 25891
rect 8202 25888 8208 25900
rect 8159 25860 8208 25888
rect 8159 25857 8171 25860
rect 8113 25851 8171 25857
rect 8202 25848 8208 25860
rect 8260 25848 8266 25900
rect 12066 25888 12072 25900
rect 12027 25860 12072 25888
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 14734 25848 14740 25900
rect 14792 25888 14798 25900
rect 15105 25891 15163 25897
rect 15105 25888 15117 25891
rect 14792 25860 15117 25888
rect 14792 25848 14798 25860
rect 15105 25857 15117 25860
rect 15151 25857 15163 25891
rect 15746 25888 15752 25900
rect 15707 25860 15752 25888
rect 15105 25851 15163 25857
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 17954 25888 17960 25900
rect 17915 25860 17960 25888
rect 17954 25848 17960 25860
rect 18012 25848 18018 25900
rect 24213 25891 24271 25897
rect 24213 25857 24225 25891
rect 24259 25888 24271 25891
rect 24394 25888 24400 25900
rect 24259 25860 24400 25888
rect 24259 25857 24271 25860
rect 24213 25851 24271 25857
rect 24394 25848 24400 25860
rect 24452 25848 24458 25900
rect 24765 25891 24823 25897
rect 24765 25857 24777 25891
rect 24811 25857 24823 25891
rect 24765 25851 24823 25857
rect 25685 25891 25743 25897
rect 25685 25857 25697 25891
rect 25731 25888 25743 25891
rect 27154 25888 27160 25900
rect 25731 25860 27160 25888
rect 25731 25857 25743 25860
rect 25685 25851 25743 25857
rect 3881 25823 3939 25829
rect 3881 25789 3893 25823
rect 3927 25820 3939 25823
rect 4798 25820 4804 25832
rect 3927 25792 4804 25820
rect 3927 25789 3939 25792
rect 3881 25783 3939 25789
rect 4798 25780 4804 25792
rect 4856 25780 4862 25832
rect 8018 25820 8024 25832
rect 7979 25792 8024 25820
rect 8018 25780 8024 25792
rect 8076 25780 8082 25832
rect 8941 25823 8999 25829
rect 8941 25789 8953 25823
rect 8987 25789 8999 25823
rect 9122 25820 9128 25832
rect 9083 25792 9128 25820
rect 8941 25783 8999 25789
rect 8956 25752 8984 25783
rect 9122 25780 9128 25792
rect 9180 25780 9186 25832
rect 12253 25823 12311 25829
rect 12253 25789 12265 25823
rect 12299 25820 12311 25823
rect 13262 25820 13268 25832
rect 12299 25792 13268 25820
rect 12299 25789 12311 25792
rect 12253 25783 12311 25789
rect 13262 25780 13268 25792
rect 13320 25780 13326 25832
rect 13446 25820 13452 25832
rect 13407 25792 13452 25820
rect 13446 25780 13452 25792
rect 13504 25820 13510 25832
rect 13504 25792 16574 25820
rect 13504 25780 13510 25792
rect 9582 25752 9588 25764
rect 8956 25724 9588 25752
rect 9582 25712 9588 25724
rect 9640 25712 9646 25764
rect 14921 25755 14979 25761
rect 14921 25721 14933 25755
rect 14967 25752 14979 25755
rect 15010 25752 15016 25764
rect 14967 25724 15016 25752
rect 14967 25721 14979 25724
rect 14921 25715 14979 25721
rect 15010 25712 15016 25724
rect 15068 25712 15074 25764
rect 15562 25752 15568 25764
rect 15523 25724 15568 25752
rect 15562 25712 15568 25724
rect 15620 25712 15626 25764
rect 16546 25752 16574 25792
rect 17678 25780 17684 25832
rect 17736 25820 17742 25832
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 17736 25792 18153 25820
rect 17736 25780 17742 25792
rect 18141 25789 18153 25792
rect 18187 25789 18199 25823
rect 19426 25820 19432 25832
rect 19387 25792 19432 25820
rect 18141 25783 18199 25789
rect 19426 25780 19432 25792
rect 19484 25780 19490 25832
rect 22554 25780 22560 25832
rect 22612 25820 22618 25832
rect 24029 25823 24087 25829
rect 24029 25820 24041 25823
rect 22612 25792 24041 25820
rect 22612 25780 22618 25792
rect 24029 25789 24041 25792
rect 24075 25789 24087 25823
rect 24029 25783 24087 25789
rect 24302 25780 24308 25832
rect 24360 25820 24366 25832
rect 24780 25820 24808 25851
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 27249 25891 27307 25897
rect 27249 25857 27261 25891
rect 27295 25888 27307 25891
rect 28276 25888 28304 25919
rect 30558 25916 30564 25928
rect 30616 25956 30622 25968
rect 31294 25956 31300 25968
rect 30616 25928 31300 25956
rect 30616 25916 30622 25928
rect 31294 25916 31300 25928
rect 31352 25916 31358 25968
rect 27295 25860 28304 25888
rect 27295 25857 27307 25860
rect 27249 25851 27307 25857
rect 29362 25848 29368 25900
rect 29420 25888 29426 25900
rect 30285 25891 30343 25897
rect 30285 25888 30297 25891
rect 29420 25860 30297 25888
rect 29420 25848 29426 25860
rect 30285 25857 30297 25860
rect 30331 25857 30343 25891
rect 34330 25888 34336 25900
rect 34291 25860 34336 25888
rect 30285 25851 30343 25857
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 34422 25848 34428 25900
rect 34480 25888 34486 25900
rect 34609 25891 34667 25897
rect 34480 25860 34525 25888
rect 34480 25848 34486 25860
rect 34609 25857 34621 25891
rect 34655 25857 34667 25891
rect 34609 25851 34667 25857
rect 25406 25820 25412 25832
rect 24360 25792 24808 25820
rect 25367 25792 25412 25820
rect 24360 25780 24366 25792
rect 25406 25780 25412 25792
rect 25464 25780 25470 25832
rect 27062 25820 27068 25832
rect 27023 25792 27068 25820
rect 27062 25780 27068 25792
rect 27120 25780 27126 25832
rect 30469 25823 30527 25829
rect 30469 25789 30481 25823
rect 30515 25789 30527 25823
rect 34624 25820 34652 25851
rect 34698 25848 34704 25900
rect 34756 25888 34762 25900
rect 35161 25891 35219 25897
rect 35161 25888 35173 25891
rect 34756 25860 35173 25888
rect 34756 25848 34762 25860
rect 35161 25857 35173 25860
rect 35207 25857 35219 25891
rect 35161 25851 35219 25857
rect 35345 25891 35403 25897
rect 35345 25857 35357 25891
rect 35391 25888 35403 25891
rect 35894 25888 35900 25900
rect 35391 25860 35900 25888
rect 35391 25857 35403 25860
rect 35345 25851 35403 25857
rect 35894 25848 35900 25860
rect 35952 25848 35958 25900
rect 35253 25823 35311 25829
rect 35253 25820 35265 25823
rect 34624 25792 35265 25820
rect 30469 25783 30527 25789
rect 35253 25789 35265 25792
rect 35299 25789 35311 25823
rect 35253 25783 35311 25789
rect 23382 25752 23388 25764
rect 16546 25724 23388 25752
rect 23382 25712 23388 25724
rect 23440 25712 23446 25764
rect 29086 25712 29092 25764
rect 29144 25752 29150 25764
rect 30484 25752 30512 25783
rect 29144 25724 30512 25752
rect 29144 25712 29150 25724
rect 33594 25712 33600 25764
rect 33652 25752 33658 25764
rect 33689 25755 33747 25761
rect 33689 25752 33701 25755
rect 33652 25724 33701 25752
rect 33652 25712 33658 25724
rect 33689 25721 33701 25724
rect 33735 25752 33747 25755
rect 34517 25755 34575 25761
rect 34517 25752 34529 25755
rect 33735 25724 34529 25752
rect 33735 25721 33747 25724
rect 33689 25715 33747 25721
rect 34517 25721 34529 25724
rect 34563 25752 34575 25755
rect 34606 25752 34612 25764
rect 34563 25724 34612 25752
rect 34563 25721 34575 25724
rect 34517 25715 34575 25721
rect 34606 25712 34612 25724
rect 34664 25712 34670 25764
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 2866 25684 2872 25696
rect 1627 25656 2872 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 2866 25644 2872 25656
rect 2924 25644 2930 25696
rect 3881 25687 3939 25693
rect 3881 25653 3893 25687
rect 3927 25684 3939 25687
rect 4706 25684 4712 25696
rect 3927 25656 4712 25684
rect 3927 25653 3939 25656
rect 3881 25647 3939 25653
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 7834 25684 7840 25696
rect 7795 25656 7840 25684
rect 7834 25644 7840 25656
rect 7892 25644 7898 25696
rect 8297 25687 8355 25693
rect 8297 25653 8309 25687
rect 8343 25684 8355 25687
rect 10042 25684 10048 25696
rect 8343 25656 10048 25684
rect 8343 25653 8355 25656
rect 8297 25647 8355 25653
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 29917 25687 29975 25693
rect 29917 25653 29929 25687
rect 29963 25684 29975 25687
rect 30098 25684 30104 25696
rect 29963 25656 30104 25684
rect 29963 25653 29975 25656
rect 29917 25647 29975 25653
rect 30098 25644 30104 25656
rect 30156 25644 30162 25696
rect 34146 25684 34152 25696
rect 34107 25656 34152 25684
rect 34146 25644 34152 25656
rect 34204 25644 34210 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1578 25440 1584 25492
rect 1636 25480 1642 25492
rect 2501 25483 2559 25489
rect 2501 25480 2513 25483
rect 1636 25452 2513 25480
rect 1636 25440 1642 25452
rect 2501 25449 2513 25452
rect 2547 25449 2559 25483
rect 2501 25443 2559 25449
rect 4065 25483 4123 25489
rect 4065 25449 4077 25483
rect 4111 25480 4123 25483
rect 4706 25480 4712 25492
rect 4111 25452 4712 25480
rect 4111 25449 4123 25452
rect 4065 25443 4123 25449
rect 4706 25440 4712 25452
rect 4764 25440 4770 25492
rect 9122 25480 9128 25492
rect 9083 25452 9128 25480
rect 9122 25440 9128 25452
rect 9180 25440 9186 25492
rect 9582 25480 9588 25492
rect 9543 25452 9588 25480
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 14918 25480 14924 25492
rect 14507 25452 14924 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 14918 25440 14924 25452
rect 14976 25440 14982 25492
rect 15194 25480 15200 25492
rect 15155 25452 15200 25480
rect 15194 25440 15200 25452
rect 15252 25440 15258 25492
rect 17678 25480 17684 25492
rect 17639 25452 17684 25480
rect 17678 25440 17684 25452
rect 17736 25440 17742 25492
rect 21913 25483 21971 25489
rect 21913 25449 21925 25483
rect 21959 25480 21971 25483
rect 22186 25480 22192 25492
rect 21959 25452 22192 25480
rect 21959 25449 21971 25452
rect 21913 25443 21971 25449
rect 22186 25440 22192 25452
rect 22244 25440 22250 25492
rect 22554 25480 22560 25492
rect 22515 25452 22560 25480
rect 22554 25440 22560 25452
rect 22612 25440 22618 25492
rect 23661 25483 23719 25489
rect 23661 25449 23673 25483
rect 23707 25480 23719 25483
rect 23750 25480 23756 25492
rect 23707 25452 23756 25480
rect 23707 25449 23719 25452
rect 23661 25443 23719 25449
rect 23750 25440 23756 25452
rect 23808 25440 23814 25492
rect 23845 25483 23903 25489
rect 23845 25449 23857 25483
rect 23891 25480 23903 25483
rect 24302 25480 24308 25492
rect 23891 25452 24308 25480
rect 23891 25449 23903 25452
rect 23845 25443 23903 25449
rect 24302 25440 24308 25452
rect 24360 25440 24366 25492
rect 24397 25483 24455 25489
rect 24397 25449 24409 25483
rect 24443 25449 24455 25483
rect 30282 25480 30288 25492
rect 30243 25452 30288 25480
rect 24397 25443 24455 25449
rect 23768 25412 23796 25440
rect 24412 25412 24440 25443
rect 30282 25440 30288 25452
rect 30340 25440 30346 25492
rect 23768 25384 24440 25412
rect 2774 25344 2780 25356
rect 2735 25316 2780 25344
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 3973 25347 4031 25353
rect 3973 25313 3985 25347
rect 4019 25344 4031 25347
rect 4798 25344 4804 25356
rect 4019 25316 4804 25344
rect 4019 25313 4031 25316
rect 3973 25307 4031 25313
rect 4798 25304 4804 25316
rect 4856 25304 4862 25356
rect 15286 25344 15292 25356
rect 15247 25316 15292 25344
rect 15286 25304 15292 25316
rect 15344 25304 15350 25356
rect 24486 25344 24492 25356
rect 24447 25316 24492 25344
rect 24486 25304 24492 25316
rect 24544 25304 24550 25356
rect 1946 25276 1952 25288
rect 1907 25248 1952 25276
rect 1946 25236 1952 25248
rect 2004 25236 2010 25288
rect 2866 25276 2872 25288
rect 2827 25248 2872 25276
rect 2866 25236 2872 25248
rect 2924 25236 2930 25288
rect 4062 25276 4068 25288
rect 4023 25248 4068 25276
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4264 25248 4905 25276
rect 2406 25208 2412 25220
rect 2367 25180 2412 25208
rect 2406 25168 2412 25180
rect 2464 25168 2470 25220
rect 3789 25211 3847 25217
rect 3789 25177 3801 25211
rect 3835 25208 3847 25211
rect 3878 25208 3884 25220
rect 3835 25180 3884 25208
rect 3835 25177 3847 25180
rect 3789 25171 3847 25177
rect 3878 25168 3884 25180
rect 3936 25168 3942 25220
rect 3050 25140 3056 25152
rect 3011 25112 3056 25140
rect 3050 25100 3056 25112
rect 3108 25100 3114 25152
rect 4264 25149 4292 25248
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 4893 25239 4951 25245
rect 7650 25236 7656 25288
rect 7708 25276 7714 25288
rect 7926 25276 7932 25288
rect 7708 25248 7932 25276
rect 7708 25236 7714 25248
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8352 25248 8953 25276
rect 8352 25236 8358 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 14642 25276 14648 25288
rect 14323 25248 14648 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 14642 25236 14648 25248
rect 14700 25236 14706 25288
rect 15010 25236 15016 25288
rect 15068 25276 15074 25288
rect 15378 25276 15384 25288
rect 15068 25248 15384 25276
rect 15068 25236 15074 25248
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 16853 25279 16911 25285
rect 16853 25276 16865 25279
rect 16546 25248 16865 25276
rect 14826 25168 14832 25220
rect 14884 25208 14890 25220
rect 15105 25211 15163 25217
rect 15105 25208 15117 25211
rect 14884 25180 15117 25208
rect 14884 25168 14890 25180
rect 15105 25177 15117 25180
rect 15151 25177 15163 25211
rect 15105 25171 15163 25177
rect 4249 25143 4307 25149
rect 4249 25109 4261 25143
rect 4295 25109 4307 25143
rect 4249 25103 4307 25109
rect 4338 25100 4344 25152
rect 4396 25140 4402 25152
rect 4709 25143 4767 25149
rect 4709 25140 4721 25143
rect 4396 25112 4721 25140
rect 4396 25100 4402 25112
rect 4709 25109 4721 25112
rect 4755 25109 4767 25143
rect 7742 25140 7748 25152
rect 7703 25112 7748 25140
rect 4709 25103 4767 25109
rect 7742 25100 7748 25112
rect 7800 25100 7806 25152
rect 15565 25143 15623 25149
rect 15565 25109 15577 25143
rect 15611 25140 15623 25143
rect 16546 25140 16574 25248
rect 16853 25245 16865 25248
rect 16899 25245 16911 25279
rect 17494 25276 17500 25288
rect 17455 25248 17500 25276
rect 16853 25239 16911 25245
rect 17494 25236 17500 25248
rect 17552 25236 17558 25288
rect 18138 25276 18144 25288
rect 18099 25248 18144 25276
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 21726 25276 21732 25288
rect 21687 25248 21732 25276
rect 21726 25236 21732 25248
rect 21784 25236 21790 25288
rect 22094 25236 22100 25288
rect 22152 25276 22158 25288
rect 22373 25279 22431 25285
rect 22373 25276 22385 25279
rect 22152 25248 22385 25276
rect 22152 25236 22158 25248
rect 22373 25245 22385 25248
rect 22419 25245 22431 25279
rect 23566 25276 23572 25288
rect 23527 25248 23572 25276
rect 22373 25239 22431 25245
rect 23566 25236 23572 25248
rect 23624 25236 23630 25288
rect 23658 25236 23664 25288
rect 23716 25276 23722 25288
rect 24026 25276 24032 25288
rect 23716 25248 24032 25276
rect 23716 25236 23722 25248
rect 24026 25236 24032 25248
rect 24084 25276 24090 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24084 25248 24685 25276
rect 24084 25236 24090 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 29914 25276 29920 25288
rect 29875 25248 29920 25276
rect 24673 25239 24731 25245
rect 29914 25236 29920 25248
rect 29972 25236 29978 25288
rect 30098 25276 30104 25288
rect 30059 25248 30104 25276
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 23385 25211 23443 25217
rect 23385 25177 23397 25211
rect 23431 25208 23443 25211
rect 23474 25208 23480 25220
rect 23431 25180 23480 25208
rect 23431 25177 23443 25180
rect 23385 25171 23443 25177
rect 23474 25168 23480 25180
rect 23532 25168 23538 25220
rect 23584 25208 23612 25236
rect 24397 25211 24455 25217
rect 24397 25208 24409 25211
rect 23584 25180 24409 25208
rect 24397 25177 24409 25180
rect 24443 25177 24455 25211
rect 24397 25171 24455 25177
rect 15611 25112 16574 25140
rect 17037 25143 17095 25149
rect 15611 25109 15623 25112
rect 15565 25103 15623 25109
rect 17037 25109 17049 25143
rect 17083 25140 17095 25143
rect 17862 25140 17868 25152
rect 17083 25112 17868 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17862 25100 17868 25112
rect 17920 25100 17926 25152
rect 24857 25143 24915 25149
rect 24857 25109 24869 25143
rect 24903 25140 24915 25143
rect 25590 25140 25596 25152
rect 24903 25112 25596 25140
rect 24903 25109 24915 25112
rect 24857 25103 24915 25109
rect 25590 25100 25596 25112
rect 25648 25100 25654 25152
rect 26878 25140 26884 25152
rect 26839 25112 26884 25140
rect 26878 25100 26884 25112
rect 26936 25100 26942 25152
rect 27062 25100 27068 25152
rect 27120 25140 27126 25152
rect 27433 25143 27491 25149
rect 27433 25140 27445 25143
rect 27120 25112 27445 25140
rect 27120 25100 27126 25112
rect 27433 25109 27445 25112
rect 27479 25140 27491 25143
rect 27798 25140 27804 25152
rect 27479 25112 27804 25140
rect 27479 25109 27491 25112
rect 27433 25103 27491 25109
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 8018 24936 8024 24948
rect 7979 24908 8024 24936
rect 8018 24896 8024 24908
rect 8076 24896 8082 24948
rect 29086 24936 29092 24948
rect 29047 24908 29092 24936
rect 29086 24896 29092 24908
rect 29144 24896 29150 24948
rect 14826 24828 14832 24880
rect 14884 24868 14890 24880
rect 15105 24871 15163 24877
rect 15105 24868 15117 24871
rect 14884 24840 15117 24868
rect 14884 24828 14890 24840
rect 15105 24837 15117 24840
rect 15151 24837 15163 24871
rect 17862 24868 17868 24880
rect 17823 24840 17868 24868
rect 15105 24831 15163 24837
rect 17862 24828 17868 24840
rect 17920 24828 17926 24880
rect 23658 24828 23664 24880
rect 23716 24868 23722 24880
rect 24486 24868 24492 24880
rect 23716 24840 24492 24868
rect 23716 24828 23722 24840
rect 24486 24828 24492 24840
rect 24544 24868 24550 24880
rect 24673 24871 24731 24877
rect 24673 24868 24685 24871
rect 24544 24840 24685 24868
rect 24544 24828 24550 24840
rect 24673 24837 24685 24840
rect 24719 24837 24731 24871
rect 24673 24831 24731 24837
rect 1946 24760 1952 24812
rect 2004 24800 2010 24812
rect 2685 24803 2743 24809
rect 2685 24800 2697 24803
rect 2004 24772 2697 24800
rect 2004 24760 2010 24772
rect 2685 24769 2697 24772
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4525 24803 4583 24809
rect 4525 24800 4537 24803
rect 4120 24772 4537 24800
rect 4120 24760 4126 24772
rect 4525 24769 4537 24772
rect 4571 24769 4583 24803
rect 4525 24763 4583 24769
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24800 5227 24803
rect 5810 24800 5816 24812
rect 5215 24772 5816 24800
rect 5215 24769 5227 24772
rect 5169 24763 5227 24769
rect 2869 24735 2927 24741
rect 2869 24701 2881 24735
rect 2915 24732 2927 24735
rect 4338 24732 4344 24744
rect 2915 24704 4344 24732
rect 2915 24701 2927 24704
rect 2869 24695 2927 24701
rect 4338 24692 4344 24704
rect 4396 24692 4402 24744
rect 4540 24732 4568 24763
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 7834 24800 7840 24812
rect 7795 24772 7840 24800
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 13262 24800 13268 24812
rect 13223 24772 13268 24800
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 15378 24800 15384 24812
rect 15339 24772 15384 24800
rect 15378 24760 15384 24772
rect 15436 24760 15442 24812
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 23474 24800 23480 24812
rect 23072 24772 23480 24800
rect 23072 24760 23078 24772
rect 23474 24760 23480 24772
rect 23532 24800 23538 24812
rect 23753 24803 23811 24809
rect 23753 24800 23765 24803
rect 23532 24772 23765 24800
rect 23532 24760 23538 24772
rect 23753 24769 23765 24772
rect 23799 24769 23811 24803
rect 24026 24800 24032 24812
rect 23987 24772 24032 24800
rect 23753 24763 23811 24769
rect 24026 24760 24032 24772
rect 24084 24760 24090 24812
rect 28905 24803 28963 24809
rect 28905 24800 28917 24803
rect 28368 24772 28917 24800
rect 10778 24732 10784 24744
rect 4540 24704 10784 24732
rect 10778 24692 10784 24704
rect 10836 24692 10842 24744
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24732 13599 24735
rect 13906 24732 13912 24744
rect 13587 24704 13912 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 15286 24732 15292 24744
rect 15247 24704 15292 24732
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 17681 24735 17739 24741
rect 17681 24701 17693 24735
rect 17727 24701 17739 24735
rect 18230 24732 18236 24744
rect 18191 24704 18236 24732
rect 17681 24695 17739 24701
rect 4798 24624 4804 24676
rect 4856 24664 4862 24676
rect 4985 24667 5043 24673
rect 4985 24664 4997 24667
rect 4856 24636 4997 24664
rect 4856 24624 4862 24636
rect 4985 24633 4997 24636
rect 5031 24633 5043 24667
rect 4985 24627 5043 24633
rect 7834 24624 7840 24676
rect 7892 24664 7898 24676
rect 8573 24667 8631 24673
rect 8573 24664 8585 24667
rect 7892 24636 8585 24664
rect 7892 24624 7898 24636
rect 8573 24633 8585 24636
rect 8619 24664 8631 24667
rect 15378 24664 15384 24676
rect 8619 24636 15384 24664
rect 8619 24633 8631 24636
rect 8573 24627 8631 24633
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 15565 24667 15623 24673
rect 15565 24633 15577 24667
rect 15611 24664 15623 24667
rect 17494 24664 17500 24676
rect 15611 24636 17500 24664
rect 15611 24633 15623 24636
rect 15565 24627 15623 24633
rect 17494 24624 17500 24636
rect 17552 24624 17558 24676
rect 17696 24664 17724 24695
rect 18230 24692 18236 24704
rect 18288 24692 18294 24744
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24701 23903 24735
rect 23845 24695 23903 24701
rect 18138 24664 18144 24676
rect 17696 24636 18144 24664
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 23474 24624 23480 24676
rect 23532 24664 23538 24676
rect 23860 24664 23888 24695
rect 23532 24636 23888 24664
rect 24213 24667 24271 24673
rect 23532 24624 23538 24636
rect 24213 24633 24225 24667
rect 24259 24664 24271 24667
rect 25406 24664 25412 24676
rect 24259 24636 25412 24664
rect 24259 24633 24271 24636
rect 24213 24627 24271 24633
rect 25406 24624 25412 24636
rect 25464 24624 25470 24676
rect 5810 24596 5816 24608
rect 5723 24568 5816 24596
rect 5810 24556 5816 24568
rect 5868 24596 5874 24608
rect 6270 24596 6276 24608
rect 5868 24568 6276 24596
rect 5868 24556 5874 24568
rect 6270 24556 6276 24568
rect 6328 24596 6334 24608
rect 6914 24596 6920 24608
rect 6328 24568 6920 24596
rect 6328 24556 6334 24568
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 15194 24596 15200 24608
rect 15155 24568 15200 24596
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 23750 24596 23756 24608
rect 23711 24568 23756 24596
rect 23750 24556 23756 24568
rect 23808 24556 23814 24608
rect 27798 24556 27804 24608
rect 27856 24596 27862 24608
rect 28368 24605 28396 24772
rect 28905 24769 28917 24772
rect 28951 24769 28963 24803
rect 28905 24763 28963 24769
rect 30190 24760 30196 24812
rect 30248 24800 30254 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 30248 24772 30573 24800
rect 30248 24760 30254 24772
rect 30561 24769 30573 24772
rect 30607 24769 30619 24803
rect 30561 24763 30619 24769
rect 35897 24803 35955 24809
rect 35897 24769 35909 24803
rect 35943 24769 35955 24803
rect 35897 24763 35955 24769
rect 35989 24803 36047 24809
rect 35989 24769 36001 24803
rect 36035 24800 36047 24803
rect 36078 24800 36084 24812
rect 36035 24772 36084 24800
rect 36035 24769 36047 24772
rect 35989 24763 36047 24769
rect 35912 24676 35940 24763
rect 36078 24760 36084 24772
rect 36136 24760 36142 24812
rect 36262 24800 36268 24812
rect 36223 24772 36268 24800
rect 36262 24760 36268 24772
rect 36320 24760 36326 24812
rect 35894 24624 35900 24676
rect 35952 24624 35958 24676
rect 28353 24599 28411 24605
rect 28353 24596 28365 24599
rect 27856 24568 28365 24596
rect 27856 24556 27862 24568
rect 28353 24565 28365 24568
rect 28399 24565 28411 24599
rect 28353 24559 28411 24565
rect 30745 24599 30803 24605
rect 30745 24565 30757 24599
rect 30791 24596 30803 24599
rect 30926 24596 30932 24608
rect 30791 24568 30932 24596
rect 30791 24565 30803 24568
rect 30745 24559 30803 24565
rect 30926 24556 30932 24568
rect 30984 24556 30990 24608
rect 34790 24596 34796 24608
rect 34751 24568 34796 24596
rect 34790 24556 34796 24568
rect 34848 24556 34854 24608
rect 35710 24596 35716 24608
rect 35671 24568 35716 24596
rect 35710 24556 35716 24568
rect 35768 24556 35774 24608
rect 36173 24599 36231 24605
rect 36173 24565 36185 24599
rect 36219 24596 36231 24599
rect 37366 24596 37372 24608
rect 36219 24568 37372 24596
rect 36219 24565 36231 24568
rect 36173 24559 36231 24565
rect 37366 24556 37372 24568
rect 37424 24556 37430 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1581 24395 1639 24401
rect 1581 24361 1593 24395
rect 1627 24392 1639 24395
rect 2406 24392 2412 24404
rect 1627 24364 2412 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 2406 24352 2412 24364
rect 2464 24352 2470 24404
rect 14461 24395 14519 24401
rect 14461 24361 14473 24395
rect 14507 24392 14519 24395
rect 15286 24392 15292 24404
rect 14507 24364 15292 24392
rect 14507 24361 14519 24364
rect 14461 24355 14519 24361
rect 15286 24352 15292 24364
rect 15344 24352 15350 24404
rect 15378 24352 15384 24404
rect 15436 24392 15442 24404
rect 22094 24392 22100 24404
rect 15436 24364 22100 24392
rect 15436 24352 15442 24364
rect 22094 24352 22100 24364
rect 22152 24352 22158 24404
rect 30190 24392 30196 24404
rect 30151 24364 30196 24392
rect 30190 24352 30196 24364
rect 30248 24352 30254 24404
rect 14826 24284 14832 24336
rect 14884 24324 14890 24336
rect 15105 24327 15163 24333
rect 15105 24324 15117 24327
rect 14884 24296 15117 24324
rect 14884 24284 14890 24296
rect 15105 24293 15117 24296
rect 15151 24293 15163 24327
rect 15105 24287 15163 24293
rect 28997 24327 29055 24333
rect 28997 24293 29009 24327
rect 29043 24324 29055 24327
rect 30466 24324 30472 24336
rect 29043 24296 30472 24324
rect 29043 24293 29055 24296
rect 28997 24287 29055 24293
rect 30466 24284 30472 24296
rect 30524 24284 30530 24336
rect 36170 24324 36176 24336
rect 32232 24296 36176 24324
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24188 1458 24200
rect 2041 24191 2099 24197
rect 2041 24188 2053 24191
rect 1452 24160 2053 24188
rect 1452 24148 1458 24160
rect 2041 24157 2053 24160
rect 2087 24157 2099 24191
rect 2041 24151 2099 24157
rect 7190 24148 7196 24200
rect 7248 24188 7254 24200
rect 7285 24191 7343 24197
rect 7285 24188 7297 24191
rect 7248 24160 7297 24188
rect 7248 24148 7254 24160
rect 7285 24157 7297 24160
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 14090 24188 14096 24200
rect 12851 24160 14096 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14642 24188 14648 24200
rect 14603 24160 14648 24188
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 15289 24191 15347 24197
rect 15289 24188 15301 24191
rect 15252 24160 15301 24188
rect 15252 24148 15258 24160
rect 15289 24157 15301 24160
rect 15335 24188 15347 24191
rect 15746 24188 15752 24200
rect 15335 24160 15752 24188
rect 15335 24157 15347 24160
rect 15289 24151 15347 24157
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 20438 24188 20444 24200
rect 19475 24160 20444 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 29914 24188 29920 24200
rect 29875 24160 29920 24188
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24188 30067 24191
rect 30282 24188 30288 24200
rect 30055 24160 30288 24188
rect 30055 24157 30067 24160
rect 30009 24151 30067 24157
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30834 24188 30840 24200
rect 30795 24160 30840 24188
rect 30834 24148 30840 24160
rect 30892 24148 30898 24200
rect 30926 24148 30932 24200
rect 30984 24188 30990 24200
rect 31093 24191 31151 24197
rect 31093 24188 31105 24191
rect 30984 24160 31105 24188
rect 30984 24148 30990 24160
rect 31093 24157 31105 24160
rect 31139 24157 31151 24191
rect 31093 24151 31151 24157
rect 28810 24120 28816 24132
rect 28771 24092 28816 24120
rect 28810 24080 28816 24092
rect 28868 24080 28874 24132
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 12621 24055 12679 24061
rect 12621 24052 12633 24055
rect 11848 24024 12633 24052
rect 11848 24012 11854 24024
rect 12621 24021 12633 24024
rect 12667 24021 12679 24055
rect 12621 24015 12679 24021
rect 22094 24012 22100 24064
rect 22152 24052 22158 24064
rect 22152 24024 22197 24052
rect 22152 24012 22158 24024
rect 29822 24012 29828 24064
rect 29880 24052 29886 24064
rect 32232 24061 32260 24296
rect 36170 24284 36176 24296
rect 36228 24284 36234 24336
rect 36081 24259 36139 24265
rect 36081 24225 36093 24259
rect 36127 24256 36139 24259
rect 36725 24259 36783 24265
rect 36725 24256 36737 24259
rect 36127 24228 36737 24256
rect 36127 24225 36139 24228
rect 36081 24219 36139 24225
rect 36725 24225 36737 24228
rect 36771 24225 36783 24259
rect 36725 24219 36783 24225
rect 33045 24191 33103 24197
rect 33045 24157 33057 24191
rect 33091 24157 33103 24191
rect 33045 24151 33103 24157
rect 33229 24191 33287 24197
rect 33229 24157 33241 24191
rect 33275 24188 33287 24191
rect 34146 24188 34152 24200
rect 33275 24160 34152 24188
rect 33275 24157 33287 24160
rect 33229 24151 33287 24157
rect 33060 24120 33088 24151
rect 34146 24148 34152 24160
rect 34204 24148 34210 24200
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34977 24191 35035 24197
rect 34977 24188 34989 24191
rect 34848 24160 34989 24188
rect 34848 24148 34854 24160
rect 34977 24157 34989 24160
rect 35023 24157 35035 24191
rect 34977 24151 35035 24157
rect 35161 24191 35219 24197
rect 35161 24157 35173 24191
rect 35207 24188 35219 24191
rect 35710 24188 35716 24200
rect 35207 24160 35716 24188
rect 35207 24157 35219 24160
rect 35161 24151 35219 24157
rect 35710 24148 35716 24160
rect 35768 24148 35774 24200
rect 35805 24191 35863 24197
rect 35805 24157 35817 24191
rect 35851 24157 35863 24191
rect 35805 24151 35863 24157
rect 35897 24191 35955 24197
rect 35897 24157 35909 24191
rect 35943 24188 35955 24191
rect 36173 24191 36231 24197
rect 35943 24160 36032 24188
rect 35943 24157 35955 24160
rect 35897 24151 35955 24157
rect 33781 24123 33839 24129
rect 33781 24120 33793 24123
rect 33060 24092 33793 24120
rect 33781 24089 33793 24092
rect 33827 24120 33839 24123
rect 34808 24120 34836 24148
rect 33827 24092 34836 24120
rect 33827 24089 33839 24092
rect 33781 24083 33839 24089
rect 34882 24080 34888 24132
rect 34940 24120 34946 24132
rect 35621 24123 35679 24129
rect 35621 24120 35633 24123
rect 34940 24092 35633 24120
rect 34940 24080 34946 24092
rect 35621 24089 35633 24092
rect 35667 24089 35679 24123
rect 35621 24083 35679 24089
rect 32217 24055 32275 24061
rect 32217 24052 32229 24055
rect 29880 24024 32229 24052
rect 29880 24012 29886 24024
rect 32217 24021 32229 24024
rect 32263 24021 32275 24055
rect 32217 24015 32275 24021
rect 32490 24012 32496 24064
rect 32548 24052 32554 24064
rect 33137 24055 33195 24061
rect 33137 24052 33149 24055
rect 32548 24024 33149 24052
rect 32548 24012 32554 24024
rect 33137 24021 33149 24024
rect 33183 24021 33195 24055
rect 33137 24015 33195 24021
rect 35069 24055 35127 24061
rect 35069 24021 35081 24055
rect 35115 24052 35127 24055
rect 35526 24052 35532 24064
rect 35115 24024 35532 24052
rect 35115 24021 35127 24024
rect 35069 24015 35127 24021
rect 35526 24012 35532 24024
rect 35584 24012 35590 24064
rect 35820 24052 35848 24151
rect 36004 24120 36032 24160
rect 36173 24157 36185 24191
rect 36219 24188 36231 24191
rect 36262 24188 36268 24200
rect 36219 24160 36268 24188
rect 36219 24157 36231 24160
rect 36173 24151 36231 24157
rect 36262 24148 36268 24160
rect 36320 24148 36326 24200
rect 36814 24188 36820 24200
rect 36775 24160 36820 24188
rect 36814 24148 36820 24160
rect 36872 24148 36878 24200
rect 36078 24120 36084 24132
rect 35991 24092 36084 24120
rect 36078 24080 36084 24092
rect 36136 24120 36142 24132
rect 36998 24120 37004 24132
rect 36136 24092 37004 24120
rect 36136 24080 36142 24092
rect 36998 24080 37004 24092
rect 37056 24080 37062 24132
rect 37274 24052 37280 24064
rect 35820 24024 37280 24052
rect 37274 24012 37280 24024
rect 37332 24012 37338 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 13906 23848 13912 23860
rect 13867 23820 13912 23848
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 28994 23848 29000 23860
rect 28955 23820 29000 23848
rect 28994 23808 29000 23820
rect 29052 23848 29058 23860
rect 29917 23851 29975 23857
rect 29917 23848 29929 23851
rect 29052 23820 29929 23848
rect 29052 23808 29058 23820
rect 29917 23817 29929 23820
rect 29963 23817 29975 23851
rect 30282 23848 30288 23860
rect 30243 23820 30288 23848
rect 29917 23811 29975 23817
rect 30282 23808 30288 23820
rect 30340 23808 30346 23860
rect 37366 23848 37372 23860
rect 37327 23820 37372 23848
rect 37366 23808 37372 23820
rect 37424 23808 37430 23860
rect 7098 23780 7104 23792
rect 6886 23752 7104 23780
rect 6365 23715 6423 23721
rect 6365 23681 6377 23715
rect 6411 23712 6423 23715
rect 6886 23712 6914 23752
rect 7098 23740 7104 23752
rect 7156 23740 7162 23792
rect 11790 23780 11796 23792
rect 11751 23752 11796 23780
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 13170 23740 13176 23792
rect 13228 23780 13234 23792
rect 14369 23783 14427 23789
rect 14369 23780 14381 23783
rect 13228 23752 14381 23780
rect 13228 23740 13234 23752
rect 14369 23749 14381 23752
rect 14415 23749 14427 23783
rect 14826 23780 14832 23792
rect 14787 23752 14832 23780
rect 14369 23743 14427 23749
rect 14826 23740 14832 23752
rect 14884 23740 14890 23792
rect 18230 23740 18236 23792
rect 18288 23780 18294 23792
rect 18601 23783 18659 23789
rect 18601 23780 18613 23783
rect 18288 23752 18613 23780
rect 18288 23740 18294 23752
rect 18601 23749 18613 23752
rect 18647 23749 18659 23783
rect 18601 23743 18659 23749
rect 26418 23740 26424 23792
rect 26476 23780 26482 23792
rect 29822 23780 29828 23792
rect 26476 23752 29828 23780
rect 26476 23740 26482 23752
rect 29822 23740 29828 23752
rect 29880 23740 29886 23792
rect 30834 23740 30840 23792
rect 30892 23780 30898 23792
rect 34514 23780 34520 23792
rect 30892 23752 34520 23780
rect 30892 23740 30898 23752
rect 7190 23712 7196 23724
rect 6411 23684 6914 23712
rect 7151 23684 7196 23712
rect 6411 23681 6423 23684
rect 6365 23675 6423 23681
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 14093 23715 14151 23721
rect 14093 23681 14105 23715
rect 14139 23712 14151 23715
rect 14182 23712 14188 23724
rect 14139 23684 14188 23712
rect 14139 23681 14151 23684
rect 14093 23675 14151 23681
rect 14182 23672 14188 23684
rect 14240 23712 14246 23724
rect 15105 23715 15163 23721
rect 15105 23712 15117 23715
rect 14240 23684 15117 23712
rect 14240 23672 14246 23684
rect 15105 23681 15117 23684
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 20438 23672 20444 23724
rect 20496 23712 20502 23724
rect 20496 23684 20541 23712
rect 20496 23672 20502 23684
rect 22094 23672 22100 23724
rect 22152 23712 22158 23724
rect 22281 23715 22339 23721
rect 22281 23712 22293 23715
rect 22152 23684 22293 23712
rect 22152 23672 22158 23684
rect 22281 23681 22293 23684
rect 22327 23681 22339 23715
rect 27154 23712 27160 23724
rect 27115 23684 27160 23712
rect 22281 23675 22339 23681
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 32232 23721 32260 23752
rect 34514 23740 34520 23752
rect 34572 23780 34578 23792
rect 34572 23752 35388 23780
rect 34572 23740 34578 23752
rect 32490 23721 32496 23724
rect 32217 23715 32275 23721
rect 32217 23681 32229 23715
rect 32263 23681 32275 23715
rect 32484 23712 32496 23721
rect 32451 23684 32496 23712
rect 32217 23675 32275 23681
rect 32484 23675 32496 23684
rect 32490 23672 32496 23675
rect 32548 23672 32554 23724
rect 34701 23715 34759 23721
rect 34701 23681 34713 23715
rect 34747 23681 34759 23715
rect 34882 23712 34888 23724
rect 34843 23684 34888 23712
rect 34701 23675 34759 23681
rect 7374 23644 7380 23656
rect 7335 23616 7380 23644
rect 7374 23604 7380 23616
rect 7432 23604 7438 23656
rect 9033 23647 9091 23653
rect 9033 23613 9045 23647
rect 9079 23613 9091 23647
rect 11606 23644 11612 23656
rect 11567 23616 11612 23644
rect 9033 23607 9091 23613
rect 3418 23536 3424 23588
rect 3476 23576 3482 23588
rect 9048 23576 9076 23607
rect 11606 23604 11612 23616
rect 11664 23604 11670 23656
rect 13449 23647 13507 23653
rect 13449 23613 13461 23647
rect 13495 23644 13507 23647
rect 13538 23644 13544 23656
rect 13495 23616 13544 23644
rect 13495 23613 13507 23616
rect 13449 23607 13507 23613
rect 13464 23576 13492 23607
rect 13538 23604 13544 23616
rect 13596 23604 13602 23656
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23644 14335 23647
rect 14458 23644 14464 23656
rect 14323 23616 14464 23644
rect 14323 23613 14335 23616
rect 14277 23607 14335 23613
rect 14458 23604 14464 23616
rect 14516 23644 14522 23656
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 14516 23616 15025 23644
rect 14516 23604 14522 23616
rect 15013 23613 15025 23616
rect 15059 23644 15071 23647
rect 15286 23644 15292 23656
rect 15059 23616 15292 23644
rect 15059 23613 15071 23616
rect 15013 23607 15071 23613
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 19484 23616 20269 23644
rect 19484 23604 19490 23616
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 20257 23607 20315 23613
rect 29086 23604 29092 23656
rect 29144 23644 29150 23656
rect 29641 23647 29699 23653
rect 29641 23644 29653 23647
rect 29144 23616 29653 23644
rect 29144 23604 29150 23616
rect 29641 23613 29653 23616
rect 29687 23644 29699 23647
rect 29730 23644 29736 23656
rect 29687 23616 29736 23644
rect 29687 23613 29699 23616
rect 29641 23607 29699 23613
rect 29730 23604 29736 23616
rect 29788 23604 29794 23656
rect 34241 23647 34299 23653
rect 34241 23613 34253 23647
rect 34287 23644 34299 23647
rect 34716 23644 34744 23675
rect 34882 23672 34888 23684
rect 34940 23672 34946 23724
rect 35360 23721 35388 23752
rect 35526 23740 35532 23792
rect 35584 23789 35590 23792
rect 35584 23783 35648 23789
rect 35584 23749 35602 23783
rect 35636 23749 35648 23783
rect 35584 23743 35648 23749
rect 35584 23740 35590 23743
rect 35345 23715 35403 23721
rect 35345 23681 35357 23715
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 37277 23715 37335 23721
rect 37277 23681 37289 23715
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 34790 23644 34796 23656
rect 34287 23616 34796 23644
rect 34287 23613 34299 23616
rect 34241 23607 34299 23613
rect 34790 23604 34796 23616
rect 34848 23604 34854 23656
rect 3476 23548 13492 23576
rect 22465 23579 22523 23585
rect 3476 23536 3482 23548
rect 22465 23545 22477 23579
rect 22511 23576 22523 23579
rect 23474 23576 23480 23588
rect 22511 23548 23480 23576
rect 22511 23545 22523 23548
rect 22465 23539 22523 23545
rect 23474 23536 23480 23548
rect 23532 23536 23538 23588
rect 36722 23576 36728 23588
rect 36635 23548 36728 23576
rect 36722 23536 36728 23548
rect 36780 23576 36786 23588
rect 37292 23576 37320 23675
rect 36780 23548 37320 23576
rect 36780 23536 36786 23548
rect 6546 23508 6552 23520
rect 6507 23480 6552 23508
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14093 23511 14151 23517
rect 14093 23508 14105 23511
rect 13872 23480 14105 23508
rect 13872 23468 13878 23480
rect 14093 23477 14105 23480
rect 14139 23508 14151 23511
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 14139 23480 14841 23508
rect 14139 23477 14151 23480
rect 14093 23471 14151 23477
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 14829 23471 14887 23477
rect 15289 23511 15347 23517
rect 15289 23477 15301 23511
rect 15335 23508 15347 23511
rect 16022 23508 16028 23520
rect 15335 23480 16028 23508
rect 15335 23477 15347 23480
rect 15289 23471 15347 23477
rect 16022 23468 16028 23480
rect 16080 23468 16086 23520
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 16945 23511 17003 23517
rect 16945 23508 16957 23511
rect 16908 23480 16957 23508
rect 16908 23468 16914 23480
rect 16945 23477 16957 23480
rect 16991 23477 17003 23511
rect 22922 23508 22928 23520
rect 22883 23480 22928 23508
rect 16945 23471 17003 23477
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 26786 23468 26792 23520
rect 26844 23508 26850 23520
rect 26973 23511 27031 23517
rect 26973 23508 26985 23511
rect 26844 23480 26985 23508
rect 26844 23468 26850 23480
rect 26973 23477 26985 23480
rect 27019 23477 27031 23511
rect 26973 23471 27031 23477
rect 33597 23511 33655 23517
rect 33597 23477 33609 23511
rect 33643 23508 33655 23511
rect 33870 23508 33876 23520
rect 33643 23480 33876 23508
rect 33643 23477 33655 23480
rect 33597 23471 33655 23477
rect 33870 23468 33876 23480
rect 33928 23468 33934 23520
rect 34885 23511 34943 23517
rect 34885 23477 34897 23511
rect 34931 23508 34943 23511
rect 35618 23508 35624 23520
rect 34931 23480 35624 23508
rect 34931 23477 34943 23480
rect 34885 23471 34943 23477
rect 35618 23468 35624 23480
rect 35676 23468 35682 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 6546 23304 6552 23316
rect 6507 23276 6552 23304
rect 6546 23264 6552 23276
rect 6604 23264 6610 23316
rect 7374 23264 7380 23316
rect 7432 23304 7438 23316
rect 7929 23307 7987 23313
rect 7929 23304 7941 23307
rect 7432 23276 7941 23304
rect 7432 23264 7438 23276
rect 7929 23273 7941 23276
rect 7975 23273 7987 23307
rect 7929 23267 7987 23273
rect 11606 23264 11612 23316
rect 11664 23304 11670 23316
rect 11701 23307 11759 23313
rect 11701 23304 11713 23307
rect 11664 23276 11713 23304
rect 11664 23264 11670 23276
rect 11701 23273 11713 23276
rect 11747 23273 11759 23307
rect 11701 23267 11759 23273
rect 13173 23307 13231 23313
rect 13173 23273 13185 23307
rect 13219 23304 13231 23307
rect 13814 23304 13820 23316
rect 13219 23276 13820 23304
rect 13219 23273 13231 23276
rect 13173 23267 13231 23273
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 14090 23304 14096 23316
rect 14051 23276 14096 23304
rect 14090 23264 14096 23276
rect 14148 23264 14154 23316
rect 14277 23307 14335 23313
rect 14277 23273 14289 23307
rect 14323 23273 14335 23307
rect 14277 23267 14335 23273
rect 5629 23239 5687 23245
rect 5629 23205 5641 23239
rect 5675 23236 5687 23239
rect 6638 23236 6644 23248
rect 5675 23208 6644 23236
rect 5675 23205 5687 23208
rect 5629 23199 5687 23205
rect 6380 23177 6408 23208
rect 6638 23196 6644 23208
rect 6696 23196 6702 23248
rect 6730 23196 6736 23248
rect 6788 23236 6794 23248
rect 7834 23236 7840 23248
rect 6788 23208 7840 23236
rect 6788 23196 6794 23208
rect 7834 23196 7840 23208
rect 7892 23196 7898 23248
rect 13832 23236 13860 23264
rect 14292 23236 14320 23267
rect 27154 23264 27160 23316
rect 27212 23304 27218 23316
rect 27525 23307 27583 23313
rect 27525 23304 27537 23307
rect 27212 23276 27537 23304
rect 27212 23264 27218 23276
rect 27525 23273 27537 23276
rect 27571 23273 27583 23307
rect 27525 23267 27583 23273
rect 36814 23264 36820 23316
rect 36872 23304 36878 23316
rect 36909 23307 36967 23313
rect 36909 23304 36921 23307
rect 36872 23276 36921 23304
rect 36872 23264 36878 23276
rect 36909 23273 36921 23276
rect 36955 23273 36967 23307
rect 36909 23267 36967 23273
rect 15013 23239 15071 23245
rect 15013 23236 15025 23239
rect 13832 23208 15025 23236
rect 15013 23205 15025 23208
rect 15059 23205 15071 23239
rect 15013 23199 15071 23205
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23137 6423 23171
rect 7742 23168 7748 23180
rect 6365 23131 6423 23137
rect 6472 23140 7748 23168
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23100 1458 23112
rect 2041 23103 2099 23109
rect 2041 23100 2053 23103
rect 1452 23072 2053 23100
rect 1452 23060 1458 23072
rect 2041 23069 2053 23072
rect 2087 23069 2099 23103
rect 2041 23063 2099 23069
rect 2774 23060 2780 23112
rect 2832 23100 2838 23112
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2832 23072 2881 23100
rect 2832 23060 2838 23072
rect 2869 23069 2881 23072
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23100 4031 23103
rect 5350 23100 5356 23112
rect 4019 23072 5356 23100
rect 4019 23069 4031 23072
rect 3973 23063 4031 23069
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23069 5871 23103
rect 5813 23063 5871 23069
rect 6273 23103 6331 23109
rect 6273 23069 6285 23103
rect 6319 23100 6331 23103
rect 6472 23100 6500 23140
rect 7742 23128 7748 23140
rect 7800 23128 7806 23180
rect 14458 23168 14464 23180
rect 14419 23140 14464 23168
rect 14458 23128 14464 23140
rect 14516 23128 14522 23180
rect 16850 23168 16856 23180
rect 16811 23140 16856 23168
rect 16850 23128 16856 23140
rect 16908 23128 16914 23180
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 22922 23168 22928 23180
rect 22051 23140 22928 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 22922 23128 22928 23140
rect 22980 23128 22986 23180
rect 23845 23171 23903 23177
rect 23845 23137 23857 23171
rect 23891 23168 23903 23171
rect 23934 23168 23940 23180
rect 23891 23140 23940 23168
rect 23891 23137 23903 23140
rect 23845 23131 23903 23137
rect 23934 23128 23940 23140
rect 23992 23128 23998 23180
rect 6319 23072 6500 23100
rect 6549 23103 6607 23109
rect 6319 23069 6331 23072
rect 6273 23063 6331 23069
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 2958 22924 2964 22976
rect 3016 22964 3022 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 3016 22936 3801 22964
rect 3016 22924 3022 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 5169 22967 5227 22973
rect 5169 22933 5181 22967
rect 5215 22964 5227 22967
rect 5626 22964 5632 22976
rect 5215 22936 5632 22964
rect 5215 22933 5227 22936
rect 5169 22927 5227 22933
rect 5626 22924 5632 22936
rect 5684 22964 5690 22976
rect 5828 22964 5856 23063
rect 6380 23044 6408 23072
rect 6549 23069 6561 23103
rect 6595 23069 6607 23103
rect 6549 23063 6607 23069
rect 6362 22992 6368 23044
rect 6420 22992 6426 23044
rect 6454 22992 6460 23044
rect 6512 23032 6518 23044
rect 6564 23032 6592 23063
rect 6730 23060 6736 23112
rect 6788 23060 6794 23112
rect 6822 23060 6828 23112
rect 6880 23100 6886 23112
rect 7285 23103 7343 23109
rect 7285 23100 7297 23103
rect 6880 23072 7297 23100
rect 6880 23060 6886 23072
rect 7285 23069 7297 23072
rect 7331 23069 7343 23103
rect 8113 23103 8171 23109
rect 8113 23100 8125 23103
rect 7285 23063 7343 23069
rect 7392 23072 8125 23100
rect 6748 23032 6776 23060
rect 6512 23004 6592 23032
rect 6656 23004 6776 23032
rect 6512 22992 6518 23004
rect 6656 22964 6684 23004
rect 5684 22936 6684 22964
rect 6733 22967 6791 22973
rect 5684 22924 5690 22936
rect 6733 22933 6745 22967
rect 6779 22964 6791 22967
rect 7392 22964 7420 23072
rect 8113 23069 8125 23072
rect 8159 23069 8171 23103
rect 8113 23063 8171 23069
rect 8941 23103 8999 23109
rect 8941 23069 8953 23103
rect 8987 23069 8999 23103
rect 12894 23100 12900 23112
rect 12855 23072 12900 23100
rect 8941 23063 8999 23069
rect 7650 22992 7656 23044
rect 7708 23032 7714 23044
rect 8956 23032 8984 23063
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 12986 23060 12992 23112
rect 13044 23100 13050 23112
rect 13170 23100 13176 23112
rect 13044 23072 13089 23100
rect 13131 23072 13176 23100
rect 13044 23060 13050 23072
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 14277 23103 14335 23109
rect 14277 23100 14289 23103
rect 14240 23072 14289 23100
rect 14240 23060 14246 23072
rect 14277 23069 14289 23072
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 14553 23103 14611 23109
rect 14553 23069 14565 23103
rect 14599 23100 14611 23103
rect 14826 23100 14832 23112
rect 14599 23072 14832 23100
rect 14599 23069 14611 23072
rect 14553 23063 14611 23069
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 15197 23103 15255 23109
rect 15197 23069 15209 23103
rect 15243 23100 15255 23103
rect 15654 23100 15660 23112
rect 15243 23072 15660 23100
rect 15243 23069 15255 23072
rect 15197 23063 15255 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 16022 23100 16028 23112
rect 15983 23072 16028 23100
rect 16022 23060 16028 23072
rect 16080 23060 16086 23112
rect 26786 23060 26792 23112
rect 26844 23109 26850 23112
rect 26844 23100 26856 23109
rect 27062 23100 27068 23112
rect 26844 23072 26889 23100
rect 27023 23072 27068 23100
rect 26844 23063 26856 23072
rect 26844 23060 26850 23063
rect 27062 23060 27068 23072
rect 27120 23060 27126 23112
rect 27522 23060 27528 23112
rect 27580 23100 27586 23112
rect 27709 23103 27767 23109
rect 27709 23100 27721 23103
rect 27580 23072 27721 23100
rect 27580 23060 27586 23072
rect 27709 23069 27721 23072
rect 27755 23069 27767 23103
rect 27890 23100 27896 23112
rect 27851 23072 27896 23100
rect 27709 23063 27767 23069
rect 27890 23060 27896 23072
rect 27948 23060 27954 23112
rect 34514 23060 34520 23112
rect 34572 23100 34578 23112
rect 35529 23103 35587 23109
rect 35529 23100 35541 23103
rect 34572 23072 35541 23100
rect 34572 23060 34578 23072
rect 35529 23069 35541 23072
rect 35575 23069 35587 23103
rect 35529 23063 35587 23069
rect 35618 23060 35624 23112
rect 35676 23100 35682 23112
rect 35785 23103 35843 23109
rect 35785 23100 35797 23103
rect 35676 23072 35797 23100
rect 35676 23060 35682 23072
rect 35785 23069 35797 23072
rect 35831 23069 35843 23103
rect 35785 23063 35843 23069
rect 17037 23035 17095 23041
rect 17037 23032 17049 23035
rect 7708 23004 8984 23032
rect 16546 23004 17049 23032
rect 7708 22992 7714 23004
rect 6779 22936 7420 22964
rect 7469 22967 7527 22973
rect 6779 22933 6791 22936
rect 6733 22927 6791 22933
rect 7469 22933 7481 22967
rect 7515 22964 7527 22967
rect 7834 22964 7840 22976
rect 7515 22936 7840 22964
rect 7515 22933 7527 22936
rect 7469 22927 7527 22933
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 12710 22964 12716 22976
rect 12671 22936 12716 22964
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 16209 22967 16267 22973
rect 16209 22933 16221 22967
rect 16255 22964 16267 22967
rect 16546 22964 16574 23004
rect 17037 23001 17049 23004
rect 17083 23001 17095 23035
rect 17037 22995 17095 23001
rect 18693 23035 18751 23041
rect 18693 23001 18705 23035
rect 18739 23032 18751 23035
rect 19334 23032 19340 23044
rect 18739 23004 19340 23032
rect 18739 23001 18751 23004
rect 18693 22995 18751 23001
rect 19334 22992 19340 23004
rect 19392 22992 19398 23044
rect 22189 23035 22247 23041
rect 22189 23001 22201 23035
rect 22235 23032 22247 23035
rect 22738 23032 22744 23044
rect 22235 23004 22744 23032
rect 22235 23001 22247 23004
rect 22189 22995 22247 23001
rect 22738 22992 22744 23004
rect 22796 22992 22802 23044
rect 25682 22964 25688 22976
rect 16255 22936 16574 22964
rect 25643 22936 25688 22964
rect 16255 22933 16267 22936
rect 16209 22927 16267 22933
rect 25682 22924 25688 22936
rect 25740 22924 25746 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 5350 22760 5356 22772
rect 5311 22732 5356 22760
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 6822 22760 6828 22772
rect 5736 22732 6684 22760
rect 6783 22732 6828 22760
rect 2958 22692 2964 22704
rect 2919 22664 2964 22692
rect 2958 22652 2964 22664
rect 3016 22652 3022 22704
rect 3602 22652 3608 22704
rect 3660 22692 3666 22704
rect 5736 22692 5764 22732
rect 3660 22664 5764 22692
rect 5813 22695 5871 22701
rect 3660 22652 3666 22664
rect 5813 22661 5825 22695
rect 5859 22692 5871 22695
rect 6362 22692 6368 22704
rect 5859 22664 6368 22692
rect 5859 22661 5871 22664
rect 5813 22655 5871 22661
rect 6362 22652 6368 22664
rect 6420 22652 6426 22704
rect 6656 22692 6684 22732
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 7668 22732 9536 22760
rect 7668 22692 7696 22732
rect 7834 22692 7840 22704
rect 6656 22664 7696 22692
rect 7795 22664 7840 22692
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 9508 22701 9536 22732
rect 12894 22720 12900 22772
rect 12952 22760 12958 22772
rect 14182 22760 14188 22772
rect 12952 22732 14188 22760
rect 12952 22720 12958 22732
rect 14182 22720 14188 22732
rect 14240 22760 14246 22772
rect 14553 22763 14611 22769
rect 14553 22760 14565 22763
rect 14240 22732 14565 22760
rect 14240 22720 14246 22732
rect 14553 22729 14565 22732
rect 14599 22729 14611 22763
rect 27522 22760 27528 22772
rect 27483 22732 27528 22760
rect 14553 22723 14611 22729
rect 27522 22720 27528 22732
rect 27580 22720 27586 22772
rect 27890 22720 27896 22772
rect 27948 22760 27954 22772
rect 30469 22763 30527 22769
rect 30469 22760 30481 22763
rect 27948 22732 30481 22760
rect 27948 22720 27954 22732
rect 30469 22729 30481 22732
rect 30515 22760 30527 22763
rect 32030 22760 32036 22772
rect 30515 22732 32036 22760
rect 30515 22729 30527 22732
rect 30469 22723 30527 22729
rect 32030 22720 32036 22732
rect 32088 22720 32094 22772
rect 35894 22720 35900 22772
rect 35952 22760 35958 22772
rect 36173 22763 36231 22769
rect 36173 22760 36185 22763
rect 35952 22732 36185 22760
rect 35952 22720 35958 22732
rect 36173 22729 36185 22732
rect 36219 22729 36231 22763
rect 36173 22723 36231 22729
rect 9493 22695 9551 22701
rect 9493 22661 9505 22695
rect 9539 22692 9551 22695
rect 19981 22695 20039 22701
rect 9539 22664 13308 22692
rect 9539 22661 9551 22664
rect 9493 22655 9551 22661
rect 2774 22624 2780 22636
rect 2735 22596 2780 22624
rect 2774 22584 2780 22596
rect 2832 22584 2838 22636
rect 4614 22624 4620 22636
rect 4575 22596 4620 22624
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22624 5595 22627
rect 6454 22624 6460 22636
rect 5583 22596 6460 22624
rect 5583 22593 5595 22596
rect 5537 22587 5595 22593
rect 6454 22584 6460 22596
rect 6512 22624 6518 22636
rect 6641 22627 6699 22633
rect 6641 22624 6653 22627
rect 6512 22596 6653 22624
rect 6512 22584 6518 22596
rect 6641 22593 6653 22596
rect 6687 22593 6699 22627
rect 7650 22624 7656 22636
rect 7611 22596 7656 22624
rect 6641 22587 6699 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 4632 22488 4660 22584
rect 13280 22568 13308 22664
rect 19981 22661 19993 22695
rect 20027 22692 20039 22695
rect 23842 22692 23848 22704
rect 20027 22664 23848 22692
rect 20027 22661 20039 22664
rect 19981 22655 20039 22661
rect 23842 22652 23848 22664
rect 23900 22652 23906 22704
rect 25682 22652 25688 22704
rect 25740 22692 25746 22704
rect 27249 22695 27307 22701
rect 27249 22692 27261 22695
rect 25740 22664 27261 22692
rect 25740 22652 25746 22664
rect 27249 22661 27261 22664
rect 27295 22661 27307 22695
rect 27249 22655 27307 22661
rect 34057 22695 34115 22701
rect 34057 22661 34069 22695
rect 34103 22692 34115 22695
rect 34698 22692 34704 22704
rect 34103 22664 34704 22692
rect 34103 22661 34115 22664
rect 34057 22655 34115 22661
rect 34698 22652 34704 22664
rect 34756 22652 34762 22704
rect 14734 22624 14740 22636
rect 14695 22596 14740 22624
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 24673 22627 24731 22633
rect 24673 22593 24685 22627
rect 24719 22624 24731 22627
rect 25700 22624 25728 22652
rect 26878 22624 26884 22636
rect 24719 22596 25728 22624
rect 26344 22596 26884 22624
rect 24719 22593 24731 22596
rect 24673 22587 24731 22593
rect 5721 22559 5779 22565
rect 5721 22525 5733 22559
rect 5767 22556 5779 22559
rect 6549 22559 6607 22565
rect 6549 22556 6561 22559
rect 5767 22528 6561 22556
rect 5767 22525 5779 22528
rect 5721 22519 5779 22525
rect 6549 22525 6561 22528
rect 6595 22556 6607 22559
rect 6730 22556 6736 22568
rect 6595 22528 6736 22556
rect 6595 22525 6607 22528
rect 6549 22519 6607 22525
rect 6730 22516 6736 22528
rect 6788 22516 6794 22568
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22556 11023 22559
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11011 22528 11529 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11698 22556 11704 22568
rect 11659 22528 11704 22556
rect 11517 22519 11575 22525
rect 11698 22516 11704 22528
rect 11756 22516 11762 22568
rect 13262 22556 13268 22568
rect 13223 22528 13268 22556
rect 13262 22516 13268 22528
rect 13320 22516 13326 22568
rect 18138 22556 18144 22568
rect 18099 22528 18144 22556
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 18322 22556 18328 22568
rect 18283 22528 18328 22556
rect 18322 22516 18328 22528
rect 18380 22516 18386 22568
rect 24213 22559 24271 22565
rect 24213 22525 24225 22559
rect 24259 22525 24271 22559
rect 24486 22556 24492 22568
rect 24447 22528 24492 22556
rect 24213 22519 24271 22525
rect 19334 22488 19340 22500
rect 4632 22460 19340 22488
rect 19334 22448 19340 22460
rect 19392 22448 19398 22500
rect 24228 22488 24256 22519
rect 24486 22516 24492 22528
rect 24544 22516 24550 22568
rect 26344 22500 26372 22596
rect 26878 22584 26884 22596
rect 26936 22624 26942 22636
rect 26973 22627 27031 22633
rect 26973 22624 26985 22627
rect 26936 22596 26985 22624
rect 26936 22584 26942 22596
rect 26973 22593 26985 22596
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22624 27399 22627
rect 29454 22624 29460 22636
rect 27387 22596 29460 22624
rect 27387 22593 27399 22596
rect 27341 22587 27399 22593
rect 27172 22556 27200 22587
rect 29454 22584 29460 22596
rect 29512 22584 29518 22636
rect 30006 22584 30012 22636
rect 30064 22624 30070 22636
rect 30561 22627 30619 22633
rect 30561 22624 30573 22627
rect 30064 22596 30573 22624
rect 30064 22584 30070 22596
rect 30561 22593 30573 22596
rect 30607 22593 30619 22627
rect 33870 22624 33876 22636
rect 33831 22596 33876 22624
rect 30561 22587 30619 22593
rect 33870 22584 33876 22596
rect 33928 22584 33934 22636
rect 35621 22627 35679 22633
rect 35621 22593 35633 22627
rect 35667 22624 35679 22627
rect 36265 22627 36323 22633
rect 36265 22624 36277 22627
rect 35667 22596 36277 22624
rect 35667 22593 35679 22596
rect 35621 22587 35679 22593
rect 36265 22593 36277 22596
rect 36311 22624 36323 22627
rect 37182 22624 37188 22636
rect 36311 22596 37188 22624
rect 36311 22593 36323 22596
rect 36265 22587 36323 22593
rect 37182 22584 37188 22596
rect 37240 22584 37246 22636
rect 28166 22556 28172 22568
rect 27172 22528 28172 22556
rect 28166 22516 28172 22528
rect 28224 22516 28230 22568
rect 26326 22488 26332 22500
rect 24228 22460 26332 22488
rect 26326 22448 26332 22460
rect 26384 22448 26390 22500
rect 5813 22423 5871 22429
rect 5813 22389 5825 22423
rect 5859 22420 5871 22423
rect 6546 22420 6552 22432
rect 5859 22392 6552 22420
rect 5859 22389 5871 22392
rect 5813 22383 5871 22389
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 6457 22219 6515 22225
rect 6457 22185 6469 22219
rect 6503 22216 6515 22219
rect 6546 22216 6552 22228
rect 6503 22188 6552 22216
rect 6503 22185 6515 22188
rect 6457 22179 6515 22185
rect 6546 22176 6552 22188
rect 6604 22176 6610 22228
rect 13173 22219 13231 22225
rect 13173 22185 13185 22219
rect 13219 22216 13231 22219
rect 13814 22216 13820 22228
rect 13219 22188 13820 22216
rect 13219 22185 13231 22188
rect 13173 22179 13231 22185
rect 13814 22176 13820 22188
rect 13872 22176 13878 22228
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18233 22219 18291 22225
rect 18233 22216 18245 22219
rect 18196 22188 18245 22216
rect 18196 22176 18202 22188
rect 18233 22185 18245 22188
rect 18279 22185 18291 22219
rect 18233 22179 18291 22185
rect 36170 22108 36176 22160
rect 36228 22148 36234 22160
rect 36228 22120 36308 22148
rect 36228 22108 36234 22120
rect 36280 22094 36308 22120
rect 6365 22083 6423 22089
rect 6365 22049 6377 22083
rect 6411 22080 6423 22083
rect 6638 22080 6644 22092
rect 6411 22052 6644 22080
rect 6411 22049 6423 22052
rect 6365 22043 6423 22049
rect 6638 22040 6644 22052
rect 6696 22040 6702 22092
rect 12986 22080 12992 22092
rect 12947 22052 12992 22080
rect 12986 22040 12992 22052
rect 13044 22040 13050 22092
rect 20809 22083 20867 22089
rect 20809 22049 20821 22083
rect 20855 22080 20867 22083
rect 20990 22080 20996 22092
rect 20855 22052 20996 22080
rect 20855 22049 20867 22052
rect 20809 22043 20867 22049
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 22738 22080 22744 22092
rect 22699 22052 22744 22080
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 25682 22080 25688 22092
rect 25643 22052 25688 22080
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 26418 22080 26424 22092
rect 26379 22052 26424 22080
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 29454 22040 29460 22092
rect 29512 22080 29518 22092
rect 36280 22089 36345 22094
rect 29917 22083 29975 22089
rect 29917 22080 29929 22083
rect 29512 22052 29929 22080
rect 29512 22040 29518 22052
rect 29917 22049 29929 22052
rect 29963 22049 29975 22083
rect 29917 22043 29975 22049
rect 36265 22083 36345 22089
rect 36265 22049 36277 22083
rect 36311 22066 36345 22083
rect 36311 22049 36323 22066
rect 36265 22043 36323 22049
rect 6454 22012 6460 22024
rect 6415 21984 6460 22012
rect 6454 21972 6460 21984
rect 6512 22012 6518 22024
rect 7282 22012 7288 22024
rect 6512 21984 7144 22012
rect 7243 21984 7288 22012
rect 6512 21972 6518 21984
rect 6181 21947 6239 21953
rect 6181 21913 6193 21947
rect 6227 21944 6239 21947
rect 6914 21944 6920 21956
rect 6227 21916 6920 21944
rect 6227 21913 6239 21916
rect 6181 21907 6239 21913
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 6641 21879 6699 21885
rect 6641 21845 6653 21879
rect 6687 21876 6699 21879
rect 7006 21876 7012 21888
rect 6687 21848 7012 21876
rect 6687 21845 6699 21848
rect 6641 21839 6699 21845
rect 7006 21836 7012 21848
rect 7064 21836 7070 21888
rect 7116 21885 7144 21984
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 10318 21972 10324 22024
rect 10376 22012 10382 22024
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 10376 21984 10425 22012
rect 10376 21972 10382 21984
rect 10413 21981 10425 21984
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 11701 22015 11759 22021
rect 11701 21981 11713 22015
rect 11747 22012 11759 22015
rect 12894 22012 12900 22024
rect 11747 21984 12434 22012
rect 12855 21984 12900 22012
rect 11747 21981 11759 21984
rect 11701 21975 11759 21981
rect 7101 21879 7159 21885
rect 7101 21845 7113 21879
rect 7147 21845 7159 21879
rect 7101 21839 7159 21845
rect 10502 21836 10508 21888
rect 10560 21876 10566 21888
rect 11517 21879 11575 21885
rect 11517 21876 11529 21879
rect 10560 21848 11529 21876
rect 10560 21836 10566 21848
rect 11517 21845 11529 21848
rect 11563 21845 11575 21879
rect 12406 21876 12434 21984
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 13170 22012 13176 22024
rect 13131 21984 13176 22012
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 19242 22012 19248 22024
rect 19203 21984 19248 22012
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 22462 22012 22468 22024
rect 22423 21984 22468 22012
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 27706 22012 27712 22024
rect 27667 21984 27712 22012
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 30374 21972 30380 22024
rect 30432 22012 30438 22024
rect 31941 22015 31999 22021
rect 31941 22012 31953 22015
rect 30432 21984 31953 22012
rect 30432 21972 30438 21984
rect 31941 21981 31953 21984
rect 31987 21981 31999 22015
rect 31941 21975 31999 21981
rect 36173 22015 36231 22021
rect 36173 21981 36185 22015
rect 36219 22012 36231 22015
rect 36354 22012 36360 22024
rect 36219 21984 36360 22012
rect 36219 21981 36231 21984
rect 36173 21975 36231 21981
rect 36354 21972 36360 21984
rect 36412 22012 36418 22024
rect 36814 22012 36820 22024
rect 36412 21984 36820 22012
rect 36412 21972 36418 21984
rect 36814 21972 36820 21984
rect 36872 21972 36878 22024
rect 37829 22015 37887 22021
rect 37829 22012 37841 22015
rect 37384 21984 37841 22012
rect 19978 21904 19984 21956
rect 20036 21944 20042 21956
rect 20625 21947 20683 21953
rect 20625 21944 20637 21947
rect 20036 21916 20637 21944
rect 20036 21904 20042 21916
rect 20625 21913 20637 21916
rect 20671 21913 20683 21947
rect 26234 21944 26240 21956
rect 26195 21916 26240 21944
rect 20625 21907 20683 21913
rect 26234 21904 26240 21916
rect 26292 21904 26298 21956
rect 28994 21944 29000 21956
rect 27356 21916 29000 21944
rect 12713 21879 12771 21885
rect 12713 21876 12725 21879
rect 12406 21848 12725 21876
rect 11517 21839 11575 21845
rect 12713 21845 12725 21848
rect 12759 21845 12771 21879
rect 19426 21876 19432 21888
rect 19387 21848 19432 21876
rect 12713 21839 12771 21845
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 25682 21836 25688 21888
rect 25740 21876 25746 21888
rect 27356 21876 27384 21916
rect 28994 21904 29000 21916
rect 29052 21904 29058 21956
rect 30098 21944 30104 21956
rect 30059 21916 30104 21944
rect 30098 21904 30104 21916
rect 30156 21904 30162 21956
rect 36081 21947 36139 21953
rect 36081 21913 36093 21947
rect 36127 21944 36139 21947
rect 36262 21944 36268 21956
rect 36127 21916 36268 21944
rect 36127 21913 36139 21916
rect 36081 21907 36139 21913
rect 36262 21904 36268 21916
rect 36320 21944 36326 21956
rect 36722 21944 36728 21956
rect 36320 21916 36728 21944
rect 36320 21904 36326 21916
rect 36722 21904 36728 21916
rect 36780 21904 36786 21956
rect 37384 21888 37412 21984
rect 37829 21981 37841 21984
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 27522 21876 27528 21888
rect 25740 21848 27384 21876
rect 27483 21848 27528 21876
rect 25740 21836 25746 21848
rect 27522 21836 27528 21848
rect 27580 21836 27586 21888
rect 32030 21876 32036 21888
rect 31991 21848 32036 21876
rect 32030 21836 32036 21848
rect 32088 21836 32094 21888
rect 35710 21876 35716 21888
rect 35671 21848 35716 21876
rect 35710 21836 35716 21848
rect 35768 21836 35774 21888
rect 37366 21876 37372 21888
rect 37327 21848 37372 21876
rect 37366 21836 37372 21848
rect 37424 21836 37430 21888
rect 38010 21876 38016 21888
rect 37971 21848 38016 21876
rect 38010 21836 38016 21848
rect 38068 21836 38074 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 11698 21632 11704 21684
rect 11756 21672 11762 21684
rect 11885 21675 11943 21681
rect 11885 21672 11897 21675
rect 11756 21644 11897 21672
rect 11756 21632 11762 21644
rect 11885 21641 11897 21644
rect 11931 21641 11943 21675
rect 11885 21635 11943 21641
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 13354 21672 13360 21684
rect 13228 21644 13360 21672
rect 13228 21632 13234 21644
rect 13354 21632 13360 21644
rect 13412 21672 13418 21684
rect 13541 21675 13599 21681
rect 13541 21672 13553 21675
rect 13412 21644 13553 21672
rect 13412 21632 13418 21644
rect 13541 21641 13553 21644
rect 13587 21641 13599 21675
rect 17126 21672 17132 21684
rect 17087 21644 17132 21672
rect 13541 21635 13599 21641
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 27706 21632 27712 21684
rect 27764 21672 27770 21684
rect 28813 21675 28871 21681
rect 28813 21672 28825 21675
rect 27764 21644 28825 21672
rect 27764 21632 27770 21644
rect 28813 21641 28825 21644
rect 28859 21641 28871 21675
rect 28813 21635 28871 21641
rect 36265 21675 36323 21681
rect 36265 21641 36277 21675
rect 36311 21672 36323 21675
rect 36354 21672 36360 21684
rect 36311 21644 36360 21672
rect 36311 21641 36323 21644
rect 36265 21635 36323 21641
rect 36354 21632 36360 21644
rect 36412 21632 36418 21684
rect 6825 21607 6883 21613
rect 6825 21573 6837 21607
rect 6871 21604 6883 21607
rect 6914 21604 6920 21616
rect 6871 21576 6920 21604
rect 6871 21573 6883 21576
rect 6825 21567 6883 21573
rect 6914 21564 6920 21576
rect 6972 21604 6978 21616
rect 7374 21604 7380 21616
rect 6972 21576 7380 21604
rect 6972 21564 6978 21576
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 27240 21607 27298 21613
rect 27240 21573 27252 21607
rect 27286 21604 27298 21607
rect 27522 21604 27528 21616
rect 27286 21576 27528 21604
rect 27286 21573 27298 21576
rect 27240 21567 27298 21573
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 36170 21564 36176 21616
rect 36228 21604 36234 21616
rect 36228 21576 36492 21604
rect 36228 21564 36234 21576
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21536 1458 21548
rect 2041 21539 2099 21545
rect 2041 21536 2053 21539
rect 1452 21508 2053 21536
rect 1452 21496 1458 21508
rect 2041 21505 2053 21508
rect 2087 21505 2099 21539
rect 2041 21499 2099 21505
rect 6454 21496 6460 21548
rect 6512 21536 6518 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6638 21496 6644 21548
rect 6696 21536 6702 21548
rect 6696 21508 6741 21536
rect 6696 21496 6702 21508
rect 7006 21496 7012 21548
rect 7064 21536 7070 21548
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 7064 21508 7481 21536
rect 7064 21496 7070 21508
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 12710 21536 12716 21548
rect 12115 21508 12716 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 13998 21536 14004 21548
rect 13771 21508 14004 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 13998 21496 14004 21508
rect 14056 21536 14062 21548
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 14056 21508 14565 21536
rect 14056 21496 14062 21508
rect 14553 21505 14565 21508
rect 14599 21536 14611 21539
rect 15194 21536 15200 21548
rect 14599 21508 15200 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 17218 21536 17224 21548
rect 17179 21508 17224 21536
rect 17218 21496 17224 21508
rect 17276 21496 17282 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20809 21539 20867 21545
rect 20809 21536 20821 21539
rect 20303 21508 20821 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20809 21505 20821 21508
rect 20855 21536 20867 21539
rect 21542 21536 21548 21548
rect 20855 21508 21548 21536
rect 20855 21505 20867 21508
rect 20809 21499 20867 21505
rect 14182 21428 14188 21480
rect 14240 21468 14246 21480
rect 14277 21471 14335 21477
rect 14277 21468 14289 21471
rect 14240 21440 14289 21468
rect 14240 21428 14246 21440
rect 14277 21437 14289 21440
rect 14323 21468 14335 21471
rect 20272 21468 20300 21499
rect 21542 21496 21548 21508
rect 21600 21496 21606 21548
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21536 22155 21539
rect 24486 21536 24492 21548
rect 22143 21508 24492 21536
rect 22143 21505 22155 21508
rect 22097 21499 22155 21505
rect 24486 21496 24492 21508
rect 24544 21496 24550 21548
rect 26973 21539 27031 21545
rect 26973 21505 26985 21539
rect 27019 21536 27031 21539
rect 27062 21536 27068 21548
rect 27019 21508 27068 21536
rect 27019 21505 27031 21508
rect 26973 21499 27031 21505
rect 27062 21496 27068 21508
rect 27120 21496 27126 21548
rect 28534 21496 28540 21548
rect 28592 21536 28598 21548
rect 28997 21539 29055 21545
rect 28997 21536 29009 21539
rect 28592 21508 29009 21536
rect 28592 21496 28598 21508
rect 28997 21505 29009 21508
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 29181 21539 29239 21545
rect 29181 21505 29193 21539
rect 29227 21536 29239 21539
rect 29914 21536 29920 21548
rect 29227 21508 29920 21536
rect 29227 21505 29239 21508
rect 29181 21499 29239 21505
rect 29914 21496 29920 21508
rect 29972 21536 29978 21548
rect 32677 21539 32735 21545
rect 29972 21508 30328 21536
rect 29972 21496 29978 21508
rect 30300 21480 30328 21508
rect 32677 21505 32689 21539
rect 32723 21536 32735 21539
rect 33870 21536 33876 21548
rect 32723 21508 33876 21536
rect 32723 21505 32735 21508
rect 32677 21499 32735 21505
rect 33870 21496 33876 21508
rect 33928 21496 33934 21548
rect 36262 21496 36268 21548
rect 36320 21536 36326 21548
rect 36357 21539 36415 21545
rect 36357 21536 36369 21539
rect 36320 21508 36369 21536
rect 36320 21496 36326 21508
rect 36357 21505 36369 21508
rect 36403 21505 36415 21539
rect 36357 21499 36415 21505
rect 14323 21440 20300 21468
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 21358 21428 21364 21480
rect 21416 21468 21422 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 21416 21440 21833 21468
rect 21416 21428 21422 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 30006 21468 30012 21480
rect 29967 21440 30012 21468
rect 21821 21431 21879 21437
rect 30006 21428 30012 21440
rect 30064 21428 30070 21480
rect 30282 21468 30288 21480
rect 30243 21440 30288 21468
rect 30282 21428 30288 21440
rect 30340 21428 30346 21480
rect 36464 21477 36492 21576
rect 36449 21471 36507 21477
rect 36449 21437 36461 21471
rect 36495 21437 36507 21471
rect 36449 21431 36507 21437
rect 5166 21360 5172 21412
rect 5224 21400 5230 21412
rect 5442 21400 5448 21412
rect 5224 21372 5448 21400
rect 5224 21360 5230 21372
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 20990 21400 20996 21412
rect 20951 21372 20996 21400
rect 20990 21360 20996 21372
rect 21048 21360 21054 21412
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 2774 21332 2780 21344
rect 1627 21304 2780 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 2774 21292 2780 21304
rect 2832 21292 2838 21344
rect 5810 21332 5816 21344
rect 5771 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 6362 21332 6368 21344
rect 6323 21304 6368 21332
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 6546 21332 6552 21344
rect 6507 21304 6552 21332
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 6730 21292 6736 21344
rect 6788 21332 6794 21344
rect 7285 21335 7343 21341
rect 7285 21332 7297 21335
rect 6788 21304 7297 21332
rect 6788 21292 6794 21304
rect 7285 21301 7297 21304
rect 7331 21301 7343 21335
rect 7285 21295 7343 21301
rect 28258 21292 28264 21344
rect 28316 21332 28322 21344
rect 28353 21335 28411 21341
rect 28353 21332 28365 21335
rect 28316 21304 28365 21332
rect 28316 21292 28322 21304
rect 28353 21301 28365 21304
rect 28399 21301 28411 21335
rect 32582 21332 32588 21344
rect 32543 21304 32588 21332
rect 28353 21295 28411 21301
rect 32582 21292 32588 21304
rect 32640 21292 32646 21344
rect 35618 21292 35624 21344
rect 35676 21332 35682 21344
rect 35897 21335 35955 21341
rect 35897 21332 35909 21335
rect 35676 21304 35909 21332
rect 35676 21292 35682 21304
rect 35897 21301 35909 21304
rect 35943 21301 35955 21335
rect 35897 21295 35955 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1578 21088 1584 21140
rect 1636 21128 1642 21140
rect 2498 21128 2504 21140
rect 1636 21100 2504 21128
rect 1636 21088 1642 21100
rect 2498 21088 2504 21100
rect 2556 21088 2562 21140
rect 14182 21128 14188 21140
rect 14143 21100 14188 21128
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 21085 21131 21143 21137
rect 21085 21097 21097 21131
rect 21131 21097 21143 21131
rect 21358 21128 21364 21140
rect 21319 21100 21364 21128
rect 21085 21091 21143 21097
rect 3418 21020 3424 21072
rect 3476 21060 3482 21072
rect 3476 21032 8432 21060
rect 3476 21020 3482 21032
rect 2774 20992 2780 21004
rect 2516 20964 2780 20992
rect 2516 20933 2544 20964
rect 2774 20952 2780 20964
rect 2832 20952 2838 21004
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 6549 20995 6607 21001
rect 6549 20992 6561 20995
rect 5868 20964 6561 20992
rect 5868 20952 5874 20964
rect 6549 20961 6561 20964
rect 6595 20961 6607 20995
rect 6730 20992 6736 21004
rect 6691 20964 6736 20992
rect 6549 20955 6607 20961
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 2501 20927 2559 20933
rect 2501 20893 2513 20927
rect 2547 20893 2559 20927
rect 2501 20887 2559 20893
rect 2590 20884 2596 20936
rect 2648 20924 2654 20936
rect 5629 20927 5687 20933
rect 2648 20896 2693 20924
rect 2648 20884 2654 20896
rect 5629 20893 5641 20927
rect 5675 20924 5687 20927
rect 6362 20924 6368 20936
rect 5675 20896 6368 20924
rect 5675 20893 5687 20896
rect 5629 20887 5687 20893
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 8404 20865 8432 21032
rect 20898 21020 20904 21072
rect 20956 21060 20962 21072
rect 21100 21060 21128 21091
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 28534 21128 28540 21140
rect 28495 21100 28540 21128
rect 28534 21088 28540 21100
rect 28592 21088 28598 21140
rect 29733 21131 29791 21137
rect 29733 21097 29745 21131
rect 29779 21128 29791 21131
rect 31478 21128 31484 21140
rect 29779 21100 31484 21128
rect 29779 21097 29791 21100
rect 29733 21091 29791 21097
rect 31478 21088 31484 21100
rect 31536 21128 31542 21140
rect 31941 21131 31999 21137
rect 31536 21100 31754 21128
rect 31536 21088 31542 21100
rect 25498 21060 25504 21072
rect 20956 21032 25504 21060
rect 20956 21020 20962 21032
rect 25498 21020 25504 21032
rect 25556 21020 25562 21072
rect 31726 21060 31754 21100
rect 31941 21097 31953 21131
rect 31987 21128 31999 21131
rect 32122 21128 32128 21140
rect 31987 21100 32128 21128
rect 31987 21097 31999 21100
rect 31941 21091 31999 21097
rect 32122 21088 32128 21100
rect 32180 21088 32186 21140
rect 32306 21060 32312 21072
rect 31726 21032 32312 21060
rect 32306 21020 32312 21032
rect 32364 21020 32370 21072
rect 10318 20992 10324 21004
rect 10279 20964 10324 20992
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 10502 20992 10508 21004
rect 10463 20964 10508 20992
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 15013 20995 15071 21001
rect 15013 20992 15025 20995
rect 14700 20964 15025 20992
rect 14700 20952 14706 20964
rect 15013 20961 15025 20964
rect 15059 20961 15071 20995
rect 15013 20955 15071 20961
rect 15194 20952 15200 21004
rect 15252 20992 15258 21004
rect 16301 20995 16359 21001
rect 16301 20992 16313 20995
rect 15252 20964 16313 20992
rect 15252 20952 15258 20964
rect 16301 20961 16313 20964
rect 16347 20961 16359 20995
rect 16574 20992 16580 21004
rect 16535 20964 16580 20992
rect 16301 20955 16359 20961
rect 16574 20952 16580 20964
rect 16632 20952 16638 21004
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20992 18199 20995
rect 18322 20992 18328 21004
rect 18187 20964 18328 20992
rect 18187 20961 18199 20964
rect 18141 20955 18199 20961
rect 18322 20952 18328 20964
rect 18380 20952 18386 21004
rect 19978 20992 19984 21004
rect 19628 20964 19984 20992
rect 14550 20884 14556 20936
rect 14608 20924 14614 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14608 20896 15301 20924
rect 14608 20884 14614 20896
rect 15289 20893 15301 20896
rect 15335 20924 15347 20927
rect 16482 20924 16488 20936
rect 15335 20896 16488 20924
rect 15335 20893 15347 20896
rect 15289 20887 15347 20893
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 18414 20924 18420 20936
rect 18375 20896 18420 20924
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19628 20933 19656 20964
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 20993 20995 21051 21001
rect 20993 20992 21005 20995
rect 20088 20964 21005 20992
rect 20088 20936 20116 20964
rect 20993 20961 21005 20964
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 24673 20995 24731 21001
rect 24673 20961 24685 20995
rect 24719 20992 24731 20995
rect 26234 20992 26240 21004
rect 24719 20964 26240 20992
rect 24719 20961 24731 20964
rect 24673 20955 24731 20961
rect 26234 20952 26240 20964
rect 26292 20952 26298 21004
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 30561 20995 30619 21001
rect 30561 20992 30573 20995
rect 27120 20964 30573 20992
rect 27120 20952 27126 20964
rect 30561 20961 30573 20964
rect 30607 20961 30619 20995
rect 30561 20955 30619 20961
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19484 20896 19625 20924
rect 19484 20884 19490 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 20070 20924 20076 20936
rect 19935 20896 20076 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 21177 20927 21235 20933
rect 21177 20924 21189 20927
rect 20772 20896 21189 20924
rect 20772 20884 20778 20896
rect 21177 20893 21189 20896
rect 21223 20893 21235 20927
rect 21818 20924 21824 20936
rect 21779 20896 21824 20924
rect 21177 20887 21235 20893
rect 8389 20859 8447 20865
rect 8389 20825 8401 20859
rect 8435 20856 8447 20859
rect 12158 20856 12164 20868
rect 8435 20828 12164 20856
rect 8435 20825 8447 20828
rect 8389 20819 8447 20825
rect 12158 20816 12164 20828
rect 12216 20816 12222 20868
rect 20438 20816 20444 20868
rect 20496 20856 20502 20868
rect 20901 20859 20959 20865
rect 20901 20856 20913 20859
rect 20496 20828 20913 20856
rect 20496 20816 20502 20828
rect 20901 20825 20913 20828
rect 20947 20825 20959 20859
rect 21192 20856 21220 20887
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 24394 20924 24400 20936
rect 24355 20896 24400 20924
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 27985 20927 28043 20933
rect 27985 20924 27997 20927
rect 27448 20896 27997 20924
rect 25774 20856 25780 20868
rect 21192 20828 25780 20856
rect 20901 20819 20959 20825
rect 25774 20816 25780 20828
rect 25832 20816 25838 20868
rect 27448 20800 27476 20896
rect 27985 20893 27997 20896
rect 28031 20893 28043 20927
rect 27985 20887 28043 20893
rect 28353 20927 28411 20933
rect 28353 20893 28365 20927
rect 28399 20924 28411 20927
rect 28399 20896 29500 20924
rect 28399 20893 28411 20896
rect 28353 20887 28411 20893
rect 28166 20856 28172 20868
rect 28079 20828 28172 20856
rect 28166 20816 28172 20828
rect 28224 20816 28230 20868
rect 28258 20816 28264 20868
rect 28316 20856 28322 20868
rect 29472 20856 29500 20896
rect 29546 20884 29552 20936
rect 29604 20924 29610 20936
rect 30576 20924 30604 20955
rect 32030 20924 32036 20936
rect 29604 20896 29649 20924
rect 30576 20896 32036 20924
rect 29604 20884 29610 20896
rect 32030 20884 32036 20896
rect 32088 20924 32094 20936
rect 34514 20924 34520 20936
rect 32088 20896 34520 20924
rect 32088 20884 32094 20896
rect 34514 20884 34520 20896
rect 34572 20884 34578 20936
rect 30098 20856 30104 20868
rect 28316 20828 28361 20856
rect 29472 20828 30104 20856
rect 28316 20816 28322 20828
rect 30098 20816 30104 20828
rect 30156 20816 30162 20868
rect 30828 20859 30886 20865
rect 30828 20825 30840 20859
rect 30874 20856 30886 20859
rect 31018 20856 31024 20868
rect 30874 20828 31024 20856
rect 30874 20825 30886 20828
rect 30828 20819 30886 20825
rect 31018 20816 31024 20828
rect 31076 20816 31082 20868
rect 1394 20788 1400 20800
rect 1355 20760 1400 20788
rect 1394 20748 1400 20760
rect 1452 20748 1458 20800
rect 2866 20788 2872 20800
rect 2827 20760 2872 20788
rect 2866 20748 2872 20760
rect 2924 20748 2930 20800
rect 4890 20748 4896 20800
rect 4948 20788 4954 20800
rect 5445 20791 5503 20797
rect 5445 20788 5457 20791
rect 4948 20760 5457 20788
rect 4948 20748 4954 20760
rect 5445 20757 5457 20760
rect 5491 20757 5503 20791
rect 5445 20751 5503 20757
rect 22005 20791 22063 20797
rect 22005 20757 22017 20791
rect 22051 20788 22063 20791
rect 23290 20788 23296 20800
rect 22051 20760 23296 20788
rect 22051 20757 22063 20760
rect 22005 20751 22063 20757
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 27430 20788 27436 20800
rect 27391 20760 27436 20788
rect 27430 20748 27436 20760
rect 27488 20748 27494 20800
rect 28184 20788 28212 20816
rect 29362 20788 29368 20800
rect 28184 20760 29368 20788
rect 29362 20748 29368 20760
rect 29420 20748 29426 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 2498 20544 2504 20596
rect 2556 20584 2562 20596
rect 17129 20587 17187 20593
rect 2556 20556 3740 20584
rect 2556 20544 2562 20556
rect 3712 20525 3740 20556
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17218 20584 17224 20596
rect 17175 20556 17224 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 19426 20584 19432 20596
rect 19387 20556 19432 20584
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 20717 20587 20775 20593
rect 20717 20553 20729 20587
rect 20763 20584 20775 20587
rect 21818 20584 21824 20596
rect 20763 20556 21824 20584
rect 20763 20553 20775 20556
rect 20717 20547 20775 20553
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 31018 20584 31024 20596
rect 30979 20556 31024 20584
rect 31018 20544 31024 20556
rect 31076 20544 31082 20596
rect 3513 20519 3571 20525
rect 3513 20516 3525 20519
rect 2792 20488 3525 20516
rect 2792 20460 2820 20488
rect 3513 20485 3525 20488
rect 3559 20485 3571 20519
rect 3513 20479 3571 20485
rect 3697 20519 3755 20525
rect 3697 20485 3709 20519
rect 3743 20485 3755 20519
rect 3697 20479 3755 20485
rect 16574 20476 16580 20528
rect 16632 20516 16638 20528
rect 16669 20519 16727 20525
rect 16669 20516 16681 20519
rect 16632 20488 16681 20516
rect 16632 20476 16638 20488
rect 16669 20485 16681 20488
rect 16715 20485 16727 20519
rect 16669 20479 16727 20485
rect 23290 20476 23296 20528
rect 23348 20516 23354 20528
rect 24489 20519 24547 20525
rect 24489 20516 24501 20519
rect 23348 20488 24501 20516
rect 23348 20476 23354 20488
rect 24489 20485 24501 20488
rect 24535 20485 24547 20519
rect 24489 20479 24547 20485
rect 30098 20476 30104 20528
rect 30156 20516 30162 20528
rect 34425 20519 34483 20525
rect 34425 20516 34437 20519
rect 30156 20488 34437 20516
rect 30156 20476 30162 20488
rect 34425 20485 34437 20488
rect 34471 20485 34483 20519
rect 36078 20516 36084 20528
rect 34425 20479 34483 20485
rect 34716 20488 36084 20516
rect 34716 20460 34744 20488
rect 36078 20476 36084 20488
rect 36136 20476 36142 20528
rect 1394 20448 1400 20460
rect 1355 20420 1400 20448
rect 1394 20408 1400 20420
rect 1452 20408 1458 20460
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 2409 20451 2467 20457
rect 2409 20448 2421 20451
rect 1636 20420 2421 20448
rect 1636 20408 1642 20420
rect 2409 20417 2421 20420
rect 2455 20448 2467 20451
rect 2590 20448 2596 20460
rect 2455 20420 2596 20448
rect 2455 20417 2467 20420
rect 2409 20411 2467 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 2774 20448 2780 20460
rect 2735 20420 2780 20448
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20417 2927 20451
rect 2869 20411 2927 20417
rect 7837 20451 7895 20457
rect 7837 20417 7849 20451
rect 7883 20448 7895 20451
rect 7926 20448 7932 20460
rect 7883 20420 7932 20448
rect 7883 20417 7895 20420
rect 7837 20411 7895 20417
rect 1581 20315 1639 20321
rect 1581 20281 1593 20315
rect 1627 20312 1639 20315
rect 1854 20312 1860 20324
rect 1627 20284 1860 20312
rect 1627 20281 1639 20284
rect 1581 20275 1639 20281
rect 1854 20272 1860 20284
rect 1912 20312 1918 20324
rect 2884 20312 2912 20411
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 16942 20448 16948 20460
rect 16903 20420 16948 20448
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 18748 20420 19533 20448
rect 18748 20408 18754 20420
rect 19521 20417 19533 20420
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20438 20448 20444 20460
rect 20303 20420 20444 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20714 20448 20720 20460
rect 20579 20420 20720 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 24673 20451 24731 20457
rect 24673 20417 24685 20451
rect 24719 20448 24731 20451
rect 28258 20448 28264 20460
rect 24719 20420 28264 20448
rect 24719 20417 24731 20420
rect 24673 20411 24731 20417
rect 28258 20408 28264 20420
rect 28316 20408 28322 20460
rect 30374 20448 30380 20460
rect 30335 20420 30380 20448
rect 30374 20408 30380 20420
rect 30432 20408 30438 20460
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 31205 20451 31263 20457
rect 31205 20448 31217 20451
rect 30607 20420 31217 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 31205 20417 31217 20420
rect 31251 20417 31263 20451
rect 31205 20411 31263 20417
rect 34609 20451 34667 20457
rect 34609 20417 34621 20451
rect 34655 20417 34667 20451
rect 34609 20411 34667 20417
rect 12986 20340 12992 20392
rect 13044 20380 13050 20392
rect 14369 20383 14427 20389
rect 14369 20380 14381 20383
rect 13044 20352 14381 20380
rect 13044 20340 13050 20352
rect 14369 20349 14381 20352
rect 14415 20349 14427 20383
rect 15838 20380 15844 20392
rect 15799 20352 15844 20380
rect 14369 20343 14427 20349
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 16117 20383 16175 20389
rect 16117 20349 16129 20383
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 1912 20284 2912 20312
rect 16132 20312 16160 20343
rect 16482 20340 16488 20392
rect 16540 20380 16546 20392
rect 16761 20383 16819 20389
rect 16761 20380 16773 20383
rect 16540 20352 16773 20380
rect 16540 20340 16546 20352
rect 16761 20349 16773 20352
rect 16807 20349 16819 20383
rect 16761 20343 16819 20349
rect 19426 20340 19432 20392
rect 19484 20380 19490 20392
rect 20070 20380 20076 20392
rect 19484 20352 20076 20380
rect 19484 20340 19490 20352
rect 20070 20340 20076 20352
rect 20128 20380 20134 20392
rect 20349 20383 20407 20389
rect 20349 20380 20361 20383
rect 20128 20352 20361 20380
rect 20128 20340 20134 20352
rect 20349 20349 20361 20352
rect 20395 20349 20407 20383
rect 20349 20343 20407 20349
rect 24213 20383 24271 20389
rect 24213 20349 24225 20383
rect 24259 20380 24271 20383
rect 27430 20380 27436 20392
rect 24259 20352 27436 20380
rect 24259 20349 24271 20352
rect 24213 20343 24271 20349
rect 27430 20340 27436 20352
rect 27488 20340 27494 20392
rect 30193 20383 30251 20389
rect 30193 20349 30205 20383
rect 30239 20380 30251 20383
rect 30282 20380 30288 20392
rect 30239 20352 30288 20380
rect 30239 20349 30251 20352
rect 30193 20343 30251 20349
rect 30282 20340 30288 20352
rect 30340 20340 30346 20392
rect 34624 20380 34652 20411
rect 34698 20408 34704 20460
rect 34756 20448 34762 20460
rect 35253 20451 35311 20457
rect 34756 20420 34801 20448
rect 34756 20408 34762 20420
rect 35253 20417 35265 20451
rect 35299 20417 35311 20451
rect 35434 20448 35440 20460
rect 35395 20420 35440 20448
rect 35253 20411 35311 20417
rect 35268 20380 35296 20411
rect 35434 20408 35440 20420
rect 35492 20408 35498 20460
rect 35710 20380 35716 20392
rect 34624 20352 35716 20380
rect 35710 20340 35716 20352
rect 35768 20380 35774 20392
rect 36354 20380 36360 20392
rect 35768 20352 36360 20380
rect 35768 20340 35774 20352
rect 36354 20340 36360 20352
rect 36412 20340 36418 20392
rect 18506 20312 18512 20324
rect 16132 20284 18512 20312
rect 1912 20272 1918 20284
rect 18506 20272 18512 20284
rect 18564 20272 18570 20324
rect 21910 20312 21916 20324
rect 21871 20284 21916 20312
rect 21910 20272 21916 20284
rect 21968 20272 21974 20324
rect 2498 20244 2504 20256
rect 2459 20216 2504 20244
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 3053 20247 3111 20253
rect 3053 20213 3065 20247
rect 3099 20244 3111 20247
rect 3234 20244 3240 20256
rect 3099 20216 3240 20244
rect 3099 20213 3111 20216
rect 3053 20207 3111 20213
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 3786 20204 3792 20256
rect 3844 20244 3850 20256
rect 3881 20247 3939 20253
rect 3881 20244 3893 20247
rect 3844 20216 3893 20244
rect 3844 20204 3850 20216
rect 3881 20213 3893 20216
rect 3927 20213 3939 20247
rect 4706 20244 4712 20256
rect 4667 20216 4712 20244
rect 3881 20207 3939 20213
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7653 20247 7711 20253
rect 7653 20244 7665 20247
rect 7432 20216 7665 20244
rect 7432 20204 7438 20216
rect 7653 20213 7665 20216
rect 7699 20213 7711 20247
rect 7653 20207 7711 20213
rect 10505 20247 10563 20253
rect 10505 20213 10517 20247
rect 10551 20244 10563 20247
rect 12066 20244 12072 20256
rect 10551 20216 12072 20244
rect 10551 20213 10563 20216
rect 10505 20207 10563 20213
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 18782 20244 18788 20256
rect 18743 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 20533 20247 20591 20253
rect 20533 20213 20545 20247
rect 20579 20244 20591 20247
rect 20898 20244 20904 20256
rect 20579 20216 20904 20244
rect 20579 20213 20591 20216
rect 20533 20207 20591 20213
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 35345 20247 35403 20253
rect 35345 20213 35357 20247
rect 35391 20244 35403 20247
rect 35894 20244 35900 20256
rect 35391 20216 35900 20244
rect 35391 20213 35403 20216
rect 35345 20207 35403 20213
rect 35894 20204 35900 20216
rect 35952 20204 35958 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2958 20000 2964 20052
rect 3016 20040 3022 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3016 20012 3801 20040
rect 3016 20000 3022 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13814 20040 13820 20052
rect 13403 20012 13820 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14660 20012 16620 20040
rect 3050 19932 3056 19984
rect 3108 19972 3114 19984
rect 3145 19975 3203 19981
rect 3145 19972 3157 19975
rect 3108 19944 3157 19972
rect 3108 19932 3114 19944
rect 3145 19941 3157 19944
rect 3191 19972 3203 19975
rect 3191 19944 3924 19972
rect 3191 19941 3203 19944
rect 3145 19935 3203 19941
rect 3896 19913 3924 19944
rect 10318 19932 10324 19984
rect 10376 19972 10382 19984
rect 12434 19972 12440 19984
rect 10376 19944 12440 19972
rect 10376 19932 10382 19944
rect 12434 19932 12440 19944
rect 12492 19972 12498 19984
rect 14660 19972 14688 20012
rect 12492 19944 14688 19972
rect 12492 19932 12498 19944
rect 14734 19932 14740 19984
rect 14792 19972 14798 19984
rect 16592 19972 16620 20012
rect 16666 20000 16672 20052
rect 16724 20040 16730 20052
rect 18049 20043 18107 20049
rect 18049 20040 18061 20043
rect 16724 20012 18061 20040
rect 16724 20000 16730 20012
rect 18049 20009 18061 20012
rect 18095 20009 18107 20043
rect 18049 20003 18107 20009
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18472 20012 18521 20040
rect 18472 20000 18478 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 20898 20040 20904 20052
rect 20859 20012 20904 20040
rect 18509 20003 18567 20009
rect 20898 20000 20904 20012
rect 20956 20000 20962 20052
rect 37642 20040 37648 20052
rect 35636 20012 37136 20040
rect 37603 20012 37648 20040
rect 35636 19984 35664 20012
rect 18690 19972 18696 19984
rect 14792 19944 16068 19972
rect 16592 19944 18696 19972
rect 14792 19932 14798 19944
rect 3881 19907 3939 19913
rect 3881 19873 3893 19907
rect 3927 19873 3939 19907
rect 4706 19904 4712 19916
rect 4667 19876 4712 19904
rect 3881 19867 3939 19873
rect 4706 19864 4712 19876
rect 4764 19864 4770 19916
rect 4890 19904 4896 19916
rect 4851 19876 4896 19904
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 4982 19864 4988 19916
rect 5040 19904 5046 19916
rect 11882 19904 11888 19916
rect 5040 19876 11888 19904
rect 5040 19864 5046 19876
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12066 19904 12072 19916
rect 12027 19876 12072 19904
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12986 19864 12992 19916
rect 13044 19904 13050 19916
rect 13173 19907 13231 19913
rect 13173 19904 13185 19907
rect 13044 19876 13185 19904
rect 13044 19864 13050 19876
rect 13173 19873 13185 19876
rect 13219 19873 13231 19907
rect 13173 19867 13231 19873
rect 15013 19907 15071 19913
rect 15013 19873 15025 19907
rect 15059 19904 15071 19907
rect 15838 19904 15844 19916
rect 15059 19876 15844 19904
rect 15059 19873 15071 19876
rect 15013 19867 15071 19873
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 16040 19913 16068 19944
rect 18690 19932 18696 19944
rect 18748 19932 18754 19984
rect 19429 19975 19487 19981
rect 19429 19941 19441 19975
rect 19475 19941 19487 19975
rect 19429 19935 19487 19941
rect 20257 19975 20315 19981
rect 20257 19941 20269 19975
rect 20303 19972 20315 19975
rect 20714 19972 20720 19984
rect 20303 19944 20720 19972
rect 20303 19941 20315 19944
rect 20257 19935 20315 19941
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16114 19904 16120 19916
rect 16071 19876 16120 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16114 19864 16120 19876
rect 16172 19904 16178 19916
rect 16761 19907 16819 19913
rect 16761 19904 16773 19907
rect 16172 19876 16773 19904
rect 16172 19864 16178 19876
rect 16761 19873 16773 19876
rect 16807 19873 16819 19907
rect 18138 19904 18144 19916
rect 18099 19876 18144 19904
rect 16761 19867 16819 19873
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 2958 19836 2964 19848
rect 2919 19808 2964 19836
rect 2958 19796 2964 19808
rect 3016 19796 3022 19848
rect 3234 19796 3240 19848
rect 3292 19836 3298 19848
rect 3786 19836 3792 19848
rect 3292 19808 3337 19836
rect 3747 19808 3792 19836
rect 3292 19796 3298 19808
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 4065 19839 4123 19845
rect 4065 19836 4077 19839
rect 3896 19808 4077 19836
rect 2590 19728 2596 19780
rect 2648 19768 2654 19780
rect 3896 19768 3924 19808
rect 4065 19805 4077 19808
rect 4111 19805 4123 19839
rect 13078 19836 13084 19848
rect 13039 19808 13084 19836
rect 4065 19799 4123 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 13872 19808 14749 19836
rect 13872 19796 13878 19808
rect 14737 19805 14749 19808
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19836 16359 19839
rect 16347 19808 16528 19836
rect 16347 19805 16359 19808
rect 16301 19799 16359 19805
rect 2648 19740 3924 19768
rect 2648 19728 2654 19740
rect 3970 19728 3976 19780
rect 4028 19768 4034 19780
rect 6549 19771 6607 19777
rect 6549 19768 6561 19771
rect 4028 19740 6561 19768
rect 4028 19728 4034 19740
rect 6549 19737 6561 19740
rect 6595 19768 6607 19771
rect 10229 19771 10287 19777
rect 10229 19768 10241 19771
rect 6595 19740 10241 19768
rect 6595 19737 6607 19740
rect 6549 19731 6607 19737
rect 10229 19737 10241 19740
rect 10275 19768 10287 19771
rect 10962 19768 10968 19780
rect 10275 19740 10968 19768
rect 10275 19737 10287 19740
rect 10229 19731 10287 19737
rect 10962 19728 10968 19740
rect 11020 19728 11026 19780
rect 11790 19728 11796 19780
rect 11848 19768 11854 19780
rect 11885 19771 11943 19777
rect 11885 19768 11897 19771
rect 11848 19740 11897 19768
rect 11848 19728 11854 19740
rect 11885 19737 11897 19740
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 1946 19700 1952 19712
rect 1907 19672 1952 19700
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 2777 19703 2835 19709
rect 2777 19669 2789 19703
rect 2823 19700 2835 19703
rect 4062 19700 4068 19712
rect 2823 19672 4068 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4249 19703 4307 19709
rect 4249 19669 4261 19703
rect 4295 19700 4307 19703
rect 4614 19700 4620 19712
rect 4295 19672 4620 19700
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 12897 19703 12955 19709
rect 12897 19700 12909 19703
rect 11664 19672 12909 19700
rect 11664 19660 11670 19672
rect 12897 19669 12909 19672
rect 12943 19669 12955 19703
rect 16500 19700 16528 19808
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 17000 19808 17049 19836
rect 17000 19796 17006 19808
rect 17037 19805 17049 19808
rect 17083 19836 17095 19839
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 17083 19808 18337 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18840 19808 19257 19836
rect 18840 19796 18846 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19444 19836 19472 19935
rect 20714 19932 20720 19944
rect 20772 19932 20778 19984
rect 32582 19972 32588 19984
rect 22066 19944 32588 19972
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 22066 19904 22094 19944
rect 32582 19932 32588 19944
rect 32640 19932 32646 19984
rect 35618 19972 35624 19984
rect 35452 19944 35624 19972
rect 20220 19876 22094 19904
rect 23845 19907 23903 19913
rect 20220 19864 20226 19876
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 25222 19904 25228 19916
rect 23891 19876 25228 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 25222 19864 25228 19876
rect 25280 19904 25286 19916
rect 28810 19904 28816 19916
rect 25280 19876 28816 19904
rect 25280 19864 25286 19876
rect 28810 19864 28816 19876
rect 28868 19864 28874 19916
rect 30282 19904 30288 19916
rect 30243 19876 30288 19904
rect 30282 19864 30288 19876
rect 30340 19864 30346 19916
rect 20530 19836 20536 19848
rect 19444 19808 20536 19836
rect 19245 19799 19303 19805
rect 20530 19796 20536 19808
rect 20588 19836 20594 19848
rect 21453 19839 21511 19845
rect 21453 19836 21465 19839
rect 20588 19808 21465 19836
rect 20588 19796 20594 19808
rect 21453 19805 21465 19808
rect 21499 19805 21511 19839
rect 21453 19799 21511 19805
rect 21910 19796 21916 19848
rect 21968 19836 21974 19848
rect 35452 19845 35480 19944
rect 35618 19932 35624 19944
rect 35676 19932 35682 19984
rect 37001 19975 37059 19981
rect 37001 19972 37013 19975
rect 35866 19944 37013 19972
rect 35866 19904 35894 19944
rect 37001 19941 37013 19944
rect 37047 19941 37059 19975
rect 37001 19935 37059 19941
rect 35820 19876 35894 19904
rect 35710 19845 35716 19848
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21968 19808 22109 19836
rect 21968 19796 21974 19808
rect 22097 19805 22109 19808
rect 22143 19805 22155 19839
rect 22097 19799 22155 19805
rect 27433 19839 27491 19845
rect 27433 19805 27445 19839
rect 27479 19836 27491 19839
rect 30469 19839 30527 19845
rect 27479 19808 28028 19836
rect 27479 19805 27491 19808
rect 27433 19799 27491 19805
rect 16574 19728 16580 19780
rect 16632 19768 16638 19780
rect 18049 19771 18107 19777
rect 18049 19768 18061 19771
rect 16632 19740 18061 19768
rect 16632 19728 16638 19740
rect 18049 19737 18061 19740
rect 18095 19737 18107 19771
rect 18049 19731 18107 19737
rect 18414 19728 18420 19780
rect 18472 19768 18478 19780
rect 20073 19771 20131 19777
rect 20073 19768 20085 19771
rect 18472 19740 20085 19768
rect 18472 19728 18478 19740
rect 20073 19737 20085 19740
rect 20119 19737 20131 19771
rect 20073 19731 20131 19737
rect 20809 19771 20867 19777
rect 20809 19737 20821 19771
rect 20855 19737 20867 19771
rect 20809 19731 20867 19737
rect 18432 19700 18460 19728
rect 16500 19672 18460 19700
rect 12897 19663 12955 19669
rect 18506 19660 18512 19712
rect 18564 19700 18570 19712
rect 20824 19700 20852 19731
rect 25406 19728 25412 19780
rect 25464 19768 25470 19780
rect 25593 19771 25651 19777
rect 25593 19768 25605 19771
rect 25464 19740 25605 19768
rect 25464 19728 25470 19740
rect 25593 19737 25605 19740
rect 25639 19768 25651 19771
rect 26326 19768 26332 19780
rect 25639 19740 26332 19768
rect 25639 19737 25651 19740
rect 25593 19731 25651 19737
rect 26326 19728 26332 19740
rect 26384 19728 26390 19780
rect 27246 19768 27252 19780
rect 27207 19740 27252 19768
rect 27246 19728 27252 19740
rect 27304 19728 27310 19780
rect 18564 19672 20852 19700
rect 21637 19703 21695 19709
rect 18564 19660 18570 19672
rect 21637 19669 21649 19703
rect 21683 19700 21695 19703
rect 22094 19700 22100 19712
rect 21683 19672 22100 19700
rect 21683 19669 21695 19672
rect 21637 19663 21695 19669
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 28000 19709 28028 19808
rect 30469 19805 30481 19839
rect 30515 19805 30527 19839
rect 30469 19799 30527 19805
rect 35437 19839 35495 19845
rect 35437 19805 35449 19839
rect 35483 19805 35495 19839
rect 35437 19799 35495 19805
rect 35667 19839 35716 19845
rect 35667 19805 35679 19839
rect 35713 19805 35716 19839
rect 35667 19799 35716 19805
rect 29730 19728 29736 19780
rect 29788 19768 29794 19780
rect 30484 19768 30512 19799
rect 35710 19796 35716 19799
rect 35768 19796 35774 19848
rect 35820 19845 35848 19876
rect 35805 19839 35863 19845
rect 35805 19805 35817 19839
rect 35851 19805 35863 19839
rect 35805 19799 35863 19805
rect 35897 19839 35955 19845
rect 35897 19805 35909 19839
rect 35943 19836 35955 19839
rect 36078 19836 36084 19848
rect 35943 19808 36084 19836
rect 35943 19805 35955 19808
rect 35897 19799 35955 19805
rect 36078 19796 36084 19808
rect 36136 19796 36142 19848
rect 36354 19836 36360 19848
rect 36315 19808 36360 19836
rect 36354 19796 36360 19808
rect 36412 19796 36418 19848
rect 37001 19839 37059 19845
rect 37001 19805 37013 19839
rect 37047 19836 37059 19839
rect 37108 19836 37136 20012
rect 37642 20000 37648 20012
rect 37700 20000 37706 20052
rect 37047 19808 37136 19836
rect 37185 19839 37243 19845
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 37185 19805 37197 19839
rect 37231 19836 37243 19839
rect 37642 19836 37648 19848
rect 37231 19808 37648 19836
rect 37231 19805 37243 19808
rect 37185 19799 37243 19805
rect 37642 19796 37648 19808
rect 37700 19796 37706 19848
rect 29788 19740 30512 19768
rect 30653 19771 30711 19777
rect 29788 19728 29794 19740
rect 30653 19737 30665 19771
rect 30699 19768 30711 19771
rect 32030 19768 32036 19780
rect 30699 19740 32036 19768
rect 30699 19737 30711 19740
rect 30653 19731 30711 19737
rect 32030 19728 32036 19740
rect 32088 19728 32094 19780
rect 35342 19728 35348 19780
rect 35400 19768 35406 19780
rect 35529 19771 35587 19777
rect 35529 19768 35541 19771
rect 35400 19740 35541 19768
rect 35400 19728 35406 19740
rect 35529 19737 35541 19740
rect 35575 19737 35587 19771
rect 35529 19731 35587 19737
rect 27985 19703 28043 19709
rect 27985 19669 27997 19703
rect 28031 19700 28043 19703
rect 30558 19700 30564 19712
rect 28031 19672 30564 19700
rect 28031 19669 28043 19672
rect 27985 19663 28043 19669
rect 30558 19660 30564 19672
rect 30616 19660 30622 19712
rect 31294 19700 31300 19712
rect 31255 19672 31300 19700
rect 31294 19660 31300 19672
rect 31352 19660 31358 19712
rect 34698 19660 34704 19712
rect 34756 19700 34762 19712
rect 35253 19703 35311 19709
rect 35253 19700 35265 19703
rect 34756 19672 35265 19700
rect 34756 19660 34762 19672
rect 35253 19669 35265 19672
rect 35299 19669 35311 19703
rect 35253 19663 35311 19669
rect 35710 19660 35716 19712
rect 35768 19700 35774 19712
rect 36449 19703 36507 19709
rect 36449 19700 36461 19703
rect 35768 19672 36461 19700
rect 35768 19660 35774 19672
rect 36449 19669 36461 19672
rect 36495 19669 36507 19703
rect 36449 19663 36507 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3513 19499 3571 19505
rect 3513 19465 3525 19499
rect 3559 19496 3571 19499
rect 4982 19496 4988 19508
rect 3559 19468 4988 19496
rect 3559 19465 3571 19468
rect 3513 19459 3571 19465
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 11790 19496 11796 19508
rect 11751 19468 11796 19496
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 11882 19456 11888 19508
rect 11940 19496 11946 19508
rect 11940 19468 18644 19496
rect 11940 19456 11946 19468
rect 2866 19388 2872 19440
rect 2924 19428 2930 19440
rect 3053 19431 3111 19437
rect 3053 19428 3065 19431
rect 2924 19400 3065 19428
rect 2924 19388 2930 19400
rect 3053 19397 3065 19400
rect 3099 19397 3111 19431
rect 3053 19391 3111 19397
rect 3602 19388 3608 19440
rect 3660 19428 3666 19440
rect 3970 19428 3976 19440
rect 3660 19400 3976 19428
rect 3660 19388 3666 19400
rect 3970 19388 3976 19400
rect 4028 19388 4034 19440
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 6730 19428 6736 19440
rect 4120 19400 6736 19428
rect 4120 19388 4126 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 7926 19388 7932 19440
rect 7984 19428 7990 19440
rect 9125 19431 9183 19437
rect 9125 19428 9137 19431
rect 7984 19400 9137 19428
rect 7984 19388 7990 19400
rect 9125 19397 9137 19400
rect 9171 19428 9183 19431
rect 10137 19431 10195 19437
rect 10137 19428 10149 19431
rect 9171 19400 10149 19428
rect 9171 19397 9183 19400
rect 9125 19391 9183 19397
rect 10137 19397 10149 19400
rect 10183 19397 10195 19431
rect 10318 19428 10324 19440
rect 10279 19400 10324 19428
rect 10137 19391 10195 19397
rect 10318 19388 10324 19400
rect 10376 19388 10382 19440
rect 12986 19388 12992 19440
rect 13044 19428 13050 19440
rect 13354 19428 13360 19440
rect 13044 19400 13216 19428
rect 13315 19400 13360 19428
rect 13044 19388 13050 19400
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 3329 19363 3387 19369
rect 3329 19360 3341 19363
rect 2004 19332 3341 19360
rect 2004 19320 2010 19332
rect 3329 19329 3341 19332
rect 3375 19360 3387 19363
rect 4154 19360 4160 19372
rect 3375 19332 4160 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 11606 19360 11612 19372
rect 11567 19332 11612 19360
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 13078 19360 13084 19372
rect 12991 19332 13084 19360
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 13188 19369 13216 19400
rect 13354 19388 13360 19400
rect 13412 19388 13418 19440
rect 13998 19428 14004 19440
rect 13959 19400 14004 19428
rect 13998 19388 14004 19400
rect 14056 19388 14062 19440
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 14700 19400 14964 19428
rect 14700 19388 14706 19400
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19360 13231 19363
rect 13906 19360 13912 19372
rect 13219 19332 13912 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 14936 19369 14964 19400
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 16669 19431 16727 19437
rect 16669 19428 16681 19431
rect 16632 19400 16681 19428
rect 16632 19388 16638 19400
rect 16669 19397 16681 19400
rect 16715 19397 16727 19431
rect 16669 19391 16727 19397
rect 18616 19428 18644 19468
rect 18690 19456 18696 19508
rect 18748 19496 18754 19508
rect 18785 19499 18843 19505
rect 18785 19496 18797 19499
rect 18748 19468 18797 19496
rect 18748 19456 18754 19468
rect 18785 19465 18797 19468
rect 18831 19496 18843 19499
rect 18966 19496 18972 19508
rect 18831 19468 18972 19496
rect 18831 19465 18843 19468
rect 18785 19459 18843 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 23293 19499 23351 19505
rect 23293 19465 23305 19499
rect 23339 19496 23351 19499
rect 24394 19496 24400 19508
rect 23339 19468 24400 19496
rect 23339 19465 23351 19468
rect 23293 19459 23351 19465
rect 24394 19456 24400 19468
rect 24452 19456 24458 19508
rect 24489 19499 24547 19505
rect 24489 19465 24501 19499
rect 24535 19465 24547 19499
rect 24489 19459 24547 19465
rect 25133 19499 25191 19505
rect 25133 19465 25145 19499
rect 25179 19496 25191 19499
rect 27246 19496 27252 19508
rect 25179 19468 27252 19496
rect 25179 19465 25191 19468
rect 25133 19459 25191 19465
rect 19429 19431 19487 19437
rect 19429 19428 19441 19431
rect 18616 19400 19441 19428
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 14921 19323 14979 19329
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16540 19332 16865 19360
rect 16540 19320 16546 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 18616 19369 18644 19400
rect 19429 19397 19441 19400
rect 19475 19397 19487 19431
rect 19429 19391 19487 19397
rect 19521 19431 19579 19437
rect 19521 19397 19533 19431
rect 19567 19428 19579 19431
rect 20254 19428 20260 19440
rect 19567 19400 20260 19428
rect 19567 19397 19579 19400
rect 19521 19391 19579 19397
rect 20254 19388 20260 19400
rect 20312 19388 20318 19440
rect 22833 19431 22891 19437
rect 22833 19397 22845 19431
rect 22879 19428 22891 19431
rect 22922 19428 22928 19440
rect 22879 19400 22928 19428
rect 22879 19397 22891 19400
rect 22833 19391 22891 19397
rect 22922 19388 22928 19400
rect 22980 19428 22986 19440
rect 24504 19428 24532 19459
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 29730 19496 29736 19508
rect 29691 19468 29736 19496
rect 29730 19456 29736 19468
rect 29788 19456 29794 19508
rect 30374 19496 30380 19508
rect 30335 19468 30380 19496
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 32122 19496 32128 19508
rect 31726 19468 32128 19496
rect 26970 19428 26976 19440
rect 22980 19400 23336 19428
rect 24504 19400 26976 19428
rect 22980 19388 22986 19400
rect 23308 19372 23336 19400
rect 26970 19388 26976 19400
rect 27028 19388 27034 19440
rect 29086 19388 29092 19440
rect 29144 19428 29150 19440
rect 29457 19431 29515 19437
rect 29457 19428 29469 19431
rect 29144 19400 29469 19428
rect 29144 19388 29150 19400
rect 29457 19397 29469 19400
rect 29503 19397 29515 19431
rect 29457 19391 29515 19397
rect 30098 19388 30104 19440
rect 30156 19428 30162 19440
rect 30837 19431 30895 19437
rect 30837 19428 30849 19431
rect 30156 19400 30849 19428
rect 30156 19388 30162 19400
rect 30837 19397 30849 19400
rect 30883 19428 30895 19431
rect 31726 19428 31754 19468
rect 32122 19456 32128 19468
rect 32180 19456 32186 19508
rect 34523 19499 34581 19505
rect 34523 19465 34535 19499
rect 34569 19496 34581 19499
rect 35342 19496 35348 19508
rect 34569 19468 35204 19496
rect 35303 19468 35348 19496
rect 34569 19465 34581 19468
rect 34523 19459 34581 19465
rect 30883 19400 31754 19428
rect 32217 19431 32275 19437
rect 30883 19397 30895 19400
rect 30837 19391 30895 19397
rect 32217 19397 32229 19431
rect 32263 19428 32275 19431
rect 34609 19431 34667 19437
rect 34609 19428 34621 19431
rect 32263 19400 34621 19428
rect 32263 19397 32275 19400
rect 32217 19391 32275 19397
rect 34609 19397 34621 19400
rect 34655 19397 34667 19431
rect 35176 19428 35204 19468
rect 35342 19456 35348 19468
rect 35400 19456 35406 19508
rect 35526 19456 35532 19508
rect 35584 19496 35590 19508
rect 36078 19496 36084 19508
rect 35584 19468 36084 19496
rect 35584 19456 35590 19468
rect 36078 19456 36084 19468
rect 36136 19456 36142 19508
rect 36446 19428 36452 19440
rect 35176 19400 36452 19428
rect 34609 19391 34667 19397
rect 36446 19388 36452 19400
rect 36504 19388 36510 19440
rect 18601 19363 18659 19369
rect 17000 19332 17045 19360
rect 17000 19320 17006 19332
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 20070 19360 20076 19372
rect 19659 19332 20076 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20162 19320 20168 19372
rect 20220 19360 20226 19372
rect 22189 19363 22247 19369
rect 20220 19332 20265 19360
rect 20220 19320 20226 19332
rect 22189 19329 22201 19363
rect 22235 19360 22247 19363
rect 22278 19360 22284 19372
rect 22235 19332 22284 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 22278 19320 22284 19332
rect 22336 19320 22342 19372
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19329 23167 19363
rect 23109 19323 23167 19329
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 3108 19264 3157 19292
rect 3108 19252 3114 19264
rect 3145 19261 3157 19264
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 13096 19224 13124 19320
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 14424 19264 14657 19292
rect 14424 19252 14430 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 19978 19292 19984 19304
rect 19939 19264 19984 19292
rect 14645 19255 14703 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 23014 19292 23020 19304
rect 22975 19264 23020 19292
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 23124 19224 23152 19323
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 24302 19360 24308 19372
rect 24263 19332 24308 19360
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 24394 19320 24400 19372
rect 24452 19360 24458 19372
rect 24949 19363 25007 19369
rect 24949 19360 24961 19363
rect 24452 19332 24961 19360
rect 24452 19320 24458 19332
rect 24949 19329 24961 19332
rect 24995 19329 25007 19363
rect 24949 19323 25007 19329
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19329 29239 19363
rect 29362 19360 29368 19372
rect 29323 19332 29368 19360
rect 29181 19323 29239 19329
rect 13096 19196 14872 19224
rect 14844 19168 14872 19196
rect 22388 19196 23152 19224
rect 28721 19227 28779 19233
rect 22388 19168 22416 19196
rect 28721 19193 28733 19227
rect 28767 19224 28779 19227
rect 29196 19224 29224 19323
rect 29362 19320 29368 19332
rect 29420 19320 29426 19372
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19360 29607 19363
rect 30006 19360 30012 19372
rect 29595 19332 30012 19360
rect 29595 19329 29607 19332
rect 29549 19323 29607 19329
rect 30006 19320 30012 19332
rect 30064 19320 30070 19372
rect 30745 19363 30803 19369
rect 30745 19329 30757 19363
rect 30791 19360 30803 19363
rect 31294 19360 31300 19372
rect 30791 19332 31300 19360
rect 30791 19329 30803 19332
rect 30745 19323 30803 19329
rect 31294 19320 31300 19332
rect 31352 19320 31358 19372
rect 32122 19360 32128 19372
rect 32083 19332 32128 19360
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19360 32370 19372
rect 32769 19363 32827 19369
rect 32769 19360 32781 19363
rect 32364 19332 32781 19360
rect 32364 19320 32370 19332
rect 32769 19329 32781 19332
rect 32815 19329 32827 19363
rect 34425 19363 34483 19369
rect 34425 19360 34437 19363
rect 32769 19323 32827 19329
rect 33888 19332 34437 19360
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 30190 19292 30196 19304
rect 29880 19264 30196 19292
rect 29880 19252 29886 19264
rect 30190 19252 30196 19264
rect 30248 19292 30254 19304
rect 30929 19295 30987 19301
rect 30929 19292 30941 19295
rect 30248 19264 30941 19292
rect 30248 19252 30254 19264
rect 30929 19261 30941 19264
rect 30975 19261 30987 19295
rect 30929 19255 30987 19261
rect 30006 19224 30012 19236
rect 28767 19196 30012 19224
rect 28767 19193 28779 19196
rect 28721 19187 28779 19193
rect 30006 19184 30012 19196
rect 30064 19184 30070 19236
rect 33888 19233 33916 19332
rect 34425 19329 34437 19332
rect 34471 19329 34483 19363
rect 34425 19323 34483 19329
rect 34698 19320 34704 19372
rect 34756 19360 34762 19372
rect 35161 19363 35219 19369
rect 34756 19332 34801 19360
rect 34756 19320 34762 19332
rect 35161 19329 35173 19363
rect 35207 19329 35219 19363
rect 35161 19323 35219 19329
rect 35345 19363 35403 19369
rect 35345 19329 35357 19363
rect 35391 19360 35403 19363
rect 35710 19360 35716 19372
rect 35391 19332 35716 19360
rect 35391 19329 35403 19332
rect 35345 19323 35403 19329
rect 35176 19292 35204 19323
rect 35710 19320 35716 19332
rect 35768 19320 35774 19372
rect 35434 19292 35440 19304
rect 35176 19264 35440 19292
rect 35434 19252 35440 19264
rect 35492 19252 35498 19304
rect 33873 19227 33931 19233
rect 33873 19224 33885 19227
rect 31726 19196 33885 19224
rect 2958 19116 2964 19168
rect 3016 19156 3022 19168
rect 3053 19159 3111 19165
rect 3053 19156 3065 19159
rect 3016 19128 3065 19156
rect 3016 19116 3022 19128
rect 3053 19125 3065 19128
rect 3099 19125 3111 19159
rect 3053 19119 3111 19125
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 4890 19156 4896 19168
rect 4764 19128 4896 19156
rect 4764 19116 4770 19128
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 6454 19156 6460 19168
rect 6415 19128 6460 19156
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 9030 19156 9036 19168
rect 8991 19128 9036 19156
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 12894 19156 12900 19168
rect 12855 19128 12900 19156
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 13357 19159 13415 19165
rect 13357 19125 13369 19159
rect 13403 19156 13415 19159
rect 13814 19156 13820 19168
rect 13403 19128 13820 19156
rect 13403 19125 13415 19128
rect 13357 19119 13415 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 14056 19128 14105 19156
rect 14056 19116 14062 19128
rect 14093 19125 14105 19128
rect 14139 19125 14151 19159
rect 14093 19119 14151 19125
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 14884 19128 15945 19156
rect 14884 19116 14890 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16632 19128 16681 19156
rect 16632 19116 16638 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 17126 19156 17132 19168
rect 17087 19128 17132 19156
rect 16669 19119 16727 19125
rect 17126 19116 17132 19128
rect 17184 19116 17190 19168
rect 17957 19159 18015 19165
rect 17957 19125 17969 19159
rect 18003 19156 18015 19159
rect 18138 19156 18144 19168
rect 18003 19128 18144 19156
rect 18003 19125 18015 19128
rect 17957 19119 18015 19125
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 22370 19156 22376 19168
rect 22331 19128 22376 19156
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 22830 19156 22836 19168
rect 22791 19128 22836 19156
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 31726 19156 31754 19196
rect 33873 19193 33885 19196
rect 33919 19193 33931 19227
rect 33873 19187 33931 19193
rect 28684 19128 31754 19156
rect 28684 19116 28690 19128
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18952 4123 18955
rect 4111 18924 6914 18952
rect 4111 18921 4123 18924
rect 4065 18915 4123 18921
rect 4249 18887 4307 18893
rect 4249 18853 4261 18887
rect 4295 18884 4307 18887
rect 5537 18887 5595 18893
rect 4295 18856 5212 18884
rect 4295 18853 4307 18856
rect 4249 18847 4307 18853
rect 4154 18816 4160 18828
rect 4115 18788 4160 18816
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 4378 18819 4436 18825
rect 4378 18785 4390 18819
rect 4424 18816 4436 18819
rect 4706 18816 4712 18828
rect 4424 18788 4712 18816
rect 4424 18785 4436 18788
rect 4378 18779 4436 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 5184 18760 5212 18856
rect 5537 18853 5549 18887
rect 5583 18884 5595 18887
rect 5626 18884 5632 18896
rect 5583 18856 5632 18884
rect 5583 18853 5595 18856
rect 5537 18847 5595 18853
rect 5626 18844 5632 18856
rect 5684 18844 5690 18896
rect 6886 18816 6914 18924
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 9088 18924 21465 18952
rect 9088 18912 9094 18924
rect 21453 18921 21465 18924
rect 21499 18952 21511 18955
rect 21910 18952 21916 18964
rect 21499 18924 21916 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 22830 18952 22836 18964
rect 22152 18924 22836 18952
rect 22152 18912 22158 18924
rect 22830 18912 22836 18924
rect 22888 18952 22894 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22888 18924 22937 18952
rect 22888 18912 22894 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23385 18955 23443 18961
rect 23385 18921 23397 18955
rect 23431 18952 23443 18955
rect 24302 18952 24308 18964
rect 23431 18924 24308 18952
rect 23431 18921 23443 18924
rect 23385 18915 23443 18921
rect 24302 18912 24308 18924
rect 24360 18912 24366 18964
rect 31573 18955 31631 18961
rect 31573 18921 31585 18955
rect 31619 18952 31631 18955
rect 32122 18952 32128 18964
rect 31619 18924 32128 18952
rect 31619 18921 31631 18924
rect 31573 18915 31631 18921
rect 32122 18912 32128 18924
rect 32180 18912 32186 18964
rect 35434 18952 35440 18964
rect 35395 18924 35440 18952
rect 35434 18912 35440 18924
rect 35492 18912 35498 18964
rect 37642 18912 37648 18964
rect 37700 18952 37706 18964
rect 37737 18955 37795 18961
rect 37737 18952 37749 18955
rect 37700 18924 37749 18952
rect 37700 18912 37706 18924
rect 37737 18921 37749 18924
rect 37783 18921 37795 18955
rect 37737 18915 37795 18921
rect 26326 18884 26332 18896
rect 12406 18856 19334 18884
rect 12406 18816 12434 18856
rect 6886 18788 12434 18816
rect 14642 18776 14648 18828
rect 14700 18816 14706 18828
rect 15013 18819 15071 18825
rect 15013 18816 15025 18819
rect 14700 18788 15025 18816
rect 14700 18776 14706 18788
rect 15013 18785 15025 18788
rect 15059 18785 15071 18819
rect 19306 18816 19334 18856
rect 22020 18856 26332 18884
rect 22020 18816 22048 18856
rect 26326 18844 26332 18856
rect 26384 18844 26390 18896
rect 19306 18788 22048 18816
rect 15013 18779 15071 18785
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22189 18819 22247 18825
rect 22189 18816 22201 18819
rect 22152 18788 22201 18816
rect 22152 18776 22158 18788
rect 22189 18785 22201 18788
rect 22235 18816 22247 18819
rect 23014 18816 23020 18828
rect 22235 18788 23020 18816
rect 22235 18785 22247 18788
rect 22189 18779 22247 18785
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 25777 18819 25835 18825
rect 25777 18785 25789 18819
rect 25823 18785 25835 18819
rect 26970 18816 26976 18828
rect 26931 18788 26976 18816
rect 25777 18779 25835 18785
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18748 1458 18760
rect 2041 18751 2099 18757
rect 2041 18748 2053 18751
rect 1452 18720 2053 18748
rect 1452 18708 1458 18720
rect 2041 18717 2053 18720
rect 2087 18717 2099 18751
rect 2041 18711 2099 18717
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4614 18748 4620 18760
rect 4571 18720 4620 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5224 18720 5365 18748
rect 5224 18708 5230 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18748 6883 18751
rect 7098 18748 7104 18760
rect 6871 18720 7104 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 7098 18708 7104 18720
rect 7156 18748 7162 18760
rect 7285 18751 7343 18757
rect 7285 18748 7297 18751
rect 7156 18720 7297 18748
rect 7156 18708 7162 18720
rect 7285 18717 7297 18720
rect 7331 18717 7343 18751
rect 7285 18711 7343 18717
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 10367 18720 10793 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10781 18717 10793 18720
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 15252 18720 15301 18748
rect 15252 18708 15258 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15896 18720 16405 18748
rect 15896 18708 15902 18720
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 18739 18720 19533 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 19521 18717 19533 18720
rect 19567 18748 19579 18751
rect 20162 18748 20168 18760
rect 19567 18720 20168 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 21910 18708 21916 18760
rect 21968 18748 21974 18760
rect 22005 18751 22063 18757
rect 22005 18748 22017 18751
rect 21968 18720 22017 18748
rect 21968 18708 21974 18720
rect 22005 18717 22017 18720
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18748 22339 18751
rect 22370 18748 22376 18760
rect 22327 18720 22376 18748
rect 22327 18717 22339 18720
rect 22281 18711 22339 18717
rect 6454 18640 6460 18692
rect 6512 18680 6518 18692
rect 6641 18683 6699 18689
rect 6641 18680 6653 18683
rect 6512 18652 6653 18680
rect 6512 18640 6518 18652
rect 6641 18649 6653 18652
rect 6687 18680 6699 18683
rect 9766 18680 9772 18692
rect 6687 18652 9772 18680
rect 6687 18649 6699 18652
rect 6641 18643 6699 18649
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 10965 18683 11023 18689
rect 10965 18649 10977 18683
rect 11011 18680 11023 18683
rect 11974 18680 11980 18692
rect 11011 18652 11980 18680
rect 11011 18649 11023 18652
rect 10965 18643 11023 18649
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 12621 18683 12679 18689
rect 12621 18680 12633 18683
rect 12308 18652 12633 18680
rect 12308 18640 12314 18652
rect 12621 18649 12633 18652
rect 12667 18649 12679 18683
rect 16574 18680 16580 18692
rect 16535 18652 16580 18680
rect 12621 18643 12679 18649
rect 16574 18640 16580 18652
rect 16632 18640 16638 18692
rect 22020 18680 22048 18711
rect 22370 18708 22376 18720
rect 22428 18748 22434 18760
rect 23106 18748 23112 18760
rect 22428 18720 23112 18748
rect 22428 18708 22434 18720
rect 23106 18708 23112 18720
rect 23164 18748 23170 18760
rect 23201 18751 23259 18757
rect 23201 18748 23213 18751
rect 23164 18720 23213 18748
rect 23164 18708 23170 18720
rect 23201 18717 23213 18720
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 22830 18680 22836 18692
rect 19352 18652 21588 18680
rect 22020 18652 22836 18680
rect 7466 18612 7472 18624
rect 7427 18584 7472 18612
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 19352 18621 19380 18652
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 14424 18584 14473 18612
rect 14424 18572 14430 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 14461 18575 14519 18581
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18581 19395 18615
rect 20070 18612 20076 18624
rect 20031 18584 20076 18612
rect 19337 18575 19395 18581
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 21560 18612 21588 18652
rect 22830 18640 22836 18652
rect 22888 18640 22894 18692
rect 22925 18683 22983 18689
rect 22925 18649 22937 18683
rect 22971 18680 22983 18683
rect 23290 18680 23296 18692
rect 22971 18652 23296 18680
rect 22971 18649 22983 18652
rect 22925 18643 22983 18649
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 25792 18680 25820 18779
rect 26970 18776 26976 18788
rect 27028 18776 27034 18828
rect 30558 18776 30564 18828
rect 30616 18816 30622 18828
rect 30929 18819 30987 18825
rect 30929 18816 30941 18819
rect 30616 18788 30941 18816
rect 30616 18776 30622 18788
rect 30929 18785 30941 18788
rect 30975 18816 30987 18819
rect 33229 18819 33287 18825
rect 33229 18816 33241 18819
rect 30975 18788 33241 18816
rect 30975 18785 30987 18788
rect 30929 18779 30987 18785
rect 33229 18785 33241 18788
rect 33275 18816 33287 18819
rect 34057 18819 34115 18825
rect 34057 18816 34069 18819
rect 33275 18788 34069 18816
rect 33275 18785 33287 18788
rect 33229 18779 33287 18785
rect 34057 18785 34069 18788
rect 34103 18816 34115 18819
rect 34793 18819 34851 18825
rect 34793 18816 34805 18819
rect 34103 18788 34805 18816
rect 34103 18785 34115 18788
rect 34057 18779 34115 18785
rect 34793 18785 34805 18788
rect 34839 18785 34851 18819
rect 34793 18779 34851 18785
rect 27157 18751 27215 18757
rect 27157 18717 27169 18751
rect 27203 18748 27215 18751
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 27203 18720 27629 18748
rect 27203 18717 27215 18720
rect 27157 18711 27215 18717
rect 27617 18717 27629 18720
rect 27663 18748 27675 18751
rect 28902 18748 28908 18760
rect 27663 18720 28908 18748
rect 27663 18717 27675 18720
rect 27617 18711 27675 18717
rect 28902 18708 28908 18720
rect 28960 18708 28966 18760
rect 31570 18748 31576 18760
rect 30024 18720 31576 18748
rect 30024 18680 30052 18720
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 32030 18748 32036 18760
rect 31991 18720 32036 18748
rect 32030 18708 32036 18720
rect 32088 18708 32094 18760
rect 35618 18708 35624 18760
rect 35676 18748 35682 18760
rect 36357 18751 36415 18757
rect 36357 18748 36369 18751
rect 35676 18720 36369 18748
rect 35676 18708 35682 18720
rect 36357 18717 36369 18720
rect 36403 18717 36415 18751
rect 36357 18711 36415 18717
rect 36446 18708 36452 18760
rect 36504 18748 36510 18760
rect 36613 18751 36671 18757
rect 36613 18748 36625 18751
rect 36504 18720 36625 18748
rect 36504 18708 36510 18720
rect 36613 18717 36625 18720
rect 36659 18717 36671 18751
rect 36613 18711 36671 18717
rect 25792 18652 30052 18680
rect 31205 18683 31263 18689
rect 31205 18649 31217 18683
rect 31251 18680 31263 18683
rect 31294 18680 31300 18692
rect 31251 18652 31300 18680
rect 31251 18649 31263 18652
rect 31205 18643 31263 18649
rect 31294 18640 31300 18652
rect 31352 18680 31358 18692
rect 31662 18680 31668 18692
rect 31352 18652 31668 18680
rect 31352 18640 31358 18652
rect 31662 18640 31668 18652
rect 31720 18680 31726 18692
rect 32677 18683 32735 18689
rect 32677 18680 32689 18683
rect 31720 18652 32689 18680
rect 31720 18640 31726 18652
rect 32677 18649 32689 18652
rect 32723 18649 32735 18683
rect 32677 18643 32735 18649
rect 22278 18612 22284 18624
rect 21560 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22465 18615 22523 18621
rect 22465 18581 22477 18615
rect 22511 18612 22523 18615
rect 24762 18612 24768 18624
rect 22511 18584 24768 18612
rect 22511 18581 22523 18584
rect 22465 18575 22523 18581
rect 24762 18572 24768 18584
rect 24820 18572 24826 18624
rect 30006 18572 30012 18624
rect 30064 18612 30070 18624
rect 30377 18615 30435 18621
rect 30377 18612 30389 18615
rect 30064 18584 30389 18612
rect 30064 18572 30070 18584
rect 30377 18581 30389 18584
rect 30423 18612 30435 18615
rect 31113 18615 31171 18621
rect 31113 18612 31125 18615
rect 30423 18584 31125 18612
rect 30423 18581 30435 18584
rect 30377 18575 30435 18581
rect 31113 18581 31125 18584
rect 31159 18581 31171 18615
rect 31113 18575 31171 18581
rect 32217 18615 32275 18621
rect 32217 18581 32229 18615
rect 32263 18612 32275 18615
rect 32306 18612 32312 18624
rect 32263 18584 32312 18612
rect 32263 18581 32275 18584
rect 32217 18575 32275 18581
rect 32306 18572 32312 18584
rect 32364 18572 32370 18624
rect 33594 18572 33600 18624
rect 33652 18612 33658 18624
rect 34977 18615 35035 18621
rect 34977 18612 34989 18615
rect 33652 18584 34989 18612
rect 33652 18572 33658 18584
rect 34977 18581 34989 18584
rect 35023 18581 35035 18615
rect 34977 18575 35035 18581
rect 35069 18615 35127 18621
rect 35069 18581 35081 18615
rect 35115 18612 35127 18615
rect 35802 18612 35808 18624
rect 35115 18584 35808 18612
rect 35115 18581 35127 18584
rect 35069 18575 35127 18581
rect 35802 18572 35808 18584
rect 35860 18572 35866 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 5721 18411 5779 18417
rect 5721 18408 5733 18411
rect 5684 18380 5733 18408
rect 5684 18368 5690 18380
rect 5721 18377 5733 18380
rect 5767 18377 5779 18411
rect 5721 18371 5779 18377
rect 7101 18411 7159 18417
rect 7101 18377 7113 18411
rect 7147 18408 7159 18411
rect 7282 18408 7288 18420
rect 7147 18380 7288 18408
rect 7147 18377 7159 18380
rect 7101 18371 7159 18377
rect 5736 18272 5764 18371
rect 7282 18368 7288 18380
rect 7340 18368 7346 18420
rect 11974 18408 11980 18420
rect 11935 18380 11980 18408
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 17589 18411 17647 18417
rect 17589 18408 17601 18411
rect 12084 18380 17601 18408
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 5736 18244 6377 18272
rect 6365 18241 6377 18244
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 6822 18232 6828 18284
rect 6880 18272 6886 18284
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 6880 18244 7205 18272
rect 6880 18232 6886 18244
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7300 18272 7328 18368
rect 9766 18300 9772 18352
rect 9824 18340 9830 18352
rect 12084 18340 12112 18380
rect 17589 18377 17601 18380
rect 17635 18408 17647 18411
rect 18782 18408 18788 18420
rect 17635 18380 18788 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 18248 18349 18276 18380
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 23293 18411 23351 18417
rect 22152 18380 22197 18408
rect 22152 18368 22158 18380
rect 23293 18377 23305 18411
rect 23339 18408 23351 18411
rect 24394 18408 24400 18420
rect 23339 18380 24400 18408
rect 23339 18377 23351 18380
rect 23293 18371 23351 18377
rect 24394 18368 24400 18380
rect 24452 18368 24458 18420
rect 26326 18408 26332 18420
rect 26287 18380 26332 18408
rect 26326 18368 26332 18380
rect 26384 18368 26390 18420
rect 27430 18408 27436 18420
rect 27391 18380 27436 18408
rect 27430 18368 27436 18380
rect 27488 18408 27494 18420
rect 27706 18408 27712 18420
rect 27488 18380 27712 18408
rect 27488 18368 27494 18380
rect 27706 18368 27712 18380
rect 27764 18408 27770 18420
rect 28261 18411 28319 18417
rect 28261 18408 28273 18411
rect 27764 18380 28273 18408
rect 27764 18368 27770 18380
rect 28261 18377 28273 18380
rect 28307 18377 28319 18411
rect 28261 18371 28319 18377
rect 29086 18368 29092 18420
rect 29144 18408 29150 18420
rect 33594 18408 33600 18420
rect 29144 18380 33600 18408
rect 29144 18368 29150 18380
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 35894 18368 35900 18420
rect 35952 18408 35958 18420
rect 35989 18411 36047 18417
rect 35989 18408 36001 18411
rect 35952 18380 36001 18408
rect 35952 18368 35958 18380
rect 35989 18377 36001 18380
rect 36035 18377 36047 18411
rect 35989 18371 36047 18377
rect 36725 18411 36783 18417
rect 36725 18377 36737 18411
rect 36771 18408 36783 18411
rect 37826 18408 37832 18420
rect 36771 18380 37832 18408
rect 36771 18377 36783 18380
rect 36725 18371 36783 18377
rect 37826 18368 37832 18380
rect 37884 18368 37890 18420
rect 18233 18343 18291 18349
rect 9824 18312 12112 18340
rect 13740 18312 14688 18340
rect 9824 18300 9830 18312
rect 7745 18275 7803 18281
rect 7745 18272 7757 18275
rect 7300 18244 7757 18272
rect 7193 18235 7251 18241
rect 7745 18241 7757 18244
rect 7791 18241 7803 18275
rect 8386 18272 8392 18284
rect 8347 18244 8392 18272
rect 7745 18235 7803 18241
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18272 12219 18275
rect 12894 18272 12900 18284
rect 12207 18244 12900 18272
rect 12207 18241 12219 18244
rect 12161 18235 12219 18241
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 13740 18281 13768 18312
rect 13725 18275 13783 18281
rect 13725 18241 13737 18275
rect 13771 18241 13783 18275
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13725 18235 13783 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14660 18281 14688 18312
rect 18233 18309 18245 18343
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 18417 18343 18475 18349
rect 18417 18309 18429 18343
rect 18463 18340 18475 18343
rect 18506 18340 18512 18352
rect 18463 18312 18512 18340
rect 18463 18309 18475 18312
rect 18417 18303 18475 18309
rect 18506 18300 18512 18312
rect 18564 18340 18570 18352
rect 19150 18340 19156 18352
rect 18564 18312 19156 18340
rect 18564 18300 18570 18312
rect 19150 18300 19156 18312
rect 19208 18300 19214 18352
rect 19978 18300 19984 18352
rect 20036 18340 20042 18352
rect 22830 18340 22836 18352
rect 20036 18312 22692 18340
rect 22791 18312 22836 18340
rect 20036 18300 20042 18312
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18272 14703 18275
rect 14826 18272 14832 18284
rect 14691 18244 14832 18272
rect 14691 18241 14703 18244
rect 14645 18235 14703 18241
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 15010 18272 15016 18284
rect 14967 18244 15016 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 21913 18275 21971 18281
rect 21913 18241 21925 18275
rect 21959 18272 21971 18275
rect 22002 18272 22008 18284
rect 21959 18244 22008 18272
rect 21959 18241 21971 18244
rect 21913 18235 21971 18241
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 3510 18164 3516 18216
rect 3568 18204 3574 18216
rect 9674 18204 9680 18216
rect 3568 18176 9680 18204
rect 3568 18164 3574 18176
rect 9674 18164 9680 18176
rect 9732 18204 9738 18216
rect 11882 18204 11888 18216
rect 9732 18176 11888 18204
rect 9732 18164 9738 18176
rect 11882 18164 11888 18176
rect 11940 18204 11946 18216
rect 12250 18204 12256 18216
rect 11940 18176 12256 18204
rect 11940 18164 11946 18176
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 13906 18204 13912 18216
rect 13867 18176 13912 18204
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 15194 18204 15200 18216
rect 14783 18176 15200 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 15194 18164 15200 18176
rect 15252 18164 15258 18216
rect 8573 18139 8631 18145
rect 8573 18105 8585 18139
rect 8619 18136 8631 18139
rect 9122 18136 9128 18148
rect 8619 18108 9128 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 22664 18136 22692 18312
rect 22830 18300 22836 18312
rect 22888 18340 22894 18352
rect 23753 18343 23811 18349
rect 23753 18340 23765 18343
rect 22888 18312 23765 18340
rect 22888 18300 22894 18312
rect 23753 18309 23765 18312
rect 23799 18309 23811 18343
rect 23753 18303 23811 18309
rect 23014 18272 23020 18284
rect 22975 18244 23020 18272
rect 23014 18232 23020 18244
rect 23072 18232 23078 18284
rect 23106 18232 23112 18284
rect 23164 18272 23170 18284
rect 24762 18272 24768 18284
rect 23164 18244 23209 18272
rect 24723 18244 24768 18272
rect 23164 18232 23170 18244
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 26344 18272 26372 18368
rect 34514 18340 34520 18352
rect 32232 18312 34520 18340
rect 27798 18272 27804 18284
rect 26344 18244 27804 18272
rect 25041 18207 25099 18213
rect 25041 18173 25053 18207
rect 25087 18204 25099 18207
rect 26510 18204 26516 18216
rect 25087 18176 26516 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 26510 18164 26516 18176
rect 26568 18164 26574 18216
rect 27172 18213 27200 18244
rect 27798 18232 27804 18244
rect 27856 18232 27862 18284
rect 32232 18281 32260 18312
rect 34514 18300 34520 18312
rect 34572 18340 34578 18352
rect 35618 18340 35624 18352
rect 34572 18312 35624 18340
rect 34572 18300 34578 18312
rect 35618 18300 35624 18312
rect 35676 18300 35682 18352
rect 32217 18275 32275 18281
rect 32217 18241 32229 18275
rect 32263 18241 32275 18275
rect 32217 18235 32275 18241
rect 32306 18232 32312 18284
rect 32364 18272 32370 18284
rect 32473 18275 32531 18281
rect 32473 18272 32485 18275
rect 32364 18244 32485 18272
rect 32364 18232 32370 18244
rect 32473 18241 32485 18244
rect 32519 18241 32531 18275
rect 32473 18235 32531 18241
rect 34698 18232 34704 18284
rect 34756 18272 34762 18284
rect 35342 18272 35348 18284
rect 34756 18244 35348 18272
rect 34756 18232 34762 18244
rect 35342 18232 35348 18244
rect 35400 18232 35406 18284
rect 35529 18275 35587 18281
rect 35529 18241 35541 18275
rect 35575 18272 35587 18275
rect 35710 18272 35716 18284
rect 35575 18244 35716 18272
rect 35575 18241 35587 18244
rect 35529 18235 35587 18241
rect 35710 18232 35716 18244
rect 35768 18232 35774 18284
rect 36538 18272 36544 18284
rect 36499 18244 36544 18272
rect 36538 18232 36544 18244
rect 36596 18232 36602 18284
rect 37274 18232 37280 18284
rect 37332 18272 37338 18284
rect 37829 18275 37887 18281
rect 37829 18272 37841 18275
rect 37332 18244 37841 18272
rect 37332 18232 37338 18244
rect 37829 18241 37841 18244
rect 37875 18241 37887 18275
rect 37829 18235 37887 18241
rect 27157 18207 27215 18213
rect 27157 18173 27169 18207
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 27341 18207 27399 18213
rect 27341 18173 27353 18207
rect 27387 18204 27399 18207
rect 27522 18204 27528 18216
rect 27387 18176 27528 18204
rect 27387 18173 27399 18176
rect 27341 18167 27399 18173
rect 27522 18164 27528 18176
rect 27580 18164 27586 18216
rect 35621 18207 35679 18213
rect 35621 18173 35633 18207
rect 35667 18204 35679 18207
rect 35802 18204 35808 18216
rect 35667 18176 35808 18204
rect 35667 18173 35679 18176
rect 35621 18167 35679 18173
rect 35802 18164 35808 18176
rect 35860 18164 35866 18216
rect 29362 18136 29368 18148
rect 13832 18108 14688 18136
rect 22664 18108 29368 18136
rect 13832 18080 13860 18108
rect 14660 18080 14688 18108
rect 29362 18096 29368 18108
rect 29420 18096 29426 18148
rect 4706 18068 4712 18080
rect 4619 18040 4712 18068
rect 4706 18028 4712 18040
rect 4764 18068 4770 18080
rect 5350 18068 5356 18080
rect 4764 18040 5356 18068
rect 4764 18028 4770 18040
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 6546 18068 6552 18080
rect 6507 18040 6552 18068
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 7926 18068 7932 18080
rect 7887 18040 7932 18068
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8996 18040 9045 18068
rect 8996 18028 9002 18040
rect 9033 18037 9045 18040
rect 9079 18037 9091 18071
rect 9033 18031 9091 18037
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13541 18071 13599 18077
rect 13541 18068 13553 18071
rect 13412 18040 13553 18068
rect 13412 18028 13418 18040
rect 13541 18037 13553 18040
rect 13587 18037 13599 18071
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13541 18031 13599 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14458 18068 14464 18080
rect 14419 18040 14464 18068
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 14642 18028 14648 18080
rect 14700 18068 14706 18080
rect 22922 18068 22928 18080
rect 14700 18040 14793 18068
rect 22883 18040 22928 18068
rect 14700 18028 14706 18040
rect 22922 18028 22928 18040
rect 22980 18028 22986 18080
rect 27798 18068 27804 18080
rect 27759 18040 27804 18068
rect 27798 18028 27804 18040
rect 27856 18028 27862 18080
rect 35342 18068 35348 18080
rect 35303 18040 35348 18068
rect 35342 18028 35348 18040
rect 35400 18028 35406 18080
rect 37274 18068 37280 18080
rect 37235 18040 37280 18068
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 38010 18068 38016 18080
rect 37971 18040 38016 18068
rect 38010 18028 38016 18040
rect 38068 18028 38074 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 8386 17864 8392 17876
rect 7975 17836 8392 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 14642 17864 14648 17876
rect 14603 17836 14648 17864
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 21821 17867 21879 17873
rect 21821 17833 21833 17867
rect 21867 17864 21879 17867
rect 22002 17864 22008 17876
rect 21867 17836 22008 17864
rect 21867 17833 21879 17836
rect 21821 17827 21879 17833
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 22922 17864 22928 17876
rect 22883 17836 22928 17864
rect 22922 17824 22928 17836
rect 22980 17824 22986 17876
rect 29270 17824 29276 17876
rect 29328 17864 29334 17876
rect 29549 17867 29607 17873
rect 29549 17864 29561 17867
rect 29328 17836 29561 17864
rect 29328 17824 29334 17836
rect 29549 17833 29561 17836
rect 29595 17833 29607 17867
rect 29549 17827 29607 17833
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 2590 17796 2596 17808
rect 1627 17768 2596 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 2590 17756 2596 17768
rect 2648 17756 2654 17808
rect 18325 17799 18383 17805
rect 18325 17765 18337 17799
rect 18371 17796 18383 17799
rect 18414 17796 18420 17808
rect 18371 17768 18420 17796
rect 18371 17765 18383 17768
rect 18325 17759 18383 17765
rect 18414 17756 18420 17768
rect 18472 17796 18478 17808
rect 18782 17796 18788 17808
rect 18472 17768 18788 17796
rect 18472 17756 18478 17768
rect 18782 17756 18788 17768
rect 18840 17756 18846 17808
rect 23014 17796 23020 17808
rect 22940 17768 23020 17796
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 7561 17731 7619 17737
rect 7561 17728 7573 17731
rect 6604 17700 7573 17728
rect 6604 17688 6610 17700
rect 7561 17697 7573 17700
rect 7607 17697 7619 17731
rect 8938 17728 8944 17740
rect 8899 17700 8944 17728
rect 7561 17691 7619 17697
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9122 17728 9128 17740
rect 9083 17700 9128 17728
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 9674 17728 9680 17740
rect 9635 17700 9680 17728
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17728 14795 17731
rect 15194 17728 15200 17740
rect 14783 17700 15200 17728
rect 14783 17697 14795 17700
rect 14737 17691 14795 17697
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 22940 17737 22968 17768
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 22925 17731 22983 17737
rect 22925 17697 22937 17731
rect 22971 17697 22983 17731
rect 26510 17728 26516 17740
rect 26471 17700 26516 17728
rect 22925 17691 22983 17697
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 27706 17728 27712 17740
rect 27667 17700 27712 17728
rect 27706 17688 27712 17700
rect 27764 17688 27770 17740
rect 30098 17728 30104 17740
rect 30059 17700 30104 17728
rect 30098 17688 30104 17700
rect 30156 17688 30162 17740
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17660 1458 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 1452 17632 2053 17660
rect 1452 17620 1458 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 7926 17660 7932 17672
rect 7791 17632 7932 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 12342 17660 12348 17672
rect 12303 17632 12348 17660
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 13354 17660 13360 17672
rect 13315 17632 13360 17660
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 14921 17663 14979 17669
rect 14921 17660 14933 17663
rect 14884 17632 14933 17660
rect 14884 17620 14890 17632
rect 14921 17629 14933 17632
rect 14967 17629 14979 17663
rect 17586 17660 17592 17672
rect 17499 17632 17592 17660
rect 14921 17623 14979 17629
rect 17586 17620 17592 17632
rect 17644 17660 17650 17672
rect 22741 17663 22799 17669
rect 17644 17632 18184 17660
rect 17644 17620 17650 17632
rect 7374 17552 7380 17604
rect 7432 17592 7438 17604
rect 7469 17595 7527 17601
rect 7469 17592 7481 17595
rect 7432 17564 7481 17592
rect 7432 17552 7438 17564
rect 7469 17561 7481 17564
rect 7515 17561 7527 17595
rect 7469 17555 7527 17561
rect 13998 17552 14004 17604
rect 14056 17592 14062 17604
rect 14645 17595 14703 17601
rect 14645 17592 14657 17595
rect 14056 17564 14657 17592
rect 14056 17552 14062 17564
rect 14645 17561 14657 17564
rect 14691 17592 14703 17595
rect 15010 17592 15016 17604
rect 14691 17564 15016 17592
rect 14691 17561 14703 17564
rect 14645 17555 14703 17561
rect 15010 17552 15016 17564
rect 15068 17592 15074 17604
rect 18156 17601 18184 17632
rect 22741 17629 22753 17663
rect 22787 17660 22799 17663
rect 22830 17660 22836 17672
rect 22787 17632 22836 17660
rect 22787 17629 22799 17632
rect 22741 17623 22799 17629
rect 22830 17620 22836 17632
rect 22888 17620 22894 17672
rect 23017 17663 23075 17669
rect 23017 17629 23029 17663
rect 23063 17660 23075 17663
rect 23106 17660 23112 17672
rect 23063 17632 23112 17660
rect 23063 17629 23075 17632
rect 23017 17623 23075 17629
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 26329 17663 26387 17669
rect 26329 17629 26341 17663
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 18141 17595 18199 17601
rect 15068 17564 17632 17592
rect 15068 17552 15074 17564
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 6917 17527 6975 17533
rect 6917 17524 6929 17527
rect 6880 17496 6929 17524
rect 6880 17484 6886 17496
rect 6917 17493 6929 17496
rect 6963 17524 6975 17527
rect 10134 17524 10140 17536
rect 6963 17496 10140 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 13173 17527 13231 17533
rect 13173 17524 13185 17527
rect 12584 17496 13185 17524
rect 12584 17484 12590 17496
rect 13173 17493 13185 17496
rect 13219 17493 13231 17527
rect 13173 17487 13231 17493
rect 15105 17527 15163 17533
rect 15105 17493 15117 17527
rect 15151 17524 15163 17527
rect 15562 17524 15568 17536
rect 15151 17496 15568 17524
rect 15151 17493 15163 17496
rect 15105 17487 15163 17493
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 17604 17524 17632 17564
rect 18141 17561 18153 17595
rect 18187 17592 18199 17595
rect 20162 17592 20168 17604
rect 18187 17564 20168 17592
rect 18187 17561 18199 17564
rect 18141 17555 18199 17561
rect 20162 17552 20168 17564
rect 20220 17552 20226 17604
rect 26344 17592 26372 17623
rect 27798 17620 27804 17672
rect 27856 17660 27862 17672
rect 28629 17663 28687 17669
rect 28629 17660 28641 17663
rect 27856 17632 28641 17660
rect 27856 17620 27862 17632
rect 28629 17629 28641 17632
rect 28675 17629 28687 17663
rect 28629 17623 28687 17629
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 29270 17660 29276 17672
rect 28868 17632 29276 17660
rect 28868 17620 28874 17632
rect 29270 17620 29276 17632
rect 29328 17620 29334 17672
rect 27522 17592 27528 17604
rect 26344 17564 27528 17592
rect 27522 17552 27528 17564
rect 27580 17552 27586 17604
rect 30282 17592 30288 17604
rect 30243 17564 30288 17592
rect 30282 17552 30288 17564
rect 30340 17552 30346 17604
rect 31662 17552 31668 17604
rect 31720 17592 31726 17604
rect 31941 17595 31999 17601
rect 31941 17592 31953 17595
rect 31720 17564 31953 17592
rect 31720 17552 31726 17564
rect 31941 17561 31953 17564
rect 31987 17592 31999 17595
rect 34514 17592 34520 17604
rect 31987 17564 34520 17592
rect 31987 17561 31999 17564
rect 31941 17555 31999 17561
rect 34514 17552 34520 17564
rect 34572 17552 34578 17604
rect 20714 17524 20720 17536
rect 17604 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 23201 17527 23259 17533
rect 23201 17493 23213 17527
rect 23247 17524 23259 17527
rect 23750 17524 23756 17536
rect 23247 17496 23756 17524
rect 23247 17493 23259 17496
rect 23201 17487 23259 17493
rect 23750 17484 23756 17496
rect 23808 17484 23814 17536
rect 27614 17484 27620 17536
rect 27672 17524 27678 17536
rect 28997 17527 29055 17533
rect 28997 17524 29009 17527
rect 27672 17496 29009 17524
rect 27672 17484 27678 17496
rect 28997 17493 29009 17496
rect 29043 17493 29055 17527
rect 28997 17487 29055 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 7374 17320 7380 17332
rect 6696 17292 7380 17320
rect 6696 17280 6702 17292
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 4890 17252 4896 17264
rect 4663 17224 4896 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 4890 17212 4896 17224
rect 4948 17212 4954 17264
rect 6840 17261 6868 17292
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 7800 17292 8769 17320
rect 7800 17280 7806 17292
rect 8757 17289 8769 17292
rect 8803 17320 8815 17323
rect 9030 17320 9036 17332
rect 8803 17292 9036 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 17586 17320 17592 17332
rect 10192 17292 17592 17320
rect 10192 17280 10198 17292
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 22830 17320 22836 17332
rect 22695 17292 22836 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 30101 17323 30159 17329
rect 30101 17289 30113 17323
rect 30147 17320 30159 17323
rect 36538 17320 36544 17332
rect 30147 17292 36544 17320
rect 30147 17289 30159 17292
rect 30101 17283 30159 17289
rect 36538 17280 36544 17292
rect 36596 17280 36602 17332
rect 6825 17255 6883 17261
rect 6825 17221 6837 17255
rect 6871 17252 6883 17255
rect 12526 17252 12532 17264
rect 6871 17224 6905 17252
rect 7116 17224 7972 17252
rect 12487 17224 12532 17252
rect 6871 17221 6883 17224
rect 6825 17215 6883 17221
rect 7116 17193 7144 17224
rect 7944 17196 7972 17224
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 28813 17255 28871 17261
rect 28813 17252 28825 17255
rect 26988 17224 28825 17252
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7558 17144 7564 17196
rect 7616 17184 7622 17196
rect 7742 17184 7748 17196
rect 7616 17156 7748 17184
rect 7616 17144 7622 17156
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7984 17156 8033 17184
rect 7984 17144 7990 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 12342 17184 12348 17196
rect 12303 17156 12348 17184
rect 8021 17147 8079 17153
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 23750 17184 23756 17196
rect 23711 17156 23756 17184
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 26988 17193 27016 17224
rect 28813 17221 28825 17224
rect 28859 17252 28871 17255
rect 28994 17252 29000 17264
rect 28859 17224 29000 17252
rect 28859 17221 28871 17224
rect 28813 17215 28871 17221
rect 28994 17212 29000 17224
rect 29052 17212 29058 17264
rect 27246 17193 27252 17196
rect 26973 17187 27031 17193
rect 26973 17153 26985 17187
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27240 17147 27252 17193
rect 27304 17184 27310 17196
rect 27304 17156 27340 17184
rect 27246 17144 27252 17147
rect 27304 17144 27310 17156
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 34609 17187 34667 17193
rect 27580 17156 28396 17184
rect 27580 17144 27586 17156
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 2958 17116 2964 17128
rect 2919 17088 2964 17116
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 7009 17119 7067 17125
rect 7009 17116 7021 17119
rect 6604 17088 7021 17116
rect 6604 17076 6610 17088
rect 7009 17085 7021 17088
rect 7055 17116 7067 17119
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7055 17088 7849 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7837 17085 7849 17088
rect 7883 17085 7895 17119
rect 13998 17116 14004 17128
rect 13959 17088 14004 17116
rect 7837 17079 7895 17085
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 17770 17116 17776 17128
rect 17731 17088 17776 17116
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 17954 17116 17960 17128
rect 17915 17088 17960 17116
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 19334 17116 19340 17128
rect 19295 17088 19340 17116
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 26142 17116 26148 17128
rect 24075 17088 26148 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 26142 17076 26148 17088
rect 26200 17076 26206 17128
rect 7466 17048 7472 17060
rect 7116 17020 7472 17048
rect 7116 16989 7144 17020
rect 7466 17008 7472 17020
rect 7524 17048 7530 17060
rect 28368 17057 28396 17156
rect 34609 17153 34621 17187
rect 34655 17184 34667 17187
rect 34698 17184 34704 17196
rect 34655 17156 34704 17184
rect 34655 17153 34667 17156
rect 34609 17147 34667 17153
rect 34698 17144 34704 17156
rect 34756 17184 34762 17196
rect 35069 17187 35127 17193
rect 35069 17184 35081 17187
rect 34756 17156 35081 17184
rect 34756 17144 34762 17156
rect 35069 17153 35081 17156
rect 35115 17153 35127 17187
rect 35069 17147 35127 17153
rect 35232 17190 35290 17196
rect 35232 17156 35244 17190
rect 35278 17156 35290 17190
rect 35348 17190 35406 17196
rect 35348 17184 35360 17190
rect 35232 17150 35290 17156
rect 35347 17156 35360 17184
rect 35394 17156 35406 17190
rect 35347 17150 35406 17156
rect 35437 17187 35495 17193
rect 35437 17153 35449 17187
rect 35483 17153 35495 17187
rect 29362 17076 29368 17128
rect 29420 17116 29426 17128
rect 29641 17119 29699 17125
rect 29641 17116 29653 17119
rect 29420 17088 29653 17116
rect 29420 17076 29426 17088
rect 29641 17085 29653 17088
rect 29687 17085 29699 17119
rect 29641 17079 29699 17085
rect 34790 17076 34796 17128
rect 34848 17116 34854 17128
rect 35247 17116 35275 17150
rect 34848 17088 35275 17116
rect 34848 17076 34854 17088
rect 35347 17060 35375 17150
rect 35437 17147 35495 17153
rect 35452 17116 35480 17147
rect 35526 17116 35532 17128
rect 35452 17088 35532 17116
rect 35526 17076 35532 17088
rect 35584 17076 35590 17128
rect 28353 17051 28411 17057
rect 7524 17020 7788 17048
rect 7524 17008 7530 17020
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16949 7159 16983
rect 7101 16943 7159 16949
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7650 16980 7656 16992
rect 7331 16952 7656 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 7760 16989 7788 17020
rect 28353 17017 28365 17051
rect 28399 17048 28411 17051
rect 29917 17051 29975 17057
rect 29917 17048 29929 17051
rect 28399 17020 29929 17048
rect 28399 17017 28411 17020
rect 28353 17011 28411 17017
rect 29917 17017 29929 17020
rect 29963 17017 29975 17051
rect 29917 17011 29975 17017
rect 35342 17008 35348 17060
rect 35400 17008 35406 17060
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16949 7803 16983
rect 7745 16943 7803 16949
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8570 16980 8576 16992
rect 8251 16952 8576 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 20162 16980 20168 16992
rect 19392 16952 20168 16980
rect 19392 16940 19398 16952
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 35713 16983 35771 16989
rect 35713 16949 35725 16983
rect 35759 16980 35771 16983
rect 35894 16980 35900 16992
rect 35759 16952 35900 16980
rect 35759 16949 35771 16952
rect 35713 16943 35771 16949
rect 35894 16940 35900 16952
rect 35952 16940 35958 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2832 16748 2881 16776
rect 2832 16736 2838 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 2869 16739 2927 16745
rect 6917 16779 6975 16785
rect 6917 16745 6929 16779
rect 6963 16776 6975 16779
rect 7466 16776 7472 16788
rect 6963 16748 7472 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7466 16736 7472 16748
rect 7524 16776 7530 16788
rect 7561 16779 7619 16785
rect 7561 16776 7573 16779
rect 7524 16748 7573 16776
rect 7524 16736 7530 16748
rect 7561 16745 7573 16748
rect 7607 16745 7619 16779
rect 9030 16776 9036 16788
rect 8991 16748 9036 16776
rect 7561 16739 7619 16745
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 17828 16748 17877 16776
rect 17828 16736 17834 16748
rect 17865 16745 17877 16748
rect 17911 16745 17923 16779
rect 17865 16739 17923 16745
rect 27246 16736 27252 16788
rect 27304 16776 27310 16788
rect 27341 16779 27399 16785
rect 27341 16776 27353 16779
rect 27304 16748 27353 16776
rect 27304 16736 27310 16748
rect 27341 16745 27353 16748
rect 27387 16745 27399 16779
rect 27341 16739 27399 16745
rect 3418 16668 3424 16720
rect 3476 16708 3482 16720
rect 8294 16708 8300 16720
rect 3476 16680 8300 16708
rect 3476 16668 3482 16680
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6604 16612 6745 16640
rect 6604 16600 6610 16612
rect 6733 16609 6745 16612
rect 6779 16640 6791 16643
rect 7653 16643 7711 16649
rect 7653 16640 7665 16643
rect 6779 16612 7665 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 7653 16609 7665 16612
rect 7699 16609 7711 16643
rect 7653 16603 7711 16609
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13906 16640 13912 16652
rect 13587 16612 13912 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 26053 16643 26111 16649
rect 26053 16640 26065 16643
rect 23808 16612 26065 16640
rect 23808 16600 23814 16612
rect 26053 16609 26065 16612
rect 26099 16609 26111 16643
rect 26053 16603 26111 16609
rect 26329 16643 26387 16649
rect 26329 16609 26341 16643
rect 26375 16640 26387 16643
rect 30282 16640 30288 16652
rect 26375 16612 30288 16640
rect 26375 16609 26387 16612
rect 26329 16603 26387 16609
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 35618 16640 35624 16652
rect 35579 16612 35624 16640
rect 35618 16600 35624 16612
rect 35676 16600 35682 16652
rect 3786 16572 3792 16584
rect 3747 16544 3792 16572
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 6638 16572 6644 16584
rect 6599 16544 6644 16572
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16541 6975 16575
rect 7558 16572 7564 16584
rect 7519 16544 7564 16572
rect 6917 16535 6975 16541
rect 6932 16504 6960 16535
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16572 7895 16575
rect 7926 16572 7932 16584
rect 7883 16544 7932 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 7852 16504 7880 16535
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 14645 16575 14703 16581
rect 14645 16572 14657 16575
rect 14516 16544 14657 16572
rect 14516 16532 14522 16544
rect 14645 16541 14657 16544
rect 14691 16541 14703 16575
rect 15562 16572 15568 16584
rect 15523 16544 15568 16572
rect 14645 16535 14703 16541
rect 15562 16532 15568 16544
rect 15620 16532 15626 16584
rect 27525 16575 27583 16581
rect 27525 16541 27537 16575
rect 27571 16572 27583 16575
rect 27614 16572 27620 16584
rect 27571 16544 27620 16572
rect 27571 16541 27583 16544
rect 27525 16535 27583 16541
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 35894 16581 35900 16584
rect 35888 16572 35900 16581
rect 35855 16544 35900 16572
rect 35888 16535 35900 16544
rect 35894 16532 35900 16535
rect 35952 16532 35958 16584
rect 6932 16476 7880 16504
rect 7098 16436 7104 16448
rect 7059 16408 7104 16436
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 14090 16396 14096 16448
rect 14148 16436 14154 16448
rect 14461 16439 14519 16445
rect 14461 16436 14473 16439
rect 14148 16408 14473 16436
rect 14148 16396 14154 16408
rect 14461 16405 14473 16408
rect 14507 16405 14519 16439
rect 14461 16399 14519 16405
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15712 16408 15761 16436
rect 15712 16396 15718 16408
rect 15749 16405 15761 16408
rect 15795 16405 15807 16439
rect 20162 16436 20168 16448
rect 20123 16408 20168 16436
rect 15749 16399 15807 16405
rect 20162 16396 20168 16408
rect 20220 16396 20226 16448
rect 35802 16396 35808 16448
rect 35860 16436 35866 16448
rect 37001 16439 37059 16445
rect 37001 16436 37013 16439
rect 35860 16408 37013 16436
rect 35860 16396 35866 16408
rect 37001 16405 37013 16408
rect 37047 16405 37059 16439
rect 37001 16399 37059 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2869 16235 2927 16241
rect 2869 16201 2881 16235
rect 2915 16232 2927 16235
rect 2958 16232 2964 16244
rect 2915 16204 2964 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3329 16235 3387 16241
rect 3329 16201 3341 16235
rect 3375 16201 3387 16235
rect 3329 16195 3387 16201
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 17954 16232 17960 16244
rect 17911 16204 17960 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16096 1458 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1452 16068 2053 16096
rect 1452 16056 1458 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 3344 16096 3372 16195
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 18969 16235 19027 16241
rect 18969 16201 18981 16235
rect 19015 16232 19027 16235
rect 19242 16232 19248 16244
rect 19015 16204 19248 16232
rect 19015 16201 19027 16204
rect 18969 16195 19027 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 22833 16235 22891 16241
rect 22833 16201 22845 16235
rect 22879 16232 22891 16235
rect 23566 16232 23572 16244
rect 22879 16204 23572 16232
rect 22879 16201 22891 16204
rect 22833 16195 22891 16201
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 23750 16232 23756 16244
rect 23711 16204 23756 16232
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 30745 16235 30803 16241
rect 30745 16201 30757 16235
rect 30791 16232 30803 16235
rect 31202 16232 31208 16244
rect 30791 16204 31208 16232
rect 30791 16201 30803 16204
rect 30745 16195 30803 16201
rect 31202 16192 31208 16204
rect 31260 16232 31266 16244
rect 31570 16232 31576 16244
rect 31260 16204 31576 16232
rect 31260 16192 31266 16204
rect 31570 16192 31576 16204
rect 31628 16192 31634 16244
rect 3789 16167 3847 16173
rect 3789 16133 3801 16167
rect 3835 16164 3847 16167
rect 3878 16164 3884 16176
rect 3835 16136 3884 16164
rect 3835 16133 3847 16136
rect 3789 16127 3847 16133
rect 3878 16124 3884 16136
rect 3936 16124 3942 16176
rect 14090 16164 14096 16176
rect 14051 16136 14096 16164
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 18509 16167 18567 16173
rect 18509 16133 18521 16167
rect 18555 16164 18567 16167
rect 18598 16164 18604 16176
rect 18555 16136 18604 16164
rect 18555 16133 18567 16136
rect 18509 16127 18567 16133
rect 18598 16124 18604 16136
rect 18656 16124 18662 16176
rect 23290 16164 23296 16176
rect 20732 16136 23296 16164
rect 2731 16068 3372 16096
rect 3513 16099 3571 16105
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 3513 16065 3525 16099
rect 3559 16096 3571 16099
rect 3602 16096 3608 16108
rect 3559 16068 3608 16096
rect 3559 16065 3571 16068
rect 3513 16059 3571 16065
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4614 16096 4620 16108
rect 4295 16068 4620 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16065 13139 16099
rect 13906 16096 13912 16108
rect 13867 16068 13912 16096
rect 13081 16059 13139 16065
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 4798 16028 4804 16040
rect 3743 16000 4804 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7653 16031 7711 16037
rect 7653 16028 7665 16031
rect 7248 16000 7665 16028
rect 7248 15988 7254 16000
rect 7653 15997 7665 16000
rect 7699 15997 7711 16031
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7653 15991 7711 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 13096 16028 13124 16059
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18230 16096 18236 16108
rect 18095 16068 18236 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18785 16099 18843 16105
rect 18785 16065 18797 16099
rect 18831 16096 18843 16099
rect 19058 16096 19064 16108
rect 18831 16068 19064 16096
rect 18831 16065 18843 16068
rect 18785 16059 18843 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 20732 16105 20760 16136
rect 23290 16124 23296 16136
rect 23348 16124 23354 16176
rect 26142 16164 26148 16176
rect 26103 16136 26148 16164
rect 26142 16124 26148 16136
rect 26200 16124 26206 16176
rect 35802 16164 35808 16176
rect 33888 16136 35808 16164
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 21821 16099 21879 16105
rect 21821 16096 21833 16099
rect 21048 16068 21833 16096
rect 21048 16056 21054 16068
rect 21821 16065 21833 16068
rect 21867 16065 21879 16099
rect 23474 16096 23480 16108
rect 23435 16068 23480 16096
rect 21821 16059 21879 16065
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 23569 16099 23627 16105
rect 23569 16065 23581 16099
rect 23615 16065 23627 16099
rect 32858 16096 32864 16108
rect 32819 16068 32864 16096
rect 23569 16059 23627 16065
rect 13814 16028 13820 16040
rect 13096 16000 13820 16028
rect 9493 15991 9551 15997
rect 2866 15920 2872 15972
rect 2924 15960 2930 15972
rect 3418 15960 3424 15972
rect 2924 15932 3424 15960
rect 2924 15920 2930 15932
rect 3418 15920 3424 15932
rect 3476 15960 3482 15972
rect 9508 15960 9536 15991
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 16028 15807 16031
rect 15930 16028 15936 16040
rect 15795 16000 15936 16028
rect 15795 15997 15807 16000
rect 15749 15991 15807 15997
rect 15764 15960 15792 15991
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 18506 15988 18512 16040
rect 18564 16028 18570 16040
rect 18601 16031 18659 16037
rect 18601 16028 18613 16031
rect 18564 16000 18613 16028
rect 18564 15988 18570 16000
rect 18601 15997 18613 16000
rect 18647 16028 18659 16031
rect 20441 16031 20499 16037
rect 20441 16028 20453 16031
rect 18647 16000 20453 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 20441 15997 20453 16000
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 23584 16028 23612 16059
rect 32858 16056 32864 16068
rect 32916 16056 32922 16108
rect 33888 16105 33916 16136
rect 35802 16124 35808 16136
rect 35860 16124 35866 16176
rect 33873 16099 33931 16105
rect 33873 16065 33885 16099
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 24670 16028 24676 16040
rect 22612 16000 23612 16028
rect 24631 16000 24676 16028
rect 22612 15988 22618 16000
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 26329 16031 26387 16037
rect 26329 15997 26341 16031
rect 26375 16028 26387 16031
rect 29362 16028 29368 16040
rect 26375 16000 29368 16028
rect 26375 15997 26387 16000
rect 26329 15991 26387 15997
rect 29362 15988 29368 16000
rect 29420 15988 29426 16040
rect 34057 16031 34115 16037
rect 34057 15997 34069 16031
rect 34103 15997 34115 16031
rect 34514 16028 34520 16040
rect 34475 16000 34520 16028
rect 34057 15991 34115 15997
rect 3476 15932 15792 15960
rect 3476 15920 3482 15932
rect 21266 15920 21272 15972
rect 21324 15960 21330 15972
rect 33045 15963 33103 15969
rect 21324 15932 32996 15960
rect 21324 15920 21330 15932
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 3789 15895 3847 15901
rect 3789 15861 3801 15895
rect 3835 15892 3847 15895
rect 4062 15892 4068 15904
rect 3835 15864 4068 15892
rect 3835 15861 3847 15864
rect 3789 15855 3847 15861
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 4706 15892 4712 15904
rect 4479 15864 4712 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 4890 15892 4896 15904
rect 4851 15864 4896 15892
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 11756 15864 12081 15892
rect 11756 15852 11762 15864
rect 12069 15861 12081 15864
rect 12115 15861 12127 15895
rect 12894 15892 12900 15904
rect 12855 15864 12900 15892
rect 12069 15855 12127 15861
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 18690 15892 18696 15904
rect 18651 15864 18696 15892
rect 18690 15852 18696 15864
rect 18748 15852 18754 15904
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 19889 15895 19947 15901
rect 19889 15892 19901 15895
rect 18932 15864 19901 15892
rect 18932 15852 18938 15864
rect 19889 15861 19901 15864
rect 19935 15861 19947 15895
rect 19889 15855 19947 15861
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21784 15864 22017 15892
rect 21784 15852 21790 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 23290 15892 23296 15904
rect 23251 15864 23296 15892
rect 22005 15855 22063 15861
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 29549 15895 29607 15901
rect 29549 15861 29561 15895
rect 29595 15892 29607 15895
rect 30006 15892 30012 15904
rect 29595 15864 30012 15892
rect 29595 15861 29607 15864
rect 29549 15855 29607 15861
rect 30006 15852 30012 15864
rect 30064 15852 30070 15904
rect 31110 15852 31116 15904
rect 31168 15892 31174 15904
rect 32122 15892 32128 15904
rect 31168 15864 32128 15892
rect 31168 15852 31174 15864
rect 32122 15852 32128 15864
rect 32180 15852 32186 15904
rect 32968 15892 32996 15932
rect 33045 15929 33057 15963
rect 33091 15960 33103 15963
rect 34072 15960 34100 15991
rect 34514 15988 34520 16000
rect 34572 15988 34578 16040
rect 33091 15932 34100 15960
rect 33091 15929 33103 15932
rect 33045 15923 33103 15929
rect 34606 15892 34612 15904
rect 32968 15864 34612 15892
rect 34606 15852 34612 15864
rect 34664 15852 34670 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 7190 15688 7196 15700
rect 7151 15660 7196 15688
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7834 15688 7840 15700
rect 7795 15660 7840 15688
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 18230 15688 18236 15700
rect 18191 15660 18236 15688
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18690 15688 18696 15700
rect 18603 15660 18696 15688
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 23385 15691 23443 15697
rect 23385 15657 23397 15691
rect 23431 15657 23443 15691
rect 28994 15688 29000 15700
rect 28955 15660 29000 15688
rect 23385 15651 23443 15657
rect 18708 15620 18736 15648
rect 18708 15592 21404 15620
rect 3786 15552 3792 15564
rect 3747 15524 3792 15552
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 3970 15512 3976 15564
rect 4028 15552 4034 15564
rect 4249 15555 4307 15561
rect 4249 15552 4261 15555
rect 4028 15524 4261 15552
rect 4028 15512 4034 15524
rect 4249 15521 4261 15524
rect 4295 15521 4307 15555
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 4249 15515 4307 15521
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 12894 15552 12900 15564
rect 11931 15524 12900 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13538 15552 13544 15564
rect 13499 15524 13544 15552
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 15654 15552 15660 15564
rect 15615 15524 15660 15552
rect 15654 15512 15660 15524
rect 15712 15512 15718 15564
rect 16666 15552 16672 15564
rect 16627 15524 16672 15552
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 19058 15552 19064 15564
rect 18432 15524 19064 15552
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 7650 15484 7656 15496
rect 7611 15456 7656 15484
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8628 15456 9137 15484
rect 8628 15444 8634 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 11238 15484 11244 15496
rect 11199 15456 11244 15484
rect 9125 15447 9183 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 15470 15484 15476 15496
rect 15431 15456 15476 15484
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 18432 15493 18460 15524
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 19150 15512 19156 15564
rect 19208 15552 19214 15564
rect 19536 15561 19564 15592
rect 21376 15564 21404 15592
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 19208 15524 19257 15552
rect 19208 15512 19214 15524
rect 19245 15521 19257 15524
rect 19291 15521 19303 15555
rect 19245 15515 19303 15521
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15521 19579 15555
rect 21266 15552 21272 15564
rect 21227 15524 21272 15552
rect 19521 15515 19579 15521
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 21358 15512 21364 15564
rect 21416 15552 21422 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21416 15524 22109 15552
rect 21416 15512 21422 15524
rect 22097 15521 22109 15524
rect 22143 15552 22155 15555
rect 23400 15552 23428 15651
rect 28994 15648 29000 15660
rect 29052 15648 29058 15700
rect 32122 15648 32128 15700
rect 32180 15688 32186 15700
rect 32180 15660 34744 15688
rect 32180 15648 32186 15660
rect 32309 15623 32367 15629
rect 32309 15620 32321 15623
rect 23768 15592 32321 15620
rect 23566 15552 23572 15564
rect 22143 15524 23428 15552
rect 23527 15524 23572 15552
rect 22143 15521 22155 15524
rect 22097 15515 22155 15521
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15453 18475 15487
rect 18417 15447 18475 15453
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 18564 15456 18609 15484
rect 18564 15444 18570 15456
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20220 15456 20545 15484
rect 20220 15444 20226 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20806 15484 20812 15496
rect 20767 15456 20812 15484
rect 20625 15447 20683 15453
rect 3973 15419 4031 15425
rect 3973 15385 3985 15419
rect 4019 15385 4031 15419
rect 18690 15416 18696 15428
rect 18651 15388 18696 15416
rect 3973 15379 4031 15385
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15348 3295 15351
rect 3988 15348 4016 15379
rect 18690 15376 18696 15388
rect 18748 15376 18754 15428
rect 18874 15376 18880 15428
rect 18932 15416 18938 15428
rect 20640 15416 20668 15447
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 22370 15484 22376 15496
rect 22283 15456 22376 15484
rect 22370 15444 22376 15456
rect 22428 15484 22434 15496
rect 23290 15484 23296 15496
rect 22428 15456 23296 15484
rect 22428 15444 22434 15456
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 23658 15484 23664 15496
rect 23619 15456 23664 15484
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 18932 15388 20668 15416
rect 23385 15419 23443 15425
rect 18932 15376 18938 15388
rect 23385 15385 23397 15419
rect 23431 15416 23443 15419
rect 23474 15416 23480 15428
rect 23431 15388 23480 15416
rect 23431 15385 23443 15388
rect 23385 15379 23443 15385
rect 23474 15376 23480 15388
rect 23532 15376 23538 15428
rect 23768 15416 23796 15592
rect 32309 15589 32321 15592
rect 32355 15620 32367 15623
rect 34716 15620 34744 15660
rect 34790 15648 34796 15700
rect 34848 15688 34854 15700
rect 34885 15691 34943 15697
rect 34885 15688 34897 15691
rect 34848 15660 34897 15688
rect 34848 15648 34854 15660
rect 34885 15657 34897 15660
rect 34931 15657 34943 15691
rect 37366 15688 37372 15700
rect 34885 15651 34943 15657
rect 35636 15660 37372 15688
rect 35636 15620 35664 15660
rect 37366 15648 37372 15660
rect 37424 15688 37430 15700
rect 37737 15691 37795 15697
rect 37737 15688 37749 15691
rect 37424 15660 37749 15688
rect 37424 15648 37430 15660
rect 37737 15657 37749 15660
rect 37783 15657 37795 15691
rect 37737 15651 37795 15657
rect 32355 15592 32904 15620
rect 34716 15592 35664 15620
rect 32355 15589 32367 15592
rect 32309 15583 32367 15589
rect 24670 15552 24676 15564
rect 24631 15524 24676 15552
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 26513 15555 26571 15561
rect 26513 15521 26525 15555
rect 26559 15552 26571 15555
rect 29086 15552 29092 15564
rect 26559 15524 29092 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 29086 15512 29092 15524
rect 29144 15512 29150 15564
rect 29362 15512 29368 15564
rect 29420 15552 29426 15564
rect 30101 15555 30159 15561
rect 30101 15552 30113 15555
rect 29420 15524 30113 15552
rect 29420 15512 29426 15524
rect 30101 15521 30113 15524
rect 30147 15521 30159 15555
rect 30101 15515 30159 15521
rect 30190 15512 30196 15564
rect 30248 15552 30254 15564
rect 32876 15561 32904 15592
rect 30929 15555 30987 15561
rect 30929 15552 30941 15555
rect 30248 15524 30941 15552
rect 30248 15512 30254 15524
rect 30929 15521 30941 15524
rect 30975 15521 30987 15555
rect 30929 15515 30987 15521
rect 32861 15555 32919 15561
rect 32861 15521 32873 15555
rect 32907 15521 32919 15555
rect 32861 15515 32919 15521
rect 34606 15512 34612 15564
rect 34664 15552 34670 15564
rect 34793 15555 34851 15561
rect 34793 15552 34805 15555
rect 34664 15524 34805 15552
rect 34664 15512 34670 15524
rect 34793 15521 34805 15524
rect 34839 15521 34851 15555
rect 34793 15515 34851 15521
rect 34977 15555 35035 15561
rect 34977 15521 34989 15555
rect 35023 15552 35035 15555
rect 35526 15552 35532 15564
rect 35023 15524 35532 15552
rect 35023 15521 35035 15524
rect 34977 15515 35035 15521
rect 35526 15512 35532 15524
rect 35584 15512 35590 15564
rect 28902 15444 28908 15496
rect 28960 15484 28966 15496
rect 31110 15484 31116 15496
rect 28960 15456 31116 15484
rect 28960 15444 28966 15456
rect 31110 15444 31116 15456
rect 31168 15444 31174 15496
rect 31202 15444 31208 15496
rect 31260 15484 31266 15496
rect 33137 15487 33195 15493
rect 31260 15456 31305 15484
rect 31260 15444 31266 15456
rect 33137 15453 33149 15487
rect 33183 15484 33195 15487
rect 34054 15484 34060 15496
rect 33183 15456 34060 15484
rect 33183 15453 33195 15456
rect 33137 15447 33195 15453
rect 34054 15444 34060 15456
rect 34112 15444 34118 15496
rect 34698 15484 34704 15496
rect 34659 15456 34704 15484
rect 34698 15444 34704 15456
rect 34756 15444 34762 15496
rect 36357 15487 36415 15493
rect 36357 15453 36369 15487
rect 36403 15453 36415 15487
rect 36357 15447 36415 15453
rect 23676 15388 23796 15416
rect 3283 15320 4016 15348
rect 3283 15317 3295 15320
rect 3237 15311 3295 15317
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8720 15320 8953 15348
rect 8720 15308 8726 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 17126 15308 17132 15360
rect 17184 15348 17190 15360
rect 23676 15348 23704 15388
rect 25498 15376 25504 15428
rect 25556 15416 25562 15428
rect 26329 15419 26387 15425
rect 26329 15416 26341 15419
rect 25556 15388 26341 15416
rect 25556 15376 25562 15388
rect 26329 15385 26341 15388
rect 26375 15385 26387 15419
rect 26329 15379 26387 15385
rect 30282 15376 30288 15428
rect 30340 15416 30346 15428
rect 35897 15419 35955 15425
rect 35897 15416 35909 15419
rect 30340 15388 35909 15416
rect 30340 15376 30346 15388
rect 35897 15385 35909 15388
rect 35943 15416 35955 15419
rect 36372 15416 36400 15447
rect 35943 15388 36400 15416
rect 35943 15385 35955 15388
rect 35897 15379 35955 15385
rect 36446 15376 36452 15428
rect 36504 15416 36510 15428
rect 36602 15419 36660 15425
rect 36602 15416 36614 15419
rect 36504 15388 36614 15416
rect 36504 15376 36510 15388
rect 36602 15385 36614 15388
rect 36648 15385 36660 15419
rect 36602 15379 36660 15385
rect 23842 15348 23848 15360
rect 17184 15320 23704 15348
rect 23803 15320 23848 15348
rect 17184 15308 17190 15320
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 29638 15348 29644 15360
rect 29599 15320 29644 15348
rect 29638 15308 29644 15320
rect 29696 15308 29702 15360
rect 30006 15348 30012 15360
rect 29967 15320 30012 15348
rect 30006 15308 30012 15320
rect 30064 15308 30070 15360
rect 31573 15351 31631 15357
rect 31573 15317 31585 15351
rect 31619 15348 31631 15351
rect 32214 15348 32220 15360
rect 31619 15320 32220 15348
rect 31619 15317 31631 15320
rect 31573 15311 31631 15317
rect 32214 15308 32220 15320
rect 32272 15308 32278 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 13814 15144 13820 15156
rect 13775 15116 13820 15144
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 20806 15144 20812 15156
rect 19024 15116 20812 15144
rect 19024 15104 19030 15116
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 22741 15147 22799 15153
rect 22741 15113 22753 15147
rect 22787 15144 22799 15147
rect 32858 15144 32864 15156
rect 22787 15116 32864 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 32858 15104 32864 15116
rect 32916 15104 32922 15156
rect 34606 15144 34612 15156
rect 34567 15116 34612 15144
rect 34606 15104 34612 15116
rect 34664 15104 34670 15156
rect 35621 15147 35679 15153
rect 35621 15113 35633 15147
rect 35667 15144 35679 15147
rect 36446 15144 36452 15156
rect 35667 15116 36452 15144
rect 35667 15113 35679 15116
rect 35621 15107 35679 15113
rect 36446 15104 36452 15116
rect 36504 15104 36510 15156
rect 4706 15076 4712 15088
rect 4667 15048 4712 15076
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 8662 15076 8668 15088
rect 8623 15048 8668 15076
rect 8662 15036 8668 15048
rect 8720 15036 8726 15088
rect 13262 15036 13268 15088
rect 13320 15076 13326 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 13320 15048 13369 15076
rect 13320 15036 13326 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 13357 15039 13415 15045
rect 21634 15036 21640 15088
rect 21692 15076 21698 15088
rect 22281 15079 22339 15085
rect 22281 15076 22293 15079
rect 21692 15048 22293 15076
rect 21692 15036 21698 15048
rect 22281 15045 22293 15048
rect 22327 15045 22339 15079
rect 23566 15076 23572 15088
rect 22281 15039 22339 15045
rect 23216 15048 23572 15076
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 15008 1458 15020
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 1452 14980 2053 15008
rect 1452 14968 1458 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 4890 14968 4896 15020
rect 4948 15008 4954 15020
rect 4948 14980 4993 15008
rect 4948 14968 4954 14980
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7156 14980 7757 15008
rect 7156 14968 7162 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11296 14980 11529 15008
rect 11296 14968 11302 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13504 14980 14013 15008
rect 13504 14968 13510 14980
rect 14001 14977 14013 14980
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14240 14980 14289 15008
rect 14240 14968 14246 14980
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 15470 15008 15476 15020
rect 15431 14980 15476 15008
rect 14277 14971 14335 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 17678 14968 17684 15020
rect 17736 15008 17742 15020
rect 20533 15011 20591 15017
rect 20533 15008 20545 15011
rect 17736 14980 20545 15008
rect 17736 14968 17742 14980
rect 20533 14977 20545 14980
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21358 15008 21364 15020
rect 21131 14980 21364 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 3326 14940 3332 14952
rect 3287 14912 3332 14940
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14940 8539 14943
rect 8938 14940 8944 14952
rect 8527 14912 8944 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14909 10379 14943
rect 11698 14940 11704 14952
rect 11659 14912 11704 14940
rect 10321 14903 10379 14909
rect 3418 14832 3424 14884
rect 3476 14872 3482 14884
rect 10226 14872 10232 14884
rect 3476 14844 10232 14872
rect 3476 14832 3482 14844
rect 10226 14832 10232 14844
rect 10284 14872 10290 14884
rect 10336 14872 10364 14903
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 14090 14940 14096 14952
rect 14051 14912 14096 14940
rect 14090 14900 14096 14912
rect 14148 14940 14154 14952
rect 18506 14940 18512 14952
rect 14148 14912 18512 14940
rect 14148 14900 14154 14912
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 18782 14940 18788 14952
rect 18743 14912 18788 14940
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 19058 14940 19064 14952
rect 19019 14912 19064 14940
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 16666 14872 16672 14884
rect 10284 14844 16672 14872
rect 10284 14832 10290 14844
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 18524 14872 18552 14900
rect 19518 14872 19524 14884
rect 18524 14844 19524 14872
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 20548 14872 20576 14971
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 22554 15008 22560 15020
rect 22515 14980 22560 15008
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 23216 15017 23244 15048
rect 23566 15036 23572 15048
rect 23624 15076 23630 15088
rect 23845 15079 23903 15085
rect 23845 15076 23857 15079
rect 23624 15048 23857 15076
rect 23624 15036 23630 15048
rect 23845 15045 23857 15048
rect 23891 15045 23903 15079
rect 23845 15039 23903 15045
rect 28994 15036 29000 15088
rect 29052 15076 29058 15088
rect 29730 15076 29736 15088
rect 29052 15048 29736 15076
rect 29052 15036 29058 15048
rect 29730 15036 29736 15048
rect 29788 15076 29794 15088
rect 30282 15076 30288 15088
rect 29788 15048 30288 15076
rect 29788 15036 29794 15048
rect 30282 15036 30288 15048
rect 30340 15076 30346 15088
rect 30340 15048 30788 15076
rect 30340 15036 30346 15048
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23201 14971 23259 14977
rect 28169 15011 28227 15017
rect 28169 14977 28181 15011
rect 28215 15008 28227 15011
rect 28629 15011 28687 15017
rect 28629 15008 28641 15011
rect 28215 14980 28641 15008
rect 28215 14977 28227 14980
rect 28169 14971 28227 14977
rect 28629 14977 28641 14980
rect 28675 15008 28687 15011
rect 28810 15008 28816 15020
rect 28675 14980 28816 15008
rect 28675 14977 28687 14980
rect 28629 14971 28687 14977
rect 28810 14968 28816 14980
rect 28868 14968 28874 15020
rect 30466 15008 30472 15020
rect 30524 15017 30530 15020
rect 30760 15017 30788 15048
rect 30436 14980 30472 15008
rect 30466 14968 30472 14980
rect 30524 14971 30536 15017
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 32125 15011 32183 15017
rect 32125 15008 32137 15011
rect 30745 14971 30803 14977
rect 31726 14980 32137 15008
rect 30524 14968 30530 14971
rect 21174 14900 21180 14952
rect 21232 14940 21238 14952
rect 22002 14940 22008 14952
rect 21232 14912 22008 14940
rect 21232 14900 21238 14912
rect 22002 14900 22008 14912
rect 22060 14940 22066 14952
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 22060 14912 22385 14940
rect 22060 14900 22066 14912
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 21634 14872 21640 14884
rect 20548 14844 21640 14872
rect 21634 14832 21640 14844
rect 21692 14832 21698 14884
rect 28626 14832 28632 14884
rect 28684 14872 28690 14884
rect 28813 14875 28871 14881
rect 28813 14872 28825 14875
rect 28684 14844 28825 14872
rect 28684 14832 28690 14844
rect 28813 14841 28825 14844
rect 28859 14872 28871 14875
rect 28902 14872 28908 14884
rect 28859 14844 28908 14872
rect 28859 14841 28871 14844
rect 28813 14835 28871 14841
rect 28902 14832 28908 14844
rect 28960 14832 28966 14884
rect 29362 14872 29368 14884
rect 29323 14844 29368 14872
rect 29362 14832 29368 14844
rect 29420 14832 29426 14884
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 2774 14804 2780 14816
rect 1627 14776 2780 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 7742 14804 7748 14816
rect 7331 14776 7748 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 7926 14804 7932 14816
rect 7887 14776 7932 14804
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 14274 14804 14280 14816
rect 14235 14776 14280 14804
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 17954 14804 17960 14816
rect 17915 14776 17960 14804
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 21269 14807 21327 14813
rect 21269 14773 21281 14807
rect 21315 14804 21327 14807
rect 21910 14804 21916 14816
rect 21315 14776 21916 14804
rect 21315 14773 21327 14776
rect 21269 14767 21327 14773
rect 21910 14764 21916 14776
rect 21968 14764 21974 14816
rect 22370 14804 22376 14816
rect 22331 14776 22376 14804
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 23382 14804 23388 14816
rect 23343 14776 23388 14804
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 30098 14764 30104 14816
rect 30156 14804 30162 14816
rect 31481 14807 31539 14813
rect 31481 14804 31493 14807
rect 30156 14776 31493 14804
rect 30156 14764 30162 14776
rect 31481 14773 31493 14776
rect 31527 14804 31539 14807
rect 31726 14804 31754 14980
rect 32125 14977 32137 14980
rect 32171 14977 32183 15011
rect 32125 14971 32183 14977
rect 32214 14968 32220 15020
rect 32272 15008 32278 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 32272 14980 32321 15008
rect 32272 14968 32278 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 32493 15011 32551 15017
rect 32493 14977 32505 15011
rect 32539 15008 32551 15011
rect 35437 15011 35495 15017
rect 35437 15008 35449 15011
rect 32539 14980 35449 15008
rect 32539 14977 32551 14980
rect 32493 14971 32551 14977
rect 35437 14977 35449 14980
rect 35483 14977 35495 15011
rect 35437 14971 35495 14977
rect 31527 14776 31754 14804
rect 31527 14773 31539 14776
rect 31481 14767 31539 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 2498 14600 2504 14612
rect 2459 14572 2504 14600
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3108 14572 3801 14600
rect 3108 14560 3114 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 4120 14572 4169 14600
rect 4120 14560 4126 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 8938 14600 8944 14612
rect 8899 14572 8944 14600
rect 4157 14563 4215 14569
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12434 14600 12440 14612
rect 12400 14572 12440 14600
rect 12400 14560 12406 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 21910 14600 21916 14612
rect 21871 14572 21916 14600
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22189 14603 22247 14609
rect 22189 14569 22201 14603
rect 22235 14600 22247 14603
rect 22462 14600 22468 14612
rect 22235 14572 22468 14600
rect 22235 14569 22247 14572
rect 22189 14563 22247 14569
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22612 14572 22845 14600
rect 22612 14560 22618 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 22833 14563 22891 14569
rect 28721 14603 28779 14609
rect 28721 14569 28733 14603
rect 28767 14600 28779 14603
rect 28810 14600 28816 14612
rect 28767 14572 28816 14600
rect 28767 14569 28779 14572
rect 28721 14563 28779 14569
rect 16758 14532 16764 14544
rect 15304 14504 16764 14532
rect 2590 14464 2596 14476
rect 2551 14436 2596 14464
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4154 14464 4160 14476
rect 4111 14436 4160 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4154 14424 4160 14436
rect 4212 14464 4218 14476
rect 4798 14464 4804 14476
rect 4212 14436 4804 14464
rect 4212 14424 4218 14436
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 13081 14467 13139 14473
rect 13081 14464 13093 14467
rect 11756 14436 13093 14464
rect 11756 14424 11762 14436
rect 13081 14433 13093 14436
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 15304 14473 15332 14504
rect 16758 14492 16764 14504
rect 16816 14532 16822 14544
rect 19150 14532 19156 14544
rect 16816 14504 19156 14532
rect 16816 14492 16822 14504
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14332 14436 15025 14464
rect 14332 14424 14338 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 19058 14424 19064 14476
rect 19116 14464 19122 14476
rect 19116 14436 21128 14464
rect 19116 14424 19122 14436
rect 1578 14356 1584 14408
rect 1636 14396 1642 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 1636 14368 2513 14396
rect 1636 14356 1642 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 2774 14396 2780 14408
rect 2735 14368 2780 14396
rect 2501 14359 2559 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 3602 14356 3608 14408
rect 3660 14396 3666 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3660 14368 3985 14396
rect 3660 14356 3666 14368
rect 3973 14365 3985 14368
rect 4019 14396 4031 14399
rect 4706 14396 4712 14408
rect 4019 14368 4712 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 8018 14396 8024 14408
rect 7979 14368 8024 14396
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13320 14368 13369 14396
rect 13320 14356 13326 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 17954 14356 17960 14408
rect 18012 14396 18018 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 18012 14368 18245 14396
rect 18012 14356 18018 14368
rect 18233 14365 18245 14368
rect 18279 14396 18291 14399
rect 18874 14396 18880 14408
rect 18279 14368 18880 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 18966 14356 18972 14408
rect 19024 14396 19030 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19024 14368 19257 14396
rect 19024 14356 19030 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19518 14396 19524 14408
rect 19479 14368 19524 14396
rect 19245 14359 19303 14365
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 21100 14405 21128 14436
rect 21358 14424 21364 14476
rect 21416 14464 21422 14476
rect 21913 14467 21971 14473
rect 21416 14436 21864 14464
rect 21416 14424 21422 14436
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14396 21143 14399
rect 21726 14396 21732 14408
rect 21131 14368 21588 14396
rect 21687 14368 21732 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 4249 14331 4307 14337
rect 4249 14328 4261 14331
rect 3936 14300 4261 14328
rect 3936 14288 3942 14300
rect 4249 14297 4261 14300
rect 4295 14297 4307 14331
rect 9582 14328 9588 14340
rect 4249 14291 4307 14297
rect 6886 14300 9588 14328
rect 2958 14260 2964 14272
rect 2919 14232 2964 14260
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 6886 14260 6914 14300
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 14182 14288 14188 14340
rect 14240 14328 14246 14340
rect 17405 14331 17463 14337
rect 17405 14328 17417 14331
rect 14240 14300 17417 14328
rect 14240 14288 14246 14300
rect 17405 14297 17417 14300
rect 17451 14328 17463 14331
rect 18690 14328 18696 14340
rect 17451 14300 18696 14328
rect 17451 14297 17463 14300
rect 17405 14291 17463 14297
rect 7834 14260 7840 14272
rect 3476 14232 6914 14260
rect 7795 14232 7840 14260
rect 3476 14220 3482 14232
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 17497 14263 17555 14269
rect 17497 14229 17509 14263
rect 17543 14260 17555 14263
rect 17678 14260 17684 14272
rect 17543 14232 17684 14260
rect 17543 14229 17555 14232
rect 17497 14223 17555 14229
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 18064 14269 18092 14300
rect 18690 14288 18696 14300
rect 18748 14288 18754 14340
rect 21560 14328 21588 14368
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 21836 14396 21864 14436
rect 21913 14433 21925 14467
rect 21959 14464 21971 14467
rect 22094 14464 22100 14476
rect 21959 14436 22100 14464
rect 21959 14433 21971 14436
rect 21913 14427 21971 14433
rect 22094 14424 22100 14436
rect 22152 14464 22158 14476
rect 23382 14464 23388 14476
rect 22152 14436 23388 14464
rect 22152 14424 22158 14436
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14464 24731 14467
rect 25498 14464 25504 14476
rect 24719 14436 25504 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 25498 14424 25504 14436
rect 25556 14424 25562 14476
rect 25590 14424 25596 14476
rect 25648 14464 25654 14476
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 25648 14436 25697 14464
rect 25648 14424 25654 14436
rect 25685 14433 25697 14436
rect 25731 14433 25743 14467
rect 25685 14427 25743 14433
rect 22005 14399 22063 14405
rect 22005 14396 22017 14399
rect 21836 14368 22017 14396
rect 22005 14365 22017 14368
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14396 22707 14399
rect 23658 14396 23664 14408
rect 22695 14368 23664 14396
rect 22695 14365 22707 14368
rect 22649 14359 22707 14365
rect 22664 14328 22692 14359
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 24394 14396 24400 14408
rect 24355 14368 24400 14396
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 25961 14399 26019 14405
rect 25961 14365 25973 14399
rect 26007 14396 26019 14399
rect 27522 14396 27528 14408
rect 26007 14368 27528 14396
rect 26007 14365 26019 14368
rect 25961 14359 26019 14365
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14396 28227 14399
rect 28736 14396 28764 14563
rect 28810 14560 28816 14572
rect 28868 14560 28874 14612
rect 30466 14560 30472 14612
rect 30524 14600 30530 14612
rect 30561 14603 30619 14609
rect 30561 14600 30573 14603
rect 30524 14572 30573 14600
rect 30524 14560 30530 14572
rect 30561 14569 30573 14572
rect 30607 14569 30619 14603
rect 30561 14563 30619 14569
rect 34698 14560 34704 14612
rect 34756 14600 34762 14612
rect 34793 14603 34851 14609
rect 34793 14600 34805 14603
rect 34756 14572 34805 14600
rect 34756 14560 34762 14572
rect 34793 14569 34805 14572
rect 34839 14569 34851 14603
rect 34793 14563 34851 14569
rect 28215 14368 28764 14396
rect 28215 14365 28227 14368
rect 28169 14359 28227 14365
rect 29362 14356 29368 14408
rect 29420 14396 29426 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 29420 14368 29561 14396
rect 29420 14356 29426 14368
rect 29549 14365 29561 14368
rect 29595 14365 29607 14399
rect 29549 14359 29607 14365
rect 29638 14356 29644 14408
rect 29696 14396 29702 14408
rect 29733 14399 29791 14405
rect 29733 14396 29745 14399
rect 29696 14368 29745 14396
rect 29696 14356 29702 14368
rect 29733 14365 29745 14368
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14396 29975 14399
rect 30377 14399 30435 14405
rect 30377 14396 30389 14399
rect 29963 14368 30389 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 30377 14365 30389 14368
rect 30423 14365 30435 14399
rect 30377 14359 30435 14365
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 34701 14399 34759 14405
rect 34701 14396 34713 14399
rect 34572 14368 34713 14396
rect 34572 14356 34578 14368
rect 34701 14365 34713 14368
rect 34747 14396 34759 14399
rect 35345 14399 35403 14405
rect 35345 14396 35357 14399
rect 34747 14368 35357 14396
rect 34747 14365 34759 14368
rect 34701 14359 34759 14365
rect 35345 14365 35357 14368
rect 35391 14396 35403 14399
rect 35526 14396 35532 14408
rect 35391 14368 35532 14396
rect 35391 14365 35403 14368
rect 35345 14359 35403 14365
rect 35526 14356 35532 14368
rect 35584 14356 35590 14408
rect 21560 14300 22692 14328
rect 37369 14331 37427 14337
rect 37369 14297 37381 14331
rect 37415 14328 37427 14331
rect 38010 14328 38016 14340
rect 37415 14300 38016 14328
rect 37415 14297 37427 14300
rect 37369 14291 37427 14297
rect 38010 14288 38016 14300
rect 38068 14288 38074 14340
rect 18049 14263 18107 14269
rect 18049 14229 18061 14263
rect 18095 14229 18107 14263
rect 18049 14223 18107 14229
rect 21269 14263 21327 14269
rect 21269 14229 21281 14263
rect 21315 14260 21327 14263
rect 21358 14260 21364 14272
rect 21315 14232 21364 14260
rect 21315 14229 21327 14232
rect 21269 14223 21327 14229
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 28074 14260 28080 14272
rect 28035 14232 28080 14260
rect 28074 14220 28080 14232
rect 28132 14220 28138 14272
rect 37918 14260 37924 14272
rect 37879 14232 37924 14260
rect 37918 14220 37924 14232
rect 37976 14220 37982 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 3421 14059 3479 14065
rect 3421 14025 3433 14059
rect 3467 14056 3479 14059
rect 4614 14056 4620 14068
rect 3467 14028 4620 14056
rect 3467 14025 3479 14028
rect 3421 14019 3479 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 5074 14056 5080 14068
rect 5035 14028 5080 14056
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 13262 14056 13268 14068
rect 13223 14028 13268 14056
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 14645 14059 14703 14065
rect 14645 14025 14657 14059
rect 14691 14025 14703 14059
rect 14645 14019 14703 14025
rect 3878 13988 3884 14000
rect 3839 13960 3884 13988
rect 3878 13948 3884 13960
rect 3936 13988 3942 14000
rect 4341 13991 4399 13997
rect 4341 13988 4353 13991
rect 3936 13960 4353 13988
rect 3936 13948 3942 13960
rect 4341 13957 4353 13960
rect 4387 13988 4399 13991
rect 7926 13988 7932 14000
rect 4387 13960 4660 13988
rect 7887 13960 7932 13988
rect 4387 13957 4399 13960
rect 4341 13951 4399 13957
rect 4632 13932 4660 13960
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 13725 13991 13783 13997
rect 13725 13957 13737 13991
rect 13771 13988 13783 13991
rect 14182 13988 14188 14000
rect 13771 13960 14188 13988
rect 13771 13957 13783 13960
rect 13725 13951 13783 13957
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 3602 13920 3608 13932
rect 3563 13892 3608 13920
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 3789 13855 3847 13861
rect 3789 13821 3801 13855
rect 3835 13852 3847 13855
rect 4154 13852 4160 13864
rect 3835 13824 4160 13852
rect 3835 13821 3847 13824
rect 3789 13815 3847 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 4540 13852 4568 13883
rect 4614 13880 4620 13932
rect 4672 13880 4678 13932
rect 7742 13920 7748 13932
rect 7703 13892 7748 13920
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 12342 13920 12348 13932
rect 12303 13892 12348 13920
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 13446 13920 13452 13932
rect 13407 13892 13452 13920
rect 13446 13880 13452 13892
rect 13504 13920 13510 13932
rect 14660 13920 14688 14019
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 22060 14028 22109 14056
rect 22060 14016 22066 14028
rect 22097 14025 22109 14028
rect 22143 14025 22155 14059
rect 32582 14056 32588 14068
rect 32495 14028 32588 14056
rect 22097 14019 22155 14025
rect 32582 14016 32588 14028
rect 32640 14056 32646 14068
rect 34790 14056 34796 14068
rect 32640 14028 34796 14056
rect 32640 14016 32646 14028
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 21358 13988 21364 14000
rect 15252 13960 18920 13988
rect 15252 13948 15258 13960
rect 13504 13892 14688 13920
rect 14829 13923 14887 13929
rect 13504 13880 13510 13892
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 14875 13892 17509 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 17497 13889 17509 13892
rect 17543 13920 17555 13923
rect 18782 13920 18788 13932
rect 17543 13892 18788 13920
rect 17543 13889 17555 13892
rect 17497 13883 17555 13889
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 4798 13852 4804 13864
rect 4540 13824 4804 13852
rect 4798 13812 4804 13824
rect 4856 13852 4862 13864
rect 5074 13852 5080 13864
rect 4856 13824 5080 13852
rect 4856 13812 4862 13824
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 8294 13852 8300 13864
rect 8255 13824 8300 13852
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 14090 13852 14096 13864
rect 13679 13824 14096 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 17218 13852 17224 13864
rect 17179 13824 17224 13852
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 18892 13852 18920 13960
rect 20548 13960 21364 13988
rect 20548 13929 20576 13960
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 34054 13988 34060 14000
rect 34015 13960 34060 13988
rect 34054 13948 34060 13960
rect 34112 13948 34118 14000
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20772 13892 20821 13920
rect 20772 13880 20778 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 23900 13892 24593 13920
rect 23900 13880 23906 13892
rect 24581 13889 24593 13892
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 29914 13880 29920 13932
rect 29972 13920 29978 13932
rect 30561 13923 30619 13929
rect 30561 13920 30573 13923
rect 29972 13892 30573 13920
rect 29972 13880 29978 13892
rect 30561 13889 30573 13892
rect 30607 13920 30619 13923
rect 32401 13923 32459 13929
rect 32401 13920 32413 13923
rect 30607 13892 32413 13920
rect 30607 13889 30619 13892
rect 30561 13883 30619 13889
rect 32401 13889 32413 13892
rect 32447 13889 32459 13923
rect 32401 13883 32459 13889
rect 20622 13852 20628 13864
rect 18892 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 24857 13855 24915 13861
rect 24857 13821 24869 13855
rect 24903 13852 24915 13855
rect 25958 13852 25964 13864
rect 24903 13824 25964 13852
rect 24903 13821 24915 13824
rect 24857 13815 24915 13821
rect 25958 13812 25964 13824
rect 26016 13812 26022 13864
rect 29362 13812 29368 13864
rect 29420 13852 29426 13864
rect 30009 13855 30067 13861
rect 30009 13852 30021 13855
rect 29420 13824 30021 13852
rect 29420 13812 29426 13824
rect 30009 13821 30021 13824
rect 30055 13852 30067 13855
rect 30098 13852 30104 13864
rect 30055 13824 30104 13852
rect 30055 13821 30067 13824
rect 30009 13815 30067 13821
rect 30098 13812 30104 13824
rect 30156 13852 30162 13864
rect 33873 13855 33931 13861
rect 30156 13824 30788 13852
rect 30156 13812 30162 13824
rect 30760 13793 30788 13824
rect 33873 13821 33885 13855
rect 33919 13852 33931 13855
rect 35434 13852 35440 13864
rect 33919 13824 35440 13852
rect 33919 13821 33931 13824
rect 33873 13815 33931 13821
rect 35434 13812 35440 13824
rect 35492 13812 35498 13864
rect 35526 13812 35532 13864
rect 35584 13852 35590 13864
rect 35584 13824 35629 13852
rect 35584 13812 35590 13824
rect 30745 13787 30803 13793
rect 30745 13753 30757 13787
rect 30791 13753 30803 13787
rect 30745 13747 30803 13753
rect 3881 13719 3939 13725
rect 3881 13685 3893 13719
rect 3927 13716 3939 13719
rect 4062 13716 4068 13728
rect 3927 13688 4068 13716
rect 3927 13685 3939 13688
rect 3881 13679 3939 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 12526 13716 12532 13728
rect 12487 13688 12532 13716
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 13725 13719 13783 13725
rect 13725 13685 13737 13719
rect 13771 13716 13783 13719
rect 13814 13716 13820 13728
rect 13771 13688 13820 13716
rect 13771 13685 13783 13688
rect 13725 13679 13783 13685
rect 13814 13676 13820 13688
rect 13872 13716 13878 13728
rect 14274 13716 14280 13728
rect 13872 13688 14280 13716
rect 13872 13676 13878 13688
rect 14274 13676 14280 13688
rect 14332 13676 14338 13728
rect 20346 13716 20352 13728
rect 20307 13688 20352 13716
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 20806 13716 20812 13728
rect 20767 13688 20812 13716
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 2498 13512 2504 13524
rect 1627 13484 2504 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 4706 13512 4712 13524
rect 4479 13484 4712 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 17402 13512 17408 13524
rect 17363 13484 17408 13512
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 20806 13472 20812 13524
rect 20864 13512 20870 13524
rect 21085 13515 21143 13521
rect 21085 13512 21097 13515
rect 20864 13484 21097 13512
rect 20864 13472 20870 13484
rect 21085 13481 21097 13484
rect 21131 13512 21143 13515
rect 21910 13512 21916 13524
rect 21131 13484 21916 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 24394 13512 24400 13524
rect 22066 13484 24400 13512
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 5077 13447 5135 13453
rect 5077 13444 5089 13447
rect 4120 13416 5089 13444
rect 4120 13404 4126 13416
rect 5077 13413 5089 13416
rect 5123 13413 5135 13447
rect 5077 13407 5135 13413
rect 17865 13447 17923 13453
rect 17865 13413 17877 13447
rect 17911 13444 17923 13447
rect 22066 13444 22094 13484
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 29914 13472 29920 13524
rect 29972 13512 29978 13524
rect 30098 13512 30104 13524
rect 29972 13484 30104 13512
rect 29972 13472 29978 13484
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 17911 13416 22094 13444
rect 22189 13447 22247 13453
rect 17911 13413 17923 13416
rect 17865 13407 17923 13413
rect 22189 13413 22201 13447
rect 22235 13444 22247 13447
rect 22235 13416 25636 13444
rect 22235 13413 22247 13416
rect 22189 13407 22247 13413
rect 5534 13376 5540 13388
rect 4632 13348 5540 13376
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13308 1458 13320
rect 4632 13317 4660 13348
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 17402 13376 17408 13388
rect 16531 13348 17408 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 17586 13376 17592 13388
rect 17547 13348 17592 13376
rect 17586 13336 17592 13348
rect 17644 13376 17650 13388
rect 19426 13376 19432 13388
rect 17644 13348 19432 13376
rect 17644 13336 17650 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 20165 13379 20223 13385
rect 20165 13345 20177 13379
rect 20211 13376 20223 13379
rect 20346 13376 20352 13388
rect 20211 13348 20352 13376
rect 20211 13345 20223 13348
rect 20165 13339 20223 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 25608 13385 25636 13416
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 20680 13348 21005 13376
rect 20680 13336 20686 13348
rect 20993 13345 21005 13348
rect 21039 13376 21051 13379
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21039 13348 21833 13376
rect 21039 13345 21051 13348
rect 20993 13339 21051 13345
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 25593 13379 25651 13385
rect 25593 13345 25605 13379
rect 25639 13345 25651 13379
rect 26878 13376 26884 13388
rect 26839 13348 26884 13376
rect 25593 13339 25651 13345
rect 26878 13336 26884 13348
rect 26936 13336 26942 13388
rect 27522 13336 27528 13388
rect 27580 13376 27586 13388
rect 28537 13379 28595 13385
rect 28537 13376 28549 13379
rect 27580 13348 28549 13376
rect 27580 13336 27586 13348
rect 28537 13345 28549 13348
rect 28583 13345 28595 13379
rect 28537 13339 28595 13345
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1452 13280 2053 13308
rect 1452 13268 1458 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4019 13280 4629 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 5258 13308 5264 13320
rect 5219 13280 5264 13308
rect 4617 13271 4675 13277
rect 5258 13268 5264 13280
rect 5316 13308 5322 13320
rect 5721 13311 5779 13317
rect 5721 13308 5733 13311
rect 5316 13280 5733 13308
rect 5316 13268 5322 13280
rect 5721 13277 5733 13280
rect 5767 13308 5779 13311
rect 6546 13308 6552 13320
rect 5767 13280 6552 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 7742 13308 7748 13320
rect 7703 13280 7748 13308
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17276 13280 17693 13308
rect 17276 13268 17282 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 19978 13308 19984 13320
rect 19935 13280 19984 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 20772 13280 20821 13308
rect 20772 13268 20778 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 21085 13271 21143 13277
rect 17405 13243 17463 13249
rect 17405 13209 17417 13243
rect 17451 13240 17463 13243
rect 17494 13240 17500 13252
rect 17451 13212 17500 13240
rect 17451 13209 17463 13212
rect 17405 13203 17463 13209
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 21100 13240 21128 13271
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 22002 13308 22008 13320
rect 21963 13280 22008 13308
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 25866 13308 25872 13320
rect 25827 13280 25872 13308
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 33410 13308 33416 13320
rect 28767 13280 33416 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 33410 13268 33416 13280
rect 33468 13268 33474 13320
rect 34698 13268 34704 13320
rect 34756 13308 34762 13320
rect 34793 13311 34851 13317
rect 34793 13308 34805 13311
rect 34756 13280 34805 13308
rect 34756 13268 34762 13280
rect 34793 13277 34805 13280
rect 34839 13277 34851 13311
rect 34793 13271 34851 13277
rect 34977 13311 35035 13317
rect 34977 13277 34989 13311
rect 35023 13277 35035 13311
rect 34977 13271 35035 13277
rect 21358 13240 21364 13252
rect 21100 13212 21364 13240
rect 21358 13200 21364 13212
rect 21416 13240 21422 13252
rect 22020 13240 22048 13268
rect 21416 13212 22048 13240
rect 21416 13200 21422 13212
rect 28074 13200 28080 13252
rect 28132 13240 28138 13252
rect 30009 13243 30067 13249
rect 30009 13240 30021 13243
rect 28132 13212 30021 13240
rect 28132 13200 28138 13212
rect 30009 13209 30021 13212
rect 30055 13209 30067 13243
rect 30009 13203 30067 13209
rect 34422 13200 34428 13252
rect 34480 13240 34486 13252
rect 34992 13240 35020 13271
rect 34480 13212 35020 13240
rect 34480 13200 34486 13212
rect 21269 13175 21327 13181
rect 21269 13141 21281 13175
rect 21315 13172 21327 13175
rect 22186 13172 22192 13184
rect 21315 13144 22192 13172
rect 21315 13141 21327 13144
rect 21269 13135 21327 13141
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 34885 13175 34943 13181
rect 34885 13141 34897 13175
rect 34931 13172 34943 13175
rect 35250 13172 35256 13184
rect 34931 13144 35256 13172
rect 34931 13141 34943 13144
rect 34885 13135 34943 13141
rect 35250 13132 35256 13144
rect 35308 13132 35314 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7834 12928 7840 12980
rect 7892 12928 7898 12980
rect 10612 12940 18184 12968
rect 7852 12900 7880 12928
rect 7929 12903 7987 12909
rect 7929 12900 7941 12903
rect 7852 12872 7941 12900
rect 7929 12869 7941 12872
rect 7975 12869 7987 12903
rect 9582 12900 9588 12912
rect 9495 12872 9588 12900
rect 7929 12863 7987 12869
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 10612 12900 10640 12940
rect 9640 12872 10640 12900
rect 12621 12903 12679 12909
rect 9640 12860 9646 12872
rect 12621 12869 12633 12903
rect 12667 12900 12679 12903
rect 13170 12900 13176 12912
rect 12667 12872 13176 12900
rect 12667 12869 12679 12872
rect 12621 12863 12679 12869
rect 13170 12860 13176 12872
rect 13228 12900 13234 12912
rect 18156 12909 18184 12940
rect 21726 12928 21732 12980
rect 21784 12968 21790 12980
rect 21784 12940 22968 12968
rect 21784 12928 21790 12940
rect 13541 12903 13599 12909
rect 13541 12900 13553 12903
rect 13228 12872 13553 12900
rect 13228 12860 13234 12872
rect 13541 12869 13553 12872
rect 13587 12869 13599 12903
rect 13541 12863 13599 12869
rect 18141 12903 18199 12909
rect 18141 12869 18153 12903
rect 18187 12900 18199 12903
rect 19058 12900 19064 12912
rect 18187 12872 19064 12900
rect 18187 12869 18199 12872
rect 18141 12863 18199 12869
rect 19058 12860 19064 12872
rect 19116 12860 19122 12912
rect 19797 12903 19855 12909
rect 19797 12869 19809 12903
rect 19843 12900 19855 12903
rect 19978 12900 19984 12912
rect 19843 12872 19984 12900
rect 19843 12869 19855 12872
rect 19797 12863 19855 12869
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 21928 12909 21956 12940
rect 21913 12903 21971 12909
rect 21913 12869 21925 12903
rect 21959 12869 21971 12903
rect 21913 12863 21971 12869
rect 22002 12860 22008 12912
rect 22060 12900 22066 12912
rect 22940 12909 22968 12940
rect 29086 12928 29092 12980
rect 29144 12968 29150 12980
rect 29730 12968 29736 12980
rect 29144 12940 29736 12968
rect 29144 12928 29150 12940
rect 29730 12928 29736 12940
rect 29788 12928 29794 12980
rect 34609 12971 34667 12977
rect 34609 12937 34621 12971
rect 34655 12968 34667 12971
rect 34790 12968 34796 12980
rect 34655 12940 34796 12968
rect 34655 12937 34667 12940
rect 34609 12931 34667 12937
rect 34790 12928 34796 12940
rect 34848 12928 34854 12980
rect 22925 12903 22983 12909
rect 22060 12860 22094 12900
rect 22925 12869 22937 12903
rect 22971 12900 22983 12903
rect 23845 12903 23903 12909
rect 23845 12900 23857 12903
rect 22971 12872 23857 12900
rect 22971 12869 22983 12872
rect 22925 12863 22983 12869
rect 23845 12869 23857 12872
rect 23891 12869 23903 12903
rect 23845 12863 23903 12869
rect 27433 12903 27491 12909
rect 27433 12869 27445 12903
rect 27479 12900 27491 12903
rect 27706 12900 27712 12912
rect 27479 12872 27712 12900
rect 27479 12869 27491 12872
rect 27433 12863 27491 12869
rect 27706 12860 27712 12872
rect 27764 12900 27770 12912
rect 28810 12900 28816 12912
rect 27764 12872 28816 12900
rect 27764 12860 27770 12872
rect 28810 12860 28816 12872
rect 28868 12860 28874 12912
rect 7742 12832 7748 12844
rect 7703 12804 7748 12832
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 12345 12835 12403 12841
rect 12345 12801 12357 12835
rect 12391 12832 12403 12835
rect 12434 12832 12440 12844
rect 12391 12804 12440 12832
rect 12391 12801 12403 12804
rect 12345 12795 12403 12801
rect 12434 12792 12440 12804
rect 12492 12832 12498 12844
rect 13265 12835 13323 12841
rect 13265 12832 13277 12835
rect 12492 12804 13277 12832
rect 12492 12792 12498 12804
rect 13265 12801 13277 12804
rect 13311 12832 13323 12835
rect 13446 12832 13452 12844
rect 13311 12804 13452 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 22066 12832 22094 12860
rect 22189 12835 22247 12841
rect 22189 12832 22201 12835
rect 22066 12804 22201 12832
rect 22189 12801 22201 12804
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22554 12792 22560 12844
rect 22612 12832 22618 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 22612 12804 23213 12832
rect 22612 12792 22618 12804
rect 23201 12801 23213 12804
rect 23247 12832 23259 12835
rect 24121 12835 24179 12841
rect 24121 12832 24133 12835
rect 23247 12804 24133 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 24121 12801 24133 12804
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 25866 12792 25872 12844
rect 25924 12832 25930 12844
rect 34808 12832 34836 12928
rect 35069 12835 35127 12841
rect 35069 12832 35081 12835
rect 25924 12804 27568 12832
rect 34808 12804 35081 12832
rect 25924 12792 25930 12804
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12764 3019 12767
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 3007 12736 3433 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3421 12733 3433 12736
rect 3467 12733 3479 12767
rect 3602 12764 3608 12776
rect 3563 12736 3608 12764
rect 3421 12727 3479 12733
rect 3602 12724 3608 12736
rect 3660 12724 3666 12776
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12764 5319 12767
rect 12526 12764 12532 12776
rect 5307 12736 6914 12764
rect 12487 12736 12532 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 6886 12696 6914 12736
rect 12526 12724 12532 12736
rect 12584 12764 12590 12776
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 12584 12736 13369 12764
rect 12584 12724 12590 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 9674 12696 9680 12708
rect 6886 12668 9680 12696
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 17681 12699 17739 12705
rect 12636 12668 13584 12696
rect 12636 12640 12664 12668
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 11698 12628 11704 12640
rect 10275 12600 11704 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11848 12600 12173 12628
rect 11848 12588 11854 12600
rect 12161 12597 12173 12600
rect 12207 12597 12219 12631
rect 12618 12628 12624 12640
rect 12531 12600 12624 12628
rect 12161 12591 12219 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 13078 12628 13084 12640
rect 13039 12600 13084 12628
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13556 12637 13584 12668
rect 17681 12665 17693 12699
rect 17727 12696 17739 12699
rect 19996 12696 20024 12727
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22152 12736 23029 12764
rect 22152 12724 22158 12736
rect 23017 12733 23029 12736
rect 23063 12764 23075 12767
rect 23937 12767 23995 12773
rect 23937 12764 23949 12767
rect 23063 12736 23949 12764
rect 23063 12733 23075 12736
rect 23017 12727 23075 12733
rect 23937 12733 23949 12736
rect 23983 12733 23995 12767
rect 27540 12764 27568 12804
rect 35069 12801 35081 12804
rect 35115 12801 35127 12835
rect 35250 12832 35256 12844
rect 35211 12804 35256 12832
rect 35069 12795 35127 12801
rect 35250 12792 35256 12804
rect 35308 12792 35314 12844
rect 35345 12835 35403 12841
rect 35345 12801 35357 12835
rect 35391 12801 35403 12835
rect 35345 12795 35403 12801
rect 29089 12767 29147 12773
rect 29089 12764 29101 12767
rect 27540 12736 29101 12764
rect 23937 12727 23995 12733
rect 29089 12733 29101 12736
rect 29135 12733 29147 12767
rect 29270 12764 29276 12776
rect 29231 12736 29276 12764
rect 29089 12727 29147 12733
rect 29270 12724 29276 12736
rect 29328 12724 29334 12776
rect 33502 12724 33508 12776
rect 33560 12764 33566 12776
rect 34422 12764 34428 12776
rect 33560 12736 34428 12764
rect 33560 12724 33566 12736
rect 34422 12724 34428 12736
rect 34480 12764 34486 12776
rect 35360 12764 35388 12795
rect 35434 12792 35440 12844
rect 35492 12832 35498 12844
rect 35492 12804 35537 12832
rect 35492 12792 35498 12804
rect 34480 12736 35388 12764
rect 34480 12724 34486 12736
rect 17727 12668 20024 12696
rect 22940 12668 23888 12696
rect 17727 12665 17739 12668
rect 17681 12659 17739 12665
rect 13541 12631 13599 12637
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 13814 12628 13820 12640
rect 13587 12600 13820 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 21910 12628 21916 12640
rect 21871 12600 21916 12628
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22373 12631 22431 12637
rect 22373 12628 22385 12631
rect 22336 12600 22385 12628
rect 22336 12588 22342 12600
rect 22373 12597 22385 12600
rect 22419 12597 22431 12631
rect 22373 12591 22431 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22940 12637 22968 12668
rect 22925 12631 22983 12637
rect 22925 12628 22937 12631
rect 22520 12600 22937 12628
rect 22520 12588 22526 12600
rect 22925 12597 22937 12600
rect 22971 12597 22983 12631
rect 22925 12591 22983 12597
rect 23385 12631 23443 12637
rect 23385 12597 23397 12631
rect 23431 12628 23443 12631
rect 23750 12628 23756 12640
rect 23431 12600 23756 12628
rect 23431 12597 23443 12600
rect 23385 12591 23443 12597
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 23860 12637 23888 12668
rect 23845 12631 23903 12637
rect 23845 12597 23857 12631
rect 23891 12597 23903 12631
rect 24302 12628 24308 12640
rect 24263 12600 24308 12628
rect 23845 12591 23903 12597
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 26878 12588 26884 12640
rect 26936 12628 26942 12640
rect 30466 12628 30472 12640
rect 26936 12600 30472 12628
rect 26936 12588 26942 12600
rect 30466 12588 30472 12600
rect 30524 12588 30530 12640
rect 35713 12631 35771 12637
rect 35713 12597 35725 12631
rect 35759 12628 35771 12631
rect 36078 12628 36084 12640
rect 35759 12600 36084 12628
rect 35759 12597 35771 12600
rect 35713 12591 35771 12597
rect 36078 12588 36084 12600
rect 36136 12588 36142 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 3602 12424 3608 12436
rect 3283 12396 3608 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 4062 12424 4068 12436
rect 4023 12396 4068 12424
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 6273 12427 6331 12433
rect 6273 12393 6285 12427
rect 6319 12424 6331 12427
rect 6454 12424 6460 12436
rect 6319 12396 6460 12424
rect 6319 12393 6331 12396
rect 6273 12387 6331 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 17034 12424 17040 12436
rect 16995 12396 17040 12424
rect 17034 12384 17040 12396
rect 17092 12424 17098 12436
rect 17402 12424 17408 12436
rect 17092 12396 17408 12424
rect 17092 12384 17098 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 20438 12424 20444 12436
rect 17552 12396 20444 12424
rect 17552 12384 17558 12396
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 12158 12356 12164 12368
rect 9732 12328 12164 12356
rect 9732 12316 9738 12328
rect 4706 12288 4712 12300
rect 3988 12260 4712 12288
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12220 1458 12232
rect 3988 12229 4016 12260
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 11256 12297 11284 12328
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 17512 12356 17540 12384
rect 16960 12328 17540 12356
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12257 11299 12291
rect 11698 12288 11704 12300
rect 11659 12260 11704 12288
rect 11241 12251 11299 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 12526 12288 12532 12300
rect 12487 12260 12532 12288
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1452 12192 2053 12220
rect 1452 12180 1458 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3973 12223 4031 12229
rect 3099 12192 3832 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 2590 12084 2596 12096
rect 1627 12056 2596 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 3804 12093 3832 12192
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4249 12223 4307 12229
rect 4120 12192 4165 12220
rect 4120 12180 4126 12192
rect 4249 12189 4261 12223
rect 4295 12220 4307 12223
rect 4614 12220 4620 12232
rect 4295 12192 4620 12220
rect 4295 12189 4307 12192
rect 4249 12183 4307 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4890 12220 4896 12232
rect 4851 12192 4896 12220
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9217 12223 9275 12229
rect 9217 12220 9229 12223
rect 9180 12192 9229 12220
rect 9180 12180 9186 12192
rect 9217 12189 9229 12192
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 16960 12229 16988 12328
rect 17126 12288 17132 12300
rect 17039 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12288 17190 12300
rect 17586 12288 17592 12300
rect 17184 12260 17592 12288
rect 17184 12248 17190 12260
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 18156 12297 18184 12396
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 21634 12424 21640 12436
rect 21595 12396 21640 12424
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22462 12424 22468 12436
rect 22423 12396 22468 12424
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 32582 12424 32588 12436
rect 32543 12396 32588 12424
rect 32582 12384 32588 12396
rect 32640 12384 32646 12436
rect 35434 12384 35440 12436
rect 35492 12424 35498 12436
rect 35802 12424 35808 12436
rect 35492 12396 35808 12424
rect 35492 12384 35498 12396
rect 35802 12384 35808 12396
rect 35860 12424 35866 12436
rect 37369 12427 37427 12433
rect 37369 12424 37381 12427
rect 35860 12396 37381 12424
rect 35860 12384 35866 12396
rect 37369 12393 37381 12396
rect 37415 12393 37427 12427
rect 37369 12387 37427 12393
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 22152 12260 22293 12288
rect 22152 12248 22158 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 25958 12288 25964 12300
rect 25919 12260 25964 12288
rect 22281 12251 22339 12257
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 27246 12288 27252 12300
rect 27207 12260 27252 12288
rect 27246 12248 27252 12260
rect 27304 12248 27310 12300
rect 29730 12248 29736 12300
rect 29788 12288 29794 12300
rect 29825 12291 29883 12297
rect 29825 12288 29837 12291
rect 29788 12260 29837 12288
rect 29788 12248 29794 12260
rect 29825 12257 29837 12260
rect 29871 12257 29883 12291
rect 29825 12251 29883 12257
rect 13357 12223 13415 12229
rect 13357 12220 13369 12223
rect 12492 12192 12537 12220
rect 12636 12192 13369 12220
rect 12492 12180 12498 12192
rect 11514 12152 11520 12164
rect 11475 12124 11520 12152
rect 11514 12112 11520 12124
rect 11572 12112 11578 12164
rect 12636 12152 12664 12192
rect 13357 12189 13369 12192
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12189 17003 12223
rect 17218 12220 17224 12232
rect 17179 12192 17224 12220
rect 16945 12183 17003 12189
rect 11624 12124 12664 12152
rect 12713 12155 12771 12161
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4709 12087 4767 12093
rect 4709 12084 4721 12087
rect 4212 12056 4721 12084
rect 4212 12044 4218 12056
rect 4709 12053 4721 12056
rect 4755 12053 4767 12087
rect 4709 12047 4767 12053
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 11624 12084 11652 12124
rect 12713 12121 12725 12155
rect 12759 12121 12771 12155
rect 13372 12152 13400 12183
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 17862 12220 17868 12232
rect 17823 12192 17868 12220
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 22189 12223 22247 12229
rect 22189 12220 22201 12223
rect 21692 12192 22201 12220
rect 21692 12180 21698 12192
rect 22189 12189 22201 12192
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 22465 12223 22523 12229
rect 22465 12189 22477 12223
rect 22511 12220 22523 12223
rect 22554 12220 22560 12232
rect 22511 12192 22560 12220
rect 22511 12189 22523 12192
rect 22465 12183 22523 12189
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 25222 12220 25228 12232
rect 25183 12192 25228 12220
rect 25222 12180 25228 12192
rect 25280 12180 25286 12232
rect 25777 12223 25835 12229
rect 25777 12189 25789 12223
rect 25823 12189 25835 12223
rect 25777 12183 25835 12189
rect 14185 12155 14243 12161
rect 14185 12152 14197 12155
rect 13372 12124 14197 12152
rect 12713 12115 12771 12121
rect 14185 12121 14197 12124
rect 14231 12152 14243 12155
rect 18874 12152 18880 12164
rect 14231 12124 18880 12152
rect 14231 12121 14243 12124
rect 14185 12115 14243 12121
rect 12250 12084 12256 12096
rect 8260 12056 11652 12084
rect 12211 12056 12256 12084
rect 8260 12044 8266 12056
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12728 12084 12756 12115
rect 18874 12112 18880 12124
rect 18932 12112 18938 12164
rect 25038 12152 25044 12164
rect 24999 12124 25044 12152
rect 25038 12112 25044 12124
rect 25096 12112 25102 12164
rect 25792 12152 25820 12183
rect 32582 12180 32588 12232
rect 32640 12220 32646 12232
rect 33045 12223 33103 12229
rect 33045 12220 33057 12223
rect 32640 12192 33057 12220
rect 32640 12180 32646 12192
rect 33045 12189 33057 12192
rect 33091 12189 33103 12223
rect 33045 12183 33103 12189
rect 33134 12180 33140 12232
rect 33192 12220 33198 12232
rect 33229 12223 33287 12229
rect 33229 12220 33241 12223
rect 33192 12192 33241 12220
rect 33192 12180 33198 12192
rect 33229 12189 33241 12192
rect 33275 12189 33287 12223
rect 33229 12183 33287 12189
rect 33321 12223 33379 12229
rect 33321 12189 33333 12223
rect 33367 12189 33379 12223
rect 33321 12183 33379 12189
rect 27430 12152 27436 12164
rect 25792 12124 27436 12152
rect 27430 12112 27436 12124
rect 27488 12112 27494 12164
rect 29914 12112 29920 12164
rect 29972 12152 29978 12164
rect 30070 12155 30128 12161
rect 30070 12152 30082 12155
rect 29972 12124 30082 12152
rect 29972 12112 29978 12124
rect 30070 12121 30082 12124
rect 30116 12121 30128 12155
rect 33336 12152 33364 12183
rect 33410 12180 33416 12232
rect 33468 12220 33474 12232
rect 35989 12223 36047 12229
rect 35989 12220 36001 12223
rect 33468 12192 33513 12220
rect 35866 12192 36001 12220
rect 33468 12180 33474 12192
rect 33502 12152 33508 12164
rect 33336 12124 33508 12152
rect 30070 12115 30128 12121
rect 33502 12112 33508 12124
rect 33560 12112 33566 12164
rect 13170 12084 13176 12096
rect 12728 12056 13176 12084
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 17405 12087 17463 12093
rect 17405 12053 17417 12087
rect 17451 12084 17463 12087
rect 18506 12084 18512 12096
rect 17451 12056 18512 12084
rect 17451 12053 17463 12056
rect 17405 12047 17463 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 22649 12087 22707 12093
rect 22649 12053 22661 12087
rect 22695 12084 22707 12087
rect 23106 12084 23112 12096
rect 22695 12056 23112 12084
rect 22695 12053 22707 12056
rect 22649 12047 22707 12053
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 31205 12087 31263 12093
rect 31205 12053 31217 12087
rect 31251 12084 31263 12087
rect 32398 12084 32404 12096
rect 31251 12056 32404 12084
rect 31251 12053 31263 12056
rect 31205 12047 31263 12053
rect 32398 12044 32404 12056
rect 32456 12044 32462 12096
rect 33686 12084 33692 12096
rect 33647 12056 33692 12084
rect 33686 12044 33692 12056
rect 33744 12044 33750 12096
rect 35342 12044 35348 12096
rect 35400 12084 35406 12096
rect 35437 12087 35495 12093
rect 35437 12084 35449 12087
rect 35400 12056 35449 12084
rect 35400 12044 35406 12056
rect 35437 12053 35449 12056
rect 35483 12084 35495 12087
rect 35866 12084 35894 12192
rect 35989 12189 36001 12192
rect 36035 12189 36047 12223
rect 35989 12183 36047 12189
rect 36078 12180 36084 12232
rect 36136 12220 36142 12232
rect 36245 12223 36303 12229
rect 36245 12220 36257 12223
rect 36136 12192 36257 12220
rect 36136 12180 36142 12192
rect 36245 12189 36257 12192
rect 36291 12189 36303 12223
rect 36245 12183 36303 12189
rect 35483 12056 35894 12084
rect 35483 12053 35495 12056
rect 35437 12047 35495 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11880 6610 11892
rect 7650 11880 7656 11892
rect 6604 11852 7656 11880
rect 6604 11840 6610 11852
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 8343 11852 17785 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 17773 11849 17785 11852
rect 17819 11880 17831 11883
rect 17862 11880 17868 11892
rect 17819 11852 17868 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 28353 11883 28411 11889
rect 28353 11849 28365 11883
rect 28399 11880 28411 11883
rect 28902 11880 28908 11892
rect 28399 11852 28908 11880
rect 28399 11849 28411 11852
rect 28353 11843 28411 11849
rect 28902 11840 28908 11852
rect 28960 11840 28966 11892
rect 29730 11840 29736 11892
rect 29788 11880 29794 11892
rect 33229 11883 33287 11889
rect 33229 11880 33241 11883
rect 29788 11852 33241 11880
rect 29788 11840 29794 11852
rect 33229 11849 33241 11852
rect 33275 11849 33287 11883
rect 33229 11843 33287 11849
rect 4154 11812 4160 11824
rect 4115 11784 4160 11812
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 10962 11812 10968 11824
rect 6886 11784 10968 11812
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11744 6423 11747
rect 6454 11744 6460 11756
rect 6411 11716 6460 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4614 11676 4620 11688
rect 4019 11648 4620 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 5813 11679 5871 11685
rect 5813 11645 5825 11679
rect 5859 11676 5871 11679
rect 6886 11676 6914 11784
rect 10962 11772 10968 11784
rect 11020 11772 11026 11824
rect 13170 11812 13176 11824
rect 13083 11784 13176 11812
rect 13170 11772 13176 11784
rect 13228 11812 13234 11824
rect 13538 11812 13544 11824
rect 13228 11784 13544 11812
rect 13228 11772 13234 11784
rect 13538 11772 13544 11784
rect 13596 11772 13602 11824
rect 17218 11812 17224 11824
rect 15856 11784 17224 11812
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7432 11716 8033 11744
rect 7432 11704 7438 11716
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 9122 11744 9128 11756
rect 9083 11716 9128 11744
rect 8021 11707 8079 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11572 11716 12081 11744
rect 11572 11704 11578 11716
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 13078 11744 13084 11756
rect 12391 11716 13084 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 15856 11744 15884 11784
rect 17052 11753 17080 11784
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 17313 11815 17371 11821
rect 17313 11781 17325 11815
rect 17359 11812 17371 11815
rect 17494 11812 17500 11824
rect 17359 11784 17500 11812
rect 17359 11781 17371 11784
rect 17313 11775 17371 11781
rect 17494 11772 17500 11784
rect 17552 11772 17558 11824
rect 13495 11716 15884 11744
rect 15933 11747 15991 11753
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 17037 11747 17095 11753
rect 15979 11716 16896 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 5859 11648 6914 11676
rect 9309 11679 9367 11685
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 10594 11676 10600 11688
rect 9355 11648 10600 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12584 11648 13277 11676
rect 12584 11636 12590 11648
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 13354 11676 13360 11688
rect 13311 11648 13360 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 13464 11608 13492 11707
rect 16868 11617 16896 11716
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17126 11704 17132 11756
rect 17184 11744 17190 11756
rect 17184 11716 17229 11744
rect 17184 11704 17190 11716
rect 23750 11704 23756 11756
rect 23808 11744 23814 11756
rect 24581 11747 24639 11753
rect 24581 11744 24593 11747
rect 23808 11716 24593 11744
rect 23808 11704 23814 11716
rect 24581 11713 24593 11716
rect 24627 11713 24639 11747
rect 28920 11744 28948 11840
rect 29914 11812 29920 11824
rect 29875 11784 29920 11812
rect 29914 11772 29920 11784
rect 29972 11772 29978 11824
rect 30466 11772 30472 11824
rect 30524 11812 30530 11824
rect 30837 11815 30895 11821
rect 30837 11812 30849 11815
rect 30524 11784 30849 11812
rect 30524 11772 30530 11784
rect 30837 11781 30849 11784
rect 30883 11781 30895 11815
rect 30837 11775 30895 11781
rect 31021 11815 31079 11821
rect 31021 11781 31033 11815
rect 31067 11812 31079 11815
rect 33134 11812 33140 11824
rect 31067 11784 33140 11812
rect 31067 11781 31079 11784
rect 31021 11775 31079 11781
rect 33134 11772 33140 11784
rect 33192 11772 33198 11824
rect 29178 11744 29184 11756
rect 28920 11716 29184 11744
rect 24581 11707 24639 11713
rect 29178 11704 29184 11716
rect 29236 11744 29242 11756
rect 29365 11747 29423 11753
rect 29365 11744 29377 11747
rect 29236 11716 29377 11744
rect 29236 11704 29242 11716
rect 29365 11713 29377 11716
rect 29411 11713 29423 11747
rect 29365 11707 29423 11713
rect 29457 11747 29515 11753
rect 29457 11713 29469 11747
rect 29503 11744 29515 11747
rect 29546 11744 29552 11756
rect 29503 11716 29552 11744
rect 29503 11713 29515 11716
rect 29457 11707 29515 11713
rect 29546 11704 29552 11716
rect 29604 11704 29610 11756
rect 29641 11747 29699 11753
rect 29641 11713 29653 11747
rect 29687 11713 29699 11747
rect 29641 11707 29699 11713
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11676 24915 11679
rect 27338 11676 27344 11688
rect 24903 11648 27344 11676
rect 24903 11645 24915 11648
rect 24857 11639 24915 11645
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 28810 11636 28816 11688
rect 28868 11676 28874 11688
rect 29656 11676 29684 11707
rect 28868 11648 29684 11676
rect 28868 11636 28874 11648
rect 16853 11611 16911 11617
rect 13280 11580 13492 11608
rect 13556 11580 16344 11608
rect 13280 11552 13308 11580
rect 13262 11500 13268 11552
rect 13320 11500 13326 11552
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11540 13510 11552
rect 13556 11540 13584 11580
rect 13504 11512 13584 11540
rect 13633 11543 13691 11549
rect 13504 11500 13510 11512
rect 13633 11509 13645 11543
rect 13679 11540 13691 11543
rect 14090 11540 14096 11552
rect 13679 11512 14096 11540
rect 13679 11509 13691 11512
rect 13633 11503 13691 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 16117 11543 16175 11549
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 16206 11540 16212 11552
rect 16163 11512 16212 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16316 11540 16344 11580
rect 16853 11577 16865 11611
rect 16899 11577 16911 11611
rect 16853 11571 16911 11577
rect 29638 11568 29644 11620
rect 29696 11608 29702 11620
rect 29748 11608 29776 11707
rect 30282 11704 30288 11756
rect 30340 11744 30346 11756
rect 30653 11747 30711 11753
rect 30653 11744 30665 11747
rect 30340 11716 30665 11744
rect 30340 11704 30346 11716
rect 30653 11713 30665 11716
rect 30699 11713 30711 11747
rect 32585 11747 32643 11753
rect 32585 11744 32597 11747
rect 30653 11707 30711 11713
rect 30760 11716 32597 11744
rect 30098 11636 30104 11688
rect 30156 11676 30162 11688
rect 30760 11676 30788 11716
rect 32585 11713 32597 11716
rect 32631 11713 32643 11747
rect 33244 11744 33272 11843
rect 33410 11840 33416 11892
rect 33468 11880 33474 11892
rect 34422 11880 34428 11892
rect 33468 11852 34428 11880
rect 33468 11840 33474 11852
rect 34422 11840 34428 11852
rect 34480 11880 34486 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 34480 11852 35173 11880
rect 34480 11840 34486 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 35161 11843 35219 11849
rect 33686 11772 33692 11824
rect 33744 11812 33750 11824
rect 34026 11815 34084 11821
rect 34026 11812 34038 11815
rect 33744 11784 34038 11812
rect 33744 11772 33750 11784
rect 34026 11781 34038 11784
rect 34072 11781 34084 11815
rect 34026 11775 34084 11781
rect 33781 11747 33839 11753
rect 33781 11744 33793 11747
rect 33244 11716 33793 11744
rect 32585 11707 32643 11713
rect 33781 11713 33793 11716
rect 33827 11713 33839 11747
rect 33781 11707 33839 11713
rect 33502 11676 33508 11688
rect 30156 11648 30788 11676
rect 31726 11648 33508 11676
rect 30156 11636 30162 11648
rect 31726 11608 31754 11648
rect 33502 11636 33508 11648
rect 33560 11636 33566 11688
rect 29696 11580 31754 11608
rect 29696 11568 29702 11580
rect 17034 11540 17040 11552
rect 16316 11512 17040 11540
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 20349 11543 20407 11549
rect 20349 11540 20361 11543
rect 20220 11512 20361 11540
rect 20220 11500 20226 11512
rect 20349 11509 20361 11512
rect 20395 11540 20407 11543
rect 20806 11540 20812 11552
rect 20395 11512 20812 11540
rect 20395 11509 20407 11512
rect 20349 11503 20407 11509
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 28350 11500 28356 11552
rect 28408 11540 28414 11552
rect 28810 11540 28816 11552
rect 28408 11512 28816 11540
rect 28408 11500 28414 11512
rect 28810 11500 28816 11512
rect 28868 11500 28874 11552
rect 32674 11540 32680 11552
rect 32635 11512 32680 11540
rect 32674 11500 32680 11512
rect 32732 11500 32738 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 3970 11336 3976 11348
rect 3931 11308 3976 11336
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4890 11336 4896 11348
rect 4295 11308 4896 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5718 11336 5724 11348
rect 5592 11308 5724 11336
rect 5592 11296 5598 11308
rect 5718 11296 5724 11308
rect 5776 11336 5782 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 5776 11308 6837 11336
rect 5776 11296 5782 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 8202 11336 8208 11348
rect 7607 11308 8208 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 10594 11336 10600 11348
rect 10555 11308 10600 11336
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 13446 11336 13452 11348
rect 13407 11308 13452 11336
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 19334 11336 19340 11348
rect 19295 11308 19340 11336
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20622 11336 20628 11348
rect 20535 11308 20628 11336
rect 20622 11296 20628 11308
rect 20680 11336 20686 11348
rect 21450 11336 21456 11348
rect 20680 11308 21456 11336
rect 20680 11296 20686 11308
rect 21450 11296 21456 11308
rect 21508 11336 21514 11348
rect 21637 11339 21695 11345
rect 21637 11336 21649 11339
rect 21508 11308 21649 11336
rect 21508 11296 21514 11308
rect 21637 11305 21649 11308
rect 21683 11305 21695 11339
rect 29546 11336 29552 11348
rect 29507 11308 29552 11336
rect 21637 11299 21695 11305
rect 29546 11296 29552 11308
rect 29604 11296 29610 11348
rect 30466 11336 30472 11348
rect 30427 11308 30472 11336
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 34422 11296 34428 11348
rect 34480 11336 34486 11348
rect 34480 11308 35296 11336
rect 34480 11296 34486 11308
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 8754 11268 8760 11280
rect 3476 11240 8760 11268
rect 3476 11228 3482 11240
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 9766 11228 9772 11280
rect 9824 11268 9830 11280
rect 19889 11271 19947 11277
rect 19889 11268 19901 11271
rect 9824 11240 19901 11268
rect 9824 11228 9830 11240
rect 19889 11237 19901 11240
rect 19935 11268 19947 11271
rect 19978 11268 19984 11280
rect 19935 11240 19984 11268
rect 19935 11237 19947 11240
rect 19889 11231 19947 11237
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 27065 11271 27123 11277
rect 27065 11237 27077 11271
rect 27111 11268 27123 11271
rect 27430 11268 27436 11280
rect 27111 11240 27436 11268
rect 27111 11237 27123 11240
rect 27065 11231 27123 11237
rect 27430 11228 27436 11240
rect 27488 11268 27494 11280
rect 27488 11240 35204 11268
rect 27488 11228 27494 11240
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 12250 11200 12256 11212
rect 4212 11172 7420 11200
rect 12211 11172 12256 11200
rect 4212 11160 4218 11172
rect 7392 11144 7420 11172
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 13354 11200 13360 11212
rect 13315 11172 13360 11200
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 16206 11200 16212 11212
rect 16167 11172 16212 11200
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 16666 11200 16672 11212
rect 16627 11172 16672 11200
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 18874 11160 18880 11212
rect 18932 11200 18938 11212
rect 20530 11200 20536 11212
rect 18932 11172 20536 11200
rect 18932 11160 18938 11172
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 22186 11200 22192 11212
rect 22147 11172 22192 11200
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 29270 11160 29276 11212
rect 29328 11200 29334 11212
rect 29917 11203 29975 11209
rect 29917 11200 29929 11203
rect 29328 11172 29929 11200
rect 29328 11160 29334 11172
rect 29917 11169 29929 11172
rect 29963 11200 29975 11203
rect 32398 11200 32404 11212
rect 29963 11172 32404 11200
rect 29963 11169 29975 11172
rect 29917 11163 29975 11169
rect 32398 11160 32404 11172
rect 32456 11160 32462 11212
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4706 11132 4712 11144
rect 4111 11104 4712 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 5258 11132 5264 11144
rect 5219 11104 5264 11132
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 5500 11104 5549 11132
rect 5500 11092 5506 11104
rect 5537 11101 5549 11104
rect 5583 11132 5595 11135
rect 5902 11132 5908 11144
rect 5583 11104 5908 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6822 11132 6828 11144
rect 6687 11104 6828 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 7374 11132 7380 11144
rect 7335 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 8260 11104 8401 11132
rect 8260 11092 8266 11104
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 11790 11132 11796 11144
rect 10827 11104 11796 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11974 11132 11980 11144
rect 11935 11104 11980 11132
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13538 11132 13544 11144
rect 13499 11104 13544 11132
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 14090 11132 14096 11144
rect 14051 11104 14096 11132
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 16025 11135 16083 11141
rect 16025 11132 16037 11135
rect 15611 11104 16037 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 16025 11101 16037 11104
rect 16071 11101 16083 11135
rect 18506 11132 18512 11144
rect 18467 11104 18512 11132
rect 16025 11095 16083 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11132 22523 11135
rect 24670 11132 24676 11144
rect 22511 11104 24676 11132
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11132 25283 11135
rect 25314 11132 25320 11144
rect 25271 11104 25320 11132
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 25314 11092 25320 11104
rect 25372 11132 25378 11144
rect 25685 11135 25743 11141
rect 25685 11132 25697 11135
rect 25372 11104 25697 11132
rect 25372 11092 25378 11104
rect 25685 11101 25697 11104
rect 25731 11101 25743 11135
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 25685 11095 25743 11101
rect 29288 11104 29745 11132
rect 29288 11076 29316 11104
rect 29733 11101 29745 11104
rect 29779 11132 29791 11135
rect 30282 11132 30288 11144
rect 29779 11104 30288 11132
rect 29779 11101 29791 11104
rect 29733 11095 29791 11101
rect 30282 11092 30288 11104
rect 30340 11092 30346 11144
rect 34882 11132 34888 11144
rect 34843 11104 34888 11132
rect 34882 11092 34888 11104
rect 34940 11092 34946 11144
rect 35176 11141 35204 11240
rect 35268 11141 35296 11308
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11101 35035 11135
rect 34977 11095 35035 11101
rect 35161 11135 35219 11141
rect 35161 11101 35173 11135
rect 35207 11101 35219 11135
rect 35161 11095 35219 11101
rect 35253 11135 35311 11141
rect 35253 11101 35265 11135
rect 35299 11101 35311 11135
rect 35253 11095 35311 11101
rect 3789 11067 3847 11073
rect 3789 11033 3801 11067
rect 3835 11064 3847 11067
rect 5166 11064 5172 11076
rect 3835 11036 5172 11064
rect 3835 11033 3847 11036
rect 3789 11027 3847 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 25952 11067 26010 11073
rect 25952 11033 25964 11067
rect 25998 11064 26010 11067
rect 26970 11064 26976 11076
rect 25998 11036 26976 11064
rect 25998 11033 26010 11036
rect 25952 11027 26010 11033
rect 26970 11024 26976 11036
rect 27028 11024 27034 11076
rect 29270 11024 29276 11076
rect 29328 11024 29334 11076
rect 34146 11024 34152 11076
rect 34204 11064 34210 11076
rect 34701 11067 34759 11073
rect 34701 11064 34713 11067
rect 34204 11036 34713 11064
rect 34204 11024 34210 11036
rect 34701 11033 34713 11036
rect 34747 11033 34759 11067
rect 34992 11064 35020 11095
rect 35894 11092 35900 11144
rect 35952 11132 35958 11144
rect 36081 11135 36139 11141
rect 35952 11104 35997 11132
rect 35952 11092 35958 11104
rect 36081 11101 36093 11135
rect 36127 11101 36139 11135
rect 36081 11095 36139 11101
rect 35713 11067 35771 11073
rect 35713 11064 35725 11067
rect 34992 11036 35725 11064
rect 34701 11027 34759 11033
rect 35713 11033 35725 11036
rect 35759 11033 35771 11067
rect 35713 11027 35771 11033
rect 35802 11024 35808 11076
rect 35860 11064 35866 11076
rect 36096 11064 36124 11095
rect 35860 11036 36124 11064
rect 35860 11024 35866 11036
rect 8202 10996 8208 11008
rect 8163 10968 8208 10996
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 13078 10996 13084 11008
rect 13039 10968 13084 10996
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 14274 10996 14280 11008
rect 14235 10968 14280 10996
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 18322 10996 18328 11008
rect 18283 10968 18328 10996
rect 18322 10956 18328 10968
rect 18380 10956 18386 11008
rect 20806 10956 20812 11008
rect 20864 10996 20870 11008
rect 21085 10999 21143 11005
rect 21085 10996 21097 10999
rect 20864 10968 21097 10996
rect 20864 10956 20870 10968
rect 21085 10965 21097 10968
rect 21131 10965 21143 10999
rect 21085 10959 21143 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 3605 10795 3663 10801
rect 3605 10761 3617 10795
rect 3651 10792 3663 10795
rect 4154 10792 4160 10804
rect 3651 10764 4160 10792
rect 3651 10761 3663 10764
rect 3605 10755 3663 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 6454 10792 6460 10804
rect 5399 10764 6460 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 6822 10752 6828 10804
rect 6880 10792 6886 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 6880 10764 7113 10792
rect 6880 10752 6886 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10792 8079 10795
rect 8110 10792 8116 10804
rect 8067 10764 8116 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 22094 10792 22100 10804
rect 12406 10764 22100 10792
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 12406 10724 12434 10764
rect 22094 10752 22100 10764
rect 22152 10792 22158 10804
rect 24578 10792 24584 10804
rect 22152 10764 24584 10792
rect 22152 10752 22158 10764
rect 24578 10752 24584 10764
rect 24636 10752 24642 10804
rect 26970 10792 26976 10804
rect 26931 10764 26976 10792
rect 26970 10752 26976 10764
rect 27028 10752 27034 10804
rect 27341 10795 27399 10801
rect 27341 10761 27353 10795
rect 27387 10792 27399 10795
rect 27430 10792 27436 10804
rect 27387 10764 27436 10792
rect 27387 10761 27399 10764
rect 27341 10755 27399 10761
rect 27430 10752 27436 10764
rect 27488 10752 27494 10804
rect 29730 10752 29736 10804
rect 29788 10792 29794 10804
rect 30282 10792 30288 10804
rect 29788 10764 30288 10792
rect 29788 10752 29794 10764
rect 30282 10752 30288 10764
rect 30340 10792 30346 10804
rect 30561 10795 30619 10801
rect 30561 10792 30573 10795
rect 30340 10764 30573 10792
rect 30340 10752 30346 10764
rect 30561 10761 30573 10764
rect 30607 10761 30619 10795
rect 30561 10755 30619 10761
rect 33226 10752 33232 10804
rect 33284 10792 33290 10804
rect 33597 10795 33655 10801
rect 33597 10792 33609 10795
rect 33284 10764 33609 10792
rect 33284 10752 33290 10764
rect 33597 10761 33609 10764
rect 33643 10792 33655 10795
rect 33643 10764 34284 10792
rect 33643 10761 33655 10764
rect 33597 10755 33655 10761
rect 3292 10696 12434 10724
rect 17405 10727 17463 10733
rect 3292 10684 3298 10696
rect 17405 10693 17417 10727
rect 17451 10724 17463 10727
rect 18322 10724 18328 10736
rect 17451 10696 18328 10724
rect 17451 10693 17463 10696
rect 17405 10687 17463 10693
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 19058 10724 19064 10736
rect 19019 10696 19064 10724
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 19889 10727 19947 10733
rect 19889 10693 19901 10727
rect 19935 10724 19947 10727
rect 20254 10724 20260 10736
rect 19935 10696 20260 10724
rect 19935 10693 19947 10696
rect 19889 10687 19947 10693
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 24670 10724 24676 10736
rect 20916 10696 22416 10724
rect 24631 10696 24676 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10656 1458 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 1452 10628 2053 10656
rect 1452 10616 1458 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 3142 10656 3148 10668
rect 3103 10628 3148 10656
rect 2041 10619 2099 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3421 10659 3479 10665
rect 3421 10656 3433 10659
rect 3384 10628 3433 10656
rect 3384 10616 3390 10628
rect 3421 10625 3433 10628
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4614 10656 4620 10668
rect 4479 10628 4620 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5169 10659 5227 10665
rect 5169 10656 5181 10659
rect 5132 10628 5181 10656
rect 5132 10616 5138 10628
rect 5169 10625 5181 10628
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 6730 10656 6736 10668
rect 6411 10628 6736 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 19392 10628 19533 10656
rect 19392 10616 19398 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 19978 10656 19984 10668
rect 19751 10628 19984 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 3108 10560 3249 10588
rect 3108 10548 3114 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 17218 10588 17224 10600
rect 17179 10560 17224 10588
rect 3237 10551 3295 10557
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 20916 10597 20944 10696
rect 20990 10616 20996 10668
rect 21048 10656 21054 10668
rect 22388 10665 22416 10696
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 25038 10684 25044 10736
rect 25096 10724 25102 10736
rect 28721 10727 28779 10733
rect 28721 10724 28733 10727
rect 25096 10696 28733 10724
rect 25096 10684 25102 10696
rect 28721 10693 28733 10696
rect 28767 10693 28779 10727
rect 28721 10687 28779 10693
rect 28905 10727 28963 10733
rect 28905 10693 28917 10727
rect 28951 10724 28963 10727
rect 29086 10724 29092 10736
rect 28951 10696 29092 10724
rect 28951 10693 28963 10696
rect 28905 10687 28963 10693
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 29638 10724 29644 10736
rect 29599 10696 29644 10724
rect 29638 10684 29644 10696
rect 29696 10684 29702 10736
rect 34256 10733 34284 10764
rect 34882 10752 34888 10804
rect 34940 10792 34946 10804
rect 35069 10795 35127 10801
rect 35069 10792 35081 10795
rect 34940 10764 35081 10792
rect 34940 10752 34946 10764
rect 35069 10761 35081 10764
rect 35115 10761 35127 10795
rect 35069 10755 35127 10761
rect 34241 10727 34299 10733
rect 34241 10693 34253 10727
rect 34287 10693 34299 10727
rect 35894 10724 35900 10736
rect 34241 10687 34299 10693
rect 35084 10696 35900 10724
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21048 10628 22017 10656
rect 21048 10616 21054 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10625 22431 10659
rect 27154 10656 27160 10668
rect 27115 10628 27160 10656
rect 22373 10619 22431 10625
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20680 10560 20913 10588
rect 20680 10548 20686 10560
rect 20901 10557 20913 10560
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 21821 10591 21879 10597
rect 21821 10557 21833 10591
rect 21867 10557 21879 10591
rect 21821 10551 21879 10557
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 6549 10523 6607 10529
rect 6549 10520 6561 10523
rect 6328 10492 6561 10520
rect 6328 10480 6334 10492
rect 6549 10489 6561 10492
rect 6595 10489 6607 10523
rect 21836 10520 21864 10551
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 22112 10588 22140 10619
rect 27154 10616 27160 10628
rect 27212 10616 27218 10668
rect 27430 10656 27436 10668
rect 27391 10628 27436 10656
rect 27430 10616 27436 10628
rect 27488 10616 27494 10668
rect 29362 10616 29368 10668
rect 29420 10656 29426 10668
rect 35084 10665 35112 10696
rect 35894 10684 35900 10696
rect 35952 10684 35958 10736
rect 29457 10659 29515 10665
rect 29457 10656 29469 10659
rect 29420 10628 29469 10656
rect 29420 10616 29426 10628
rect 29457 10625 29469 10628
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 35069 10659 35127 10665
rect 35069 10625 35081 10659
rect 35115 10625 35127 10659
rect 35069 10619 35127 10625
rect 35253 10659 35311 10665
rect 35253 10625 35265 10659
rect 35299 10656 35311 10659
rect 35802 10656 35808 10668
rect 35299 10628 35808 10656
rect 35299 10625 35311 10628
rect 35253 10619 35311 10625
rect 35802 10616 35808 10628
rect 35860 10616 35866 10668
rect 21968 10560 22140 10588
rect 24397 10591 24455 10597
rect 21968 10548 21974 10560
rect 24397 10557 24409 10591
rect 24443 10588 24455 10591
rect 24578 10588 24584 10600
rect 24443 10560 24584 10588
rect 24443 10557 24455 10560
rect 24397 10551 24455 10557
rect 24578 10548 24584 10560
rect 24636 10548 24642 10600
rect 24857 10591 24915 10597
rect 24857 10557 24869 10591
rect 24903 10588 24915 10591
rect 30190 10588 30196 10600
rect 24903 10560 30196 10588
rect 24903 10557 24915 10560
rect 24857 10551 24915 10557
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 34517 10591 34575 10597
rect 34517 10557 34529 10591
rect 34563 10588 34575 10591
rect 34790 10588 34796 10600
rect 34563 10560 34796 10588
rect 34563 10557 34575 10560
rect 34517 10551 34575 10557
rect 34790 10548 34796 10560
rect 34848 10588 34854 10600
rect 35710 10588 35716 10600
rect 34848 10560 35716 10588
rect 34848 10548 34854 10560
rect 35710 10548 35716 10560
rect 35768 10548 35774 10600
rect 26418 10520 26424 10532
rect 21836 10492 26424 10520
rect 6549 10483 6607 10489
rect 26418 10480 26424 10492
rect 26476 10480 26482 10532
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 2406 10452 2412 10464
rect 1627 10424 2412 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 3016 10424 3157 10452
rect 3016 10412 3022 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 10410 10452 10416 10464
rect 10371 10424 10416 10452
rect 3145 10415 3203 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12492 10424 12909 10452
rect 12492 10412 12498 10424
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 13725 10455 13783 10461
rect 13725 10421 13737 10455
rect 13771 10452 13783 10455
rect 14090 10452 14096 10464
rect 13771 10424 14096 10452
rect 13771 10421 13783 10424
rect 13725 10415 13783 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 20714 10412 20720 10464
rect 20772 10452 20778 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20772 10424 20821 10452
rect 20772 10412 20778 10424
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 20809 10415 20867 10421
rect 21177 10455 21235 10461
rect 21177 10421 21189 10455
rect 21223 10452 21235 10455
rect 27982 10452 27988 10464
rect 21223 10424 27988 10452
rect 21223 10421 21235 10424
rect 21177 10415 21235 10421
rect 27982 10412 27988 10424
rect 28040 10412 28046 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2958 10248 2964 10260
rect 2919 10220 2964 10248
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 5258 10248 5264 10260
rect 4448 10220 5264 10248
rect 2777 10183 2835 10189
rect 2777 10149 2789 10183
rect 2823 10180 2835 10183
rect 4448 10180 4476 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6822 10248 6828 10260
rect 6043 10220 6828 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 17276 10220 17325 10248
rect 17276 10208 17282 10220
rect 17313 10217 17325 10220
rect 17359 10217 17371 10251
rect 17313 10211 17371 10217
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20809 10251 20867 10257
rect 20809 10248 20821 10251
rect 20588 10220 20821 10248
rect 20588 10208 20594 10220
rect 20809 10217 20821 10220
rect 20855 10217 20867 10251
rect 20809 10211 20867 10217
rect 27430 10208 27436 10260
rect 27488 10248 27494 10260
rect 28169 10251 28227 10257
rect 28169 10248 28181 10251
rect 27488 10220 28181 10248
rect 27488 10208 27494 10220
rect 28169 10217 28181 10220
rect 28215 10217 28227 10251
rect 28169 10211 28227 10217
rect 29454 10208 29460 10260
rect 29512 10248 29518 10260
rect 29730 10248 29736 10260
rect 29512 10220 29736 10248
rect 29512 10208 29518 10220
rect 29730 10208 29736 10220
rect 29788 10208 29794 10260
rect 2823 10152 4476 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 4798 10140 4804 10192
rect 4856 10140 4862 10192
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10180 6699 10183
rect 6730 10180 6736 10192
rect 6687 10152 6736 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 6730 10140 6736 10152
rect 6788 10180 6794 10192
rect 14366 10180 14372 10192
rect 6788 10152 14372 10180
rect 6788 10140 6794 10152
rect 14366 10140 14372 10152
rect 14424 10180 14430 10192
rect 18598 10180 18604 10192
rect 14424 10152 18604 10180
rect 14424 10140 14430 10152
rect 18598 10140 18604 10152
rect 18656 10180 18662 10192
rect 19521 10183 19579 10189
rect 19521 10180 19533 10183
rect 18656 10152 19533 10180
rect 18656 10140 18662 10152
rect 19521 10149 19533 10152
rect 19567 10149 19579 10183
rect 19521 10143 19579 10149
rect 20257 10183 20315 10189
rect 20257 10149 20269 10183
rect 20303 10149 20315 10183
rect 20257 10143 20315 10149
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4816 10112 4844 10140
rect 5626 10112 5632 10124
rect 4571 10084 5632 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 14090 10112 14096 10124
rect 5960 10084 12434 10112
rect 14051 10084 14096 10112
rect 5960 10072 5966 10084
rect 2222 10004 2228 10056
rect 2280 10044 2286 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2280 10016 2973 10044
rect 2280 10004 2286 10016
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 3050 10004 3056 10056
rect 3108 10044 3114 10056
rect 4801 10047 4859 10053
rect 3108 10016 3153 10044
rect 3108 10004 3114 10016
rect 4801 10013 4813 10047
rect 4847 10044 4859 10047
rect 5166 10044 5172 10056
rect 4847 10016 5172 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5592 10016 5825 10044
rect 5592 10004 5598 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 7466 10044 7472 10056
rect 6328 10016 7472 10044
rect 6328 10004 6334 10016
rect 7466 10004 7472 10016
rect 7524 10044 7530 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7524 10016 7665 10044
rect 7524 10004 7530 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 10410 10044 10416 10056
rect 10371 10016 10416 10044
rect 7653 10007 7711 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11882 10004 11888 10056
rect 11940 10044 11946 10056
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 11940 10016 12265 10044
rect 11940 10004 11946 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 3142 9936 3148 9988
rect 3200 9976 3206 9988
rect 3237 9979 3295 9985
rect 3237 9976 3249 9979
rect 3200 9948 3249 9976
rect 3200 9936 3206 9948
rect 3237 9945 3249 9948
rect 3283 9976 3295 9979
rect 4246 9976 4252 9988
rect 3283 9948 4252 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 7837 9979 7895 9985
rect 7837 9945 7849 9979
rect 7883 9976 7895 9979
rect 8846 9976 8852 9988
rect 7883 9948 8852 9976
rect 7883 9945 7895 9948
rect 7837 9939 7895 9945
rect 8846 9936 8852 9948
rect 8904 9936 8910 9988
rect 10597 9979 10655 9985
rect 10597 9945 10609 9979
rect 10643 9976 10655 9979
rect 11974 9976 11980 9988
rect 10643 9948 11980 9976
rect 10643 9945 10655 9948
rect 10597 9939 10655 9945
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 12406 9976 12434 10084
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 14274 10112 14280 10124
rect 14235 10084 14280 10112
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 15930 10112 15936 10124
rect 15891 10084 15936 10112
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 19334 10044 19340 10056
rect 18524 10016 19340 10044
rect 18524 9976 18552 10016
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19536 10044 19564 10143
rect 20272 10112 20300 10143
rect 20714 10140 20720 10192
rect 20772 10180 20778 10192
rect 21542 10180 21548 10192
rect 20772 10152 21548 10180
rect 20772 10140 20778 10152
rect 21542 10140 21548 10152
rect 21600 10180 21606 10192
rect 21729 10183 21787 10189
rect 21729 10180 21741 10183
rect 21600 10152 21741 10180
rect 21600 10140 21606 10152
rect 21729 10149 21741 10152
rect 21775 10180 21787 10183
rect 21910 10180 21916 10192
rect 21775 10152 21916 10180
rect 21775 10149 21787 10152
rect 21729 10143 21787 10149
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 29638 10140 29644 10192
rect 29696 10140 29702 10192
rect 20622 10112 20628 10124
rect 20272 10084 20628 10112
rect 20622 10072 20628 10084
rect 20680 10112 20686 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20680 10084 20913 10112
rect 20680 10072 20686 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 27338 10112 27344 10124
rect 27299 10084 27344 10112
rect 20901 10075 20959 10081
rect 27338 10072 27344 10084
rect 27396 10072 27402 10124
rect 29656 10112 29684 10140
rect 29656 10084 29960 10112
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 19536 10016 20085 10044
rect 20073 10013 20085 10016
rect 20119 10013 20131 10047
rect 20806 10044 20812 10056
rect 20719 10016 20812 10044
rect 20073 10007 20131 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 22278 10044 22284 10056
rect 22239 10016 22284 10044
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 23106 10044 23112 10056
rect 23067 10016 23112 10044
rect 23106 10004 23112 10016
rect 23164 10004 23170 10056
rect 27522 10004 27528 10056
rect 27580 10044 27586 10056
rect 29454 10044 29460 10056
rect 27580 10016 29460 10044
rect 27580 10004 27586 10016
rect 29454 10004 29460 10016
rect 29512 10004 29518 10056
rect 29638 10044 29644 10056
rect 29599 10016 29644 10044
rect 29638 10004 29644 10016
rect 29696 10004 29702 10056
rect 29822 10044 29828 10056
rect 29783 10016 29828 10044
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 29932 10053 29960 10084
rect 30282 10072 30288 10124
rect 30340 10112 30346 10124
rect 30745 10115 30803 10121
rect 30745 10112 30757 10115
rect 30340 10084 30757 10112
rect 30340 10072 30346 10084
rect 30745 10081 30757 10084
rect 30791 10081 30803 10115
rect 30745 10075 30803 10081
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30009 10047 30067 10053
rect 30009 10013 30021 10047
rect 30055 10013 30067 10047
rect 38102 10044 38108 10056
rect 38063 10016 38108 10044
rect 30009 10007 30067 10013
rect 20824 9976 20852 10004
rect 25682 9976 25688 9988
rect 12406 9948 18552 9976
rect 18616 9948 20852 9976
rect 25643 9948 25688 9976
rect 16485 9911 16543 9917
rect 16485 9877 16497 9911
rect 16531 9908 16543 9911
rect 16574 9908 16580 9920
rect 16531 9880 16580 9908
rect 16531 9877 16543 9880
rect 16485 9871 16543 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 18616 9917 18644 9948
rect 25682 9936 25688 9948
rect 25740 9936 25746 9988
rect 27982 9936 27988 9988
rect 28040 9976 28046 9988
rect 28077 9979 28135 9985
rect 28077 9976 28089 9979
rect 28040 9948 28089 9976
rect 28040 9936 28046 9948
rect 28077 9945 28089 9948
rect 28123 9976 28135 9979
rect 29270 9976 29276 9988
rect 28123 9948 29276 9976
rect 28123 9945 28135 9948
rect 28077 9939 28135 9945
rect 29270 9936 29276 9948
rect 29328 9936 29334 9988
rect 29472 9976 29500 10004
rect 30024 9976 30052 10007
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 29472 9948 30052 9976
rect 30742 9936 30748 9988
rect 30800 9976 30806 9988
rect 30990 9979 31048 9985
rect 30990 9976 31002 9979
rect 30800 9948 31002 9976
rect 30800 9936 30806 9948
rect 30990 9945 31002 9948
rect 31036 9945 31048 9979
rect 30990 9939 31048 9945
rect 18601 9911 18659 9917
rect 18601 9908 18613 9911
rect 18564 9880 18613 9908
rect 18564 9868 18570 9880
rect 18601 9877 18613 9880
rect 18647 9877 18659 9911
rect 21174 9908 21180 9920
rect 21135 9880 21180 9908
rect 18601 9871 18659 9877
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 22465 9911 22523 9917
rect 22465 9877 22477 9911
rect 22511 9908 22523 9911
rect 22830 9908 22836 9920
rect 22511 9880 22836 9908
rect 22511 9877 22523 9880
rect 22465 9871 22523 9877
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 30285 9911 30343 9917
rect 22980 9880 23025 9908
rect 22980 9868 22986 9880
rect 30285 9877 30297 9911
rect 30331 9908 30343 9911
rect 30650 9908 30656 9920
rect 30331 9880 30656 9908
rect 30331 9877 30343 9880
rect 30285 9871 30343 9877
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 32122 9908 32128 9920
rect 32083 9880 32128 9908
rect 32122 9868 32128 9880
rect 32180 9868 32186 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 10778 9704 10784 9716
rect 3476 9676 10784 9704
rect 3476 9664 3482 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 17678 9704 17684 9716
rect 16632 9676 17684 9704
rect 16632 9664 16638 9676
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 4246 9636 4252 9648
rect 3016 9608 3372 9636
rect 4159 9608 4252 9636
rect 3016 9596 3022 9608
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 3145 9571 3203 9577
rect 3145 9568 3157 9571
rect 2363 9540 3157 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 3145 9537 3157 9540
rect 3191 9568 3203 9571
rect 3234 9568 3240 9580
rect 3191 9540 3240 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3344 9577 3372 9608
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4172 9568 4200 9608
rect 4246 9596 4252 9608
rect 4304 9636 4310 9648
rect 4890 9636 4896 9648
rect 4304 9608 4896 9636
rect 4304 9596 4310 9608
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 7282 9636 7288 9648
rect 5684 9608 7288 9636
rect 5684 9596 5690 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7466 9636 7472 9648
rect 7427 9608 7472 9636
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 12537 9636
rect 12492 9596 12498 9608
rect 13998 9596 14004 9648
rect 14056 9636 14062 9648
rect 17604 9645 17632 9676
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 19337 9707 19395 9713
rect 19337 9673 19349 9707
rect 19383 9704 19395 9707
rect 20254 9704 20260 9716
rect 19383 9676 20260 9704
rect 19383 9673 19395 9676
rect 19337 9667 19395 9673
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 20622 9664 20628 9716
rect 20680 9704 20686 9716
rect 20993 9707 21051 9713
rect 20993 9704 21005 9707
rect 20680 9676 21005 9704
rect 20680 9664 20686 9676
rect 20993 9673 21005 9676
rect 21039 9673 21051 9707
rect 20993 9667 21051 9673
rect 26973 9707 27031 9713
rect 26973 9673 26985 9707
rect 27019 9704 27031 9707
rect 27154 9704 27160 9716
rect 27019 9676 27160 9704
rect 27019 9673 27031 9676
rect 26973 9667 27031 9673
rect 27154 9664 27160 9676
rect 27212 9664 27218 9716
rect 29641 9707 29699 9713
rect 29641 9673 29653 9707
rect 29687 9704 29699 9707
rect 29822 9704 29828 9716
rect 29687 9676 29828 9704
rect 29687 9673 29699 9676
rect 29641 9667 29699 9673
rect 29822 9664 29828 9676
rect 29880 9664 29886 9716
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 14056 9608 14105 9636
rect 14056 9596 14062 9608
rect 14093 9605 14105 9608
rect 14139 9605 14151 9639
rect 17589 9639 17647 9645
rect 14093 9599 14151 9605
rect 15948 9608 16988 9636
rect 4111 9540 4200 9568
rect 4801 9571 4859 9577
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5810 9568 5816 9580
rect 4847 9540 5816 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3712 9500 3740 9531
rect 5810 9528 5816 9540
rect 5868 9568 5874 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5868 9540 6377 9568
rect 5868 9528 5874 9540
rect 6365 9537 6377 9540
rect 6411 9568 6423 9571
rect 7484 9568 7512 9596
rect 15654 9568 15660 9580
rect 6411 9540 7512 9568
rect 15615 9540 15660 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 15654 9528 15660 9540
rect 15712 9568 15718 9580
rect 15948 9577 15976 9608
rect 16960 9580 16988 9608
rect 17589 9605 17601 9639
rect 17635 9605 17647 9639
rect 18598 9636 18604 9648
rect 18559 9608 18604 9636
rect 17589 9599 17647 9605
rect 18598 9596 18604 9608
rect 18656 9636 18662 9648
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 18656 9608 19257 9636
rect 18656 9596 18662 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 19245 9599 19303 9605
rect 22097 9639 22155 9645
rect 22097 9605 22109 9639
rect 22143 9636 22155 9639
rect 25038 9636 25044 9648
rect 22143 9608 25044 9636
rect 22143 9605 22155 9608
rect 22097 9599 22155 9605
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 25406 9636 25412 9648
rect 25319 9608 25412 9636
rect 25406 9596 25412 9608
rect 25464 9636 25470 9648
rect 26329 9639 26387 9645
rect 26329 9636 26341 9639
rect 25464 9608 26341 9636
rect 25464 9596 25470 9608
rect 26329 9605 26341 9608
rect 26375 9605 26387 9639
rect 29362 9636 29368 9648
rect 26329 9599 26387 9605
rect 26436 9608 29368 9636
rect 15933 9571 15991 9577
rect 15712 9540 15884 9568
rect 15712 9528 15718 9540
rect 3108 9472 3740 9500
rect 3108 9460 3114 9472
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4982 9500 4988 9512
rect 4212 9472 4988 9500
rect 4212 9460 4218 9472
rect 4982 9460 4988 9472
rect 5040 9500 5046 9512
rect 5077 9503 5135 9509
rect 5077 9500 5089 9503
rect 5040 9472 5089 9500
rect 5040 9460 5046 9472
rect 5077 9469 5089 9472
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12710 9500 12716 9512
rect 12299 9472 12716 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15746 9500 15752 9512
rect 15243 9472 15752 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9432 4307 9435
rect 15102 9432 15108 9444
rect 4295 9404 15108 9432
rect 4295 9401 4307 9404
rect 4249 9395 4307 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 15212 9364 15240 9463
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 15856 9500 15884 9540
rect 15933 9537 15945 9571
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 16669 9571 16727 9577
rect 16669 9537 16681 9571
rect 16715 9537 16727 9571
rect 16942 9568 16948 9580
rect 16903 9540 16948 9568
rect 16669 9531 16727 9537
rect 16574 9500 16580 9512
rect 15856 9472 16580 9500
rect 16574 9460 16580 9472
rect 16632 9500 16638 9512
rect 16684 9500 16712 9531
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 19426 9568 19432 9580
rect 19387 9540 19432 9568
rect 19426 9528 19432 9540
rect 19484 9568 19490 9580
rect 20070 9568 20076 9580
rect 19484 9540 20076 9568
rect 19484 9528 19490 9540
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 16632 9472 16712 9500
rect 16632 9460 16638 9472
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 18138 9500 18144 9512
rect 16908 9472 18144 9500
rect 16908 9460 16914 9472
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19116 9472 19809 9500
rect 19116 9460 19122 9472
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20806 9500 20812 9512
rect 20027 9472 20812 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 22649 9503 22707 9509
rect 22649 9469 22661 9503
rect 22695 9469 22707 9503
rect 22830 9500 22836 9512
rect 22791 9472 22836 9500
rect 22649 9463 22707 9469
rect 15948 9404 16712 9432
rect 15948 9373 15976 9404
rect 16684 9376 16712 9404
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 19392 9404 20453 9432
rect 19392 9392 19398 9404
rect 20441 9401 20453 9404
rect 20487 9432 20499 9435
rect 20714 9432 20720 9444
rect 20487 9404 20720 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 22664 9432 22692 9463
rect 22830 9460 22836 9472
rect 22888 9460 22894 9512
rect 23658 9500 23664 9512
rect 23619 9472 23664 9500
rect 23658 9460 23664 9472
rect 23716 9500 23722 9512
rect 25424 9509 25452 9596
rect 26436 9580 26464 9608
rect 26145 9571 26203 9577
rect 26145 9537 26157 9571
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 25409 9503 25467 9509
rect 25409 9500 25421 9503
rect 23716 9472 25421 9500
rect 23716 9460 23722 9472
rect 25409 9469 25421 9472
rect 25455 9469 25467 9503
rect 26160 9500 26188 9531
rect 26418 9528 26424 9580
rect 26476 9568 26482 9580
rect 27157 9571 27215 9577
rect 26476 9540 26521 9568
rect 26476 9528 26482 9540
rect 27157 9537 27169 9571
rect 27203 9537 27215 9571
rect 27338 9568 27344 9580
rect 27299 9540 27344 9568
rect 27157 9531 27215 9537
rect 26970 9500 26976 9512
rect 26160 9472 26976 9500
rect 25409 9463 25467 9469
rect 26970 9460 26976 9472
rect 27028 9500 27034 9512
rect 27172 9500 27200 9531
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 27448 9577 27476 9608
rect 29362 9596 29368 9608
rect 29420 9636 29426 9648
rect 30101 9639 30159 9645
rect 30101 9636 30113 9639
rect 29420 9608 30113 9636
rect 29420 9596 29426 9608
rect 30101 9605 30113 9608
rect 30147 9605 30159 9639
rect 30101 9599 30159 9605
rect 30190 9596 30196 9648
rect 30248 9636 30254 9648
rect 30285 9639 30343 9645
rect 30285 9636 30297 9639
rect 30248 9608 30297 9636
rect 30248 9596 30254 9608
rect 30285 9605 30297 9608
rect 30331 9636 30343 9639
rect 32122 9636 32128 9648
rect 30331 9608 32128 9636
rect 30331 9605 30343 9608
rect 30285 9599 30343 9605
rect 32122 9596 32128 9608
rect 32180 9596 32186 9648
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 29270 9568 29276 9580
rect 29231 9540 29276 9568
rect 27433 9531 27491 9537
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29457 9571 29515 9577
rect 29457 9537 29469 9571
rect 29503 9568 29515 9571
rect 29546 9568 29552 9580
rect 29503 9540 29552 9568
rect 29503 9537 29515 9540
rect 29457 9531 29515 9537
rect 29546 9528 29552 9540
rect 29604 9528 29610 9580
rect 35434 9528 35440 9580
rect 35492 9568 35498 9580
rect 35601 9571 35659 9577
rect 35601 9568 35613 9571
rect 35492 9540 35613 9568
rect 35492 9528 35498 9540
rect 35601 9537 35613 9540
rect 35647 9537 35659 9571
rect 35601 9531 35659 9537
rect 28537 9503 28595 9509
rect 28537 9500 28549 9503
rect 27028 9472 28549 9500
rect 27028 9460 27034 9472
rect 28537 9469 28549 9472
rect 28583 9500 28595 9503
rect 33226 9500 33232 9512
rect 28583 9472 33232 9500
rect 28583 9469 28595 9472
rect 28537 9463 28595 9469
rect 33226 9460 33232 9472
rect 33284 9460 33290 9512
rect 35342 9500 35348 9512
rect 34808 9472 35348 9500
rect 23382 9432 23388 9444
rect 22664 9404 23388 9432
rect 23382 9392 23388 9404
rect 23440 9392 23446 9444
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 27893 9435 27951 9441
rect 27893 9432 27905 9435
rect 27396 9404 27905 9432
rect 27396 9392 27402 9404
rect 27893 9401 27905 9404
rect 27939 9401 27951 9435
rect 32398 9432 32404 9444
rect 32359 9404 32404 9432
rect 27893 9395 27951 9401
rect 32398 9392 32404 9404
rect 32456 9392 32462 9444
rect 8904 9336 15240 9364
rect 15933 9367 15991 9373
rect 8904 9324 8910 9336
rect 15933 9333 15945 9367
rect 15979 9333 15991 9367
rect 15933 9327 15991 9333
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16574 9364 16580 9376
rect 16163 9336 16580 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 17126 9364 17132 9376
rect 16724 9336 16769 9364
rect 17087 9336 17132 9364
rect 16724 9324 16730 9336
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9364 22063 9367
rect 25314 9364 25320 9376
rect 22051 9336 25320 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 25961 9367 26019 9373
rect 25961 9333 25973 9367
rect 26007 9364 26019 9367
rect 26142 9364 26148 9376
rect 26007 9336 26148 9364
rect 26007 9333 26019 9336
rect 25961 9327 26019 9333
rect 26142 9324 26148 9336
rect 26200 9324 26206 9376
rect 30282 9324 30288 9376
rect 30340 9364 30346 9376
rect 30469 9367 30527 9373
rect 30469 9364 30481 9367
rect 30340 9336 30481 9364
rect 30340 9324 30346 9336
rect 30469 9333 30481 9336
rect 30515 9333 30527 9367
rect 32582 9364 32588 9376
rect 32543 9336 32588 9364
rect 30469 9327 30527 9333
rect 32582 9324 32588 9336
rect 32640 9324 32646 9376
rect 34606 9324 34612 9376
rect 34664 9364 34670 9376
rect 34808 9373 34836 9472
rect 35342 9460 35348 9472
rect 35400 9460 35406 9512
rect 34793 9367 34851 9373
rect 34793 9364 34805 9367
rect 34664 9336 34805 9364
rect 34664 9324 34670 9336
rect 34793 9333 34805 9336
rect 34839 9333 34851 9367
rect 34793 9327 34851 9333
rect 35986 9324 35992 9376
rect 36044 9364 36050 9376
rect 36725 9367 36783 9373
rect 36725 9364 36737 9367
rect 36044 9336 36737 9364
rect 36044 9324 36050 9336
rect 36725 9333 36737 9336
rect 36771 9333 36783 9367
rect 36725 9327 36783 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3050 9160 3056 9172
rect 3007 9132 3056 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5350 9160 5356 9172
rect 4939 9132 5356 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5350 9120 5356 9132
rect 5408 9160 5414 9172
rect 8202 9160 8208 9172
rect 5408 9132 6914 9160
rect 8163 9132 8208 9160
rect 5408 9120 5414 9132
rect 1394 9092 1400 9104
rect 1355 9064 1400 9092
rect 1394 9052 1400 9064
rect 1452 9052 1458 9104
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 5258 9024 5264 9036
rect 4448 8996 5264 9024
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 4448 8965 4476 8996
rect 5258 8984 5264 8996
rect 5316 9024 5322 9036
rect 5534 9024 5540 9036
rect 5316 8996 5540 9024
rect 5316 8984 5322 8996
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 6886 9024 6914 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16577 9163 16635 9169
rect 16577 9160 16589 9163
rect 15804 9132 16589 9160
rect 15804 9120 15810 9132
rect 16577 9129 16589 9132
rect 16623 9160 16635 9163
rect 16850 9160 16856 9172
rect 16623 9132 16856 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 20530 9160 20536 9172
rect 20491 9132 20536 9160
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 26970 9160 26976 9172
rect 26931 9132 26976 9160
rect 26970 9120 26976 9132
rect 27028 9120 27034 9172
rect 28994 9160 29000 9172
rect 28955 9132 29000 9160
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29454 9120 29460 9172
rect 29512 9160 29518 9172
rect 29641 9163 29699 9169
rect 29641 9160 29653 9163
rect 29512 9132 29653 9160
rect 29512 9120 29518 9132
rect 29641 9129 29653 9132
rect 29687 9129 29699 9163
rect 29641 9123 29699 9129
rect 35345 9163 35403 9169
rect 35345 9129 35357 9163
rect 35391 9160 35403 9163
rect 35434 9160 35440 9172
rect 35391 9132 35440 9160
rect 35391 9129 35403 9132
rect 35345 9123 35403 9129
rect 35434 9120 35440 9132
rect 35492 9120 35498 9172
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 19337 9095 19395 9101
rect 19337 9092 19349 9095
rect 15160 9064 19349 9092
rect 15160 9052 15166 9064
rect 19337 9061 19349 9064
rect 19383 9092 19395 9095
rect 19426 9092 19432 9104
rect 19383 9064 19432 9092
rect 19383 9061 19395 9064
rect 19337 9055 19395 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 18506 9024 18512 9036
rect 6886 8996 18512 9024
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 32674 8984 32680 9036
rect 32732 9024 32738 9036
rect 35342 9024 35348 9036
rect 32732 8996 35348 9024
rect 32732 8984 32738 8996
rect 2777 8959 2835 8965
rect 2777 8956 2789 8959
rect 1636 8928 2789 8956
rect 1636 8916 1642 8928
rect 2777 8925 2789 8928
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5074 8956 5080 8968
rect 5031 8928 5080 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8202 8956 8208 8968
rect 7699 8928 8208 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2501 8891 2559 8897
rect 2501 8888 2513 8891
rect 2464 8860 2513 8888
rect 2464 8848 2470 8860
rect 2501 8857 2513 8860
rect 2547 8857 2559 8891
rect 2501 8851 2559 8857
rect 5537 8891 5595 8897
rect 5537 8857 5549 8891
rect 5583 8888 5595 8891
rect 5626 8888 5632 8900
rect 5583 8860 5632 8888
rect 5583 8857 5595 8860
rect 5537 8851 5595 8857
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7668 8888 7696 8919
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 26142 8956 26148 8968
rect 26103 8928 26148 8956
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8956 26479 8959
rect 27430 8956 27436 8968
rect 26467 8928 27436 8956
rect 26467 8925 26479 8928
rect 26421 8919 26479 8925
rect 27430 8916 27436 8928
rect 27488 8916 27494 8968
rect 29086 8916 29092 8968
rect 29144 8956 29150 8968
rect 31021 8959 31079 8965
rect 31021 8956 31033 8959
rect 29144 8928 31033 8956
rect 29144 8916 29150 8928
rect 31021 8925 31033 8928
rect 31067 8956 31079 8959
rect 34606 8956 34612 8968
rect 31067 8928 34612 8956
rect 31067 8925 31079 8928
rect 31021 8919 31079 8925
rect 34606 8916 34612 8928
rect 34664 8916 34670 8968
rect 34716 8965 34744 8996
rect 35342 8984 35348 8996
rect 35400 8984 35406 9036
rect 34701 8959 34759 8965
rect 34701 8925 34713 8959
rect 34747 8925 34759 8959
rect 34882 8956 34888 8968
rect 34843 8928 34888 8956
rect 34701 8919 34759 8925
rect 34882 8916 34888 8928
rect 34940 8916 34946 8968
rect 34977 8959 35035 8965
rect 34977 8925 34989 8959
rect 35023 8925 35035 8959
rect 34977 8919 35035 8925
rect 35069 8959 35127 8965
rect 35069 8925 35081 8959
rect 35115 8956 35127 8959
rect 35894 8956 35900 8968
rect 35115 8928 35900 8956
rect 35115 8925 35127 8928
rect 35069 8919 35127 8925
rect 7340 8860 7696 8888
rect 27448 8888 27476 8916
rect 30466 8888 30472 8900
rect 27448 8860 30472 8888
rect 7340 8848 7346 8860
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 30650 8848 30656 8900
rect 30708 8888 30714 8900
rect 30754 8891 30812 8897
rect 30754 8888 30766 8891
rect 30708 8860 30766 8888
rect 30708 8848 30714 8860
rect 30754 8857 30766 8860
rect 30800 8857 30812 8891
rect 30754 8851 30812 8857
rect 34422 8848 34428 8900
rect 34480 8888 34486 8900
rect 34992 8888 35020 8919
rect 35894 8916 35900 8928
rect 35952 8916 35958 8968
rect 34480 8860 35020 8888
rect 34480 8848 34486 8860
rect 25958 8820 25964 8832
rect 25919 8792 25964 8820
rect 25958 8780 25964 8792
rect 26016 8780 26022 8832
rect 26326 8820 26332 8832
rect 26287 8792 26332 8820
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 28994 8780 29000 8832
rect 29052 8820 29058 8832
rect 35526 8820 35532 8832
rect 29052 8792 35532 8820
rect 29052 8780 29058 8792
rect 35526 8780 35532 8792
rect 35584 8780 35590 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 5810 8616 5816 8628
rect 5771 8588 5816 8616
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 8846 8616 8852 8628
rect 8807 8588 8852 8616
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 9416 8588 10425 8616
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 9416 8557 9444 8588
rect 10413 8585 10425 8588
rect 10459 8616 10471 8619
rect 15654 8616 15660 8628
rect 10459 8588 15660 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 29086 8616 29092 8628
rect 29047 8588 29092 8616
rect 29086 8576 29092 8588
rect 29144 8576 29150 8628
rect 29641 8619 29699 8625
rect 29641 8585 29653 8619
rect 29687 8616 29699 8619
rect 30006 8616 30012 8628
rect 29687 8588 30012 8616
rect 29687 8585 29699 8588
rect 29641 8579 29699 8585
rect 30006 8576 30012 8588
rect 30064 8576 30070 8628
rect 30466 8576 30472 8628
rect 30524 8576 30530 8628
rect 30742 8616 30748 8628
rect 30703 8588 30748 8616
rect 30742 8576 30748 8588
rect 30800 8576 30806 8628
rect 34425 8619 34483 8625
rect 34425 8585 34437 8619
rect 34471 8616 34483 8619
rect 34882 8616 34888 8628
rect 34471 8588 34888 8616
rect 34471 8585 34483 8588
rect 34425 8579 34483 8585
rect 34882 8576 34888 8588
rect 34940 8576 34946 8628
rect 9401 8551 9459 8557
rect 3476 8520 9352 8548
rect 3476 8508 3482 8520
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 5718 8480 5724 8492
rect 4479 8452 5724 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 5868 8452 7205 8480
rect 5868 8440 5874 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7650 8480 7656 8492
rect 7611 8452 7656 8480
rect 7193 8443 7251 8449
rect 7650 8440 7656 8452
rect 7708 8480 7714 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 7708 8452 8309 8480
rect 7708 8440 7714 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 9324 8480 9352 8520
rect 9401 8517 9413 8551
rect 9447 8517 9459 8551
rect 11974 8548 11980 8560
rect 9401 8511 9459 8517
rect 9508 8520 11980 8548
rect 9508 8480 9536 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 22465 8551 22523 8557
rect 22465 8517 22477 8551
rect 22511 8548 22523 8551
rect 22922 8548 22928 8560
rect 22511 8520 22928 8548
rect 22511 8517 22523 8520
rect 22465 8511 22523 8517
rect 22922 8508 22928 8520
rect 22980 8508 22986 8560
rect 24121 8551 24179 8557
rect 24121 8517 24133 8551
rect 24167 8548 24179 8551
rect 24486 8548 24492 8560
rect 24167 8520 24492 8548
rect 24167 8517 24179 8520
rect 24121 8511 24179 8517
rect 24486 8508 24492 8520
rect 24544 8548 24550 8560
rect 28994 8548 29000 8560
rect 24544 8520 29000 8548
rect 24544 8508 24550 8520
rect 28994 8508 29000 8520
rect 29052 8508 29058 8560
rect 30484 8548 30512 8576
rect 30392 8520 30512 8548
rect 9674 8480 9680 8492
rect 9324 8452 9536 8480
rect 9635 8452 9680 8480
rect 8297 8443 8355 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 24302 8440 24308 8492
rect 24360 8480 24366 8492
rect 25593 8483 25651 8489
rect 25593 8480 25605 8483
rect 24360 8452 25605 8480
rect 24360 8440 24366 8452
rect 25593 8449 25605 8452
rect 25639 8449 25651 8483
rect 25593 8443 25651 8449
rect 29638 8440 29644 8492
rect 29696 8480 29702 8492
rect 30098 8480 30104 8492
rect 29696 8452 30104 8480
rect 29696 8440 29702 8452
rect 30098 8440 30104 8452
rect 30156 8440 30162 8492
rect 30282 8480 30288 8492
rect 30243 8452 30288 8480
rect 30282 8440 30288 8452
rect 30340 8440 30346 8492
rect 30392 8489 30420 8520
rect 32582 8508 32588 8560
rect 32640 8548 32646 8560
rect 32640 8520 37320 8548
rect 32640 8508 32646 8520
rect 30377 8483 30435 8489
rect 30377 8449 30389 8483
rect 30423 8449 30435 8483
rect 30377 8443 30435 8449
rect 30469 8483 30527 8489
rect 30469 8449 30481 8483
rect 30515 8449 30527 8483
rect 30469 8443 30527 8449
rect 34701 8483 34759 8489
rect 34701 8449 34713 8483
rect 34747 8480 34759 8483
rect 35894 8480 35900 8492
rect 34747 8452 35900 8480
rect 34747 8449 34759 8452
rect 34701 8443 34759 8449
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8412 6975 8415
rect 8018 8412 8024 8424
rect 6963 8384 8024 8412
rect 6963 8381 6975 8384
rect 6917 8375 6975 8381
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 8904 8384 9505 8412
rect 8904 8372 8910 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 22278 8412 22284 8424
rect 22239 8384 22284 8412
rect 9493 8375 9551 8381
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 25869 8415 25927 8421
rect 25869 8381 25881 8415
rect 25915 8412 25927 8415
rect 27522 8412 27528 8424
rect 25915 8384 27528 8412
rect 25915 8381 25927 8384
rect 25869 8375 25927 8381
rect 27522 8372 27528 8384
rect 27580 8372 27586 8424
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 11054 8344 11060 8356
rect 9907 8316 11060 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 26326 8344 26332 8356
rect 23440 8316 26332 8344
rect 23440 8304 23446 8316
rect 26326 8304 26332 8316
rect 26384 8304 26390 8356
rect 30006 8304 30012 8356
rect 30064 8344 30070 8356
rect 30484 8344 30512 8443
rect 35894 8440 35900 8452
rect 35952 8440 35958 8492
rect 37292 8489 37320 8520
rect 37277 8483 37335 8489
rect 37277 8449 37289 8483
rect 37323 8449 37335 8483
rect 37277 8443 37335 8449
rect 33686 8372 33692 8424
rect 33744 8412 33750 8424
rect 34422 8412 34428 8424
rect 33744 8384 34428 8412
rect 33744 8372 33750 8384
rect 34422 8372 34428 8384
rect 34480 8372 34486 8424
rect 30064 8316 30512 8344
rect 30064 8304 30070 8316
rect 34330 8304 34336 8356
rect 34388 8344 34394 8356
rect 34609 8347 34667 8353
rect 34609 8344 34621 8347
rect 34388 8316 34621 8344
rect 34388 8304 34394 8316
rect 34609 8313 34621 8316
rect 34655 8313 34667 8347
rect 34609 8307 34667 8313
rect 37461 8347 37519 8353
rect 37461 8313 37473 8347
rect 37507 8344 37519 8347
rect 37826 8344 37832 8356
rect 37507 8316 37832 8344
rect 37507 8313 37519 8316
rect 37461 8307 37519 8313
rect 37826 8304 37832 8316
rect 37884 8304 37890 8356
rect 3694 8276 3700 8288
rect 3655 8248 3700 8276
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 7834 8276 7840 8288
rect 7795 8248 7840 8276
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 9401 8279 9459 8285
rect 9401 8276 9413 8279
rect 9272 8248 9413 8276
rect 9272 8236 9278 8248
rect 9401 8245 9413 8248
rect 9447 8245 9459 8279
rect 9401 8239 9459 8245
rect 17313 8279 17371 8285
rect 17313 8245 17325 8279
rect 17359 8276 17371 8279
rect 17586 8276 17592 8288
rect 17359 8248 17592 8276
rect 17359 8245 17371 8248
rect 17313 8239 17371 8245
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2498 8072 2504 8084
rect 1627 8044 2504 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6638 8072 6644 8084
rect 5776 8044 6644 8072
rect 5776 8032 5782 8044
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7892 8044 8217 8072
rect 7892 8032 7898 8044
rect 8205 8041 8217 8044
rect 8251 8072 8263 8075
rect 9214 8072 9220 8084
rect 8251 8044 9220 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 26326 8032 26332 8084
rect 26384 8072 26390 8084
rect 26697 8075 26755 8081
rect 26697 8072 26709 8075
rect 26384 8044 26709 8072
rect 26384 8032 26390 8044
rect 26697 8041 26709 8044
rect 26743 8041 26755 8075
rect 26697 8035 26755 8041
rect 8294 8004 8300 8016
rect 6886 7976 8300 8004
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 3752 7908 3801 7936
rect 3752 7896 3758 7908
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 3789 7899 3847 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6886 7936 6914 7976
rect 8294 7964 8300 7976
rect 8352 8004 8358 8016
rect 13998 8004 14004 8016
rect 8352 7976 14004 8004
rect 8352 7964 8358 7976
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 8018 7936 8024 7948
rect 5675 7908 6914 7936
rect 7979 7908 8024 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8904 7908 9045 7936
rect 8904 7896 8910 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 11054 7936 11060 7948
rect 11015 7908 11060 7936
rect 9033 7899 9091 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 24854 7936 24860 7948
rect 24767 7908 24860 7936
rect 24854 7896 24860 7908
rect 24912 7936 24918 7948
rect 25314 7936 25320 7948
rect 24912 7908 25320 7936
rect 24912 7896 24918 7908
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7868 1458 7880
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 1452 7840 2053 7868
rect 1452 7828 1458 7840
rect 2041 7837 2053 7840
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6696 7840 7205 7868
rect 6696 7828 6702 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7742 7868 7748 7880
rect 7432 7840 7748 7868
rect 7432 7828 7438 7840
rect 7742 7828 7748 7840
rect 7800 7868 7806 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7800 7840 7941 7868
rect 7800 7828 7806 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 8202 7868 8208 7880
rect 8115 7840 8208 7868
rect 7929 7831 7987 7837
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 3973 7803 4031 7809
rect 3973 7800 3985 7803
rect 3660 7772 3985 7800
rect 3660 7760 3666 7772
rect 3973 7769 3985 7772
rect 4019 7769 4031 7803
rect 7944 7800 7972 7831
rect 8202 7828 8208 7840
rect 8260 7868 8266 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 8260 7840 9229 7868
rect 8260 7828 8266 7840
rect 9217 7837 9229 7840
rect 9263 7868 9275 7871
rect 9674 7868 9680 7880
rect 9263 7840 9680 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 13998 7868 14004 7880
rect 11379 7840 14004 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 16574 7868 16580 7880
rect 16535 7840 16580 7868
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 20714 7868 20720 7880
rect 20675 7840 20720 7868
rect 20714 7828 20720 7840
rect 20772 7868 20778 7880
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 20772 7840 21465 7868
rect 20772 7828 20778 7840
rect 21453 7837 21465 7840
rect 21499 7868 21511 7871
rect 22094 7868 22100 7880
rect 21499 7840 22100 7868
rect 21499 7837 21511 7840
rect 21453 7831 21511 7837
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 25584 7871 25642 7877
rect 25584 7837 25596 7871
rect 25630 7868 25642 7871
rect 25958 7868 25964 7880
rect 25630 7840 25964 7868
rect 25630 7837 25642 7840
rect 25584 7831 25642 7837
rect 25958 7828 25964 7840
rect 26016 7828 26022 7880
rect 8941 7803 8999 7809
rect 8941 7800 8953 7803
rect 7944 7772 8953 7800
rect 3973 7763 4031 7769
rect 8941 7769 8953 7772
rect 8987 7769 8999 7803
rect 30006 7800 30012 7812
rect 8941 7763 8999 7769
rect 20916 7772 30012 7800
rect 20916 7744 20944 7772
rect 30006 7760 30012 7772
rect 30064 7760 30070 7812
rect 7377 7735 7435 7741
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 8202 7732 8208 7744
rect 7423 7704 8208 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 10594 7732 10600 7744
rect 9447 7704 10600 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 14090 7732 14096 7744
rect 14051 7704 14096 7732
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 16758 7732 16764 7744
rect 16719 7704 16764 7732
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 20898 7732 20904 7744
rect 20811 7704 20904 7732
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 3602 7528 3608 7540
rect 3563 7500 3608 7528
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 7742 7460 7748 7472
rect 7703 7432 7748 7460
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 9677 7463 9735 7469
rect 9677 7460 9689 7463
rect 8444 7432 9689 7460
rect 8444 7420 8450 7432
rect 9677 7429 9689 7432
rect 9723 7429 9735 7463
rect 13998 7460 14004 7472
rect 13959 7432 14004 7460
rect 9677 7423 9735 7429
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 17586 7460 17592 7472
rect 17547 7432 17592 7460
rect 17586 7420 17592 7432
rect 17644 7420 17650 7472
rect 18874 7420 18880 7472
rect 18932 7460 18938 7472
rect 26878 7460 26884 7472
rect 18932 7432 26884 7460
rect 18932 7420 18938 7432
rect 26878 7420 26884 7432
rect 26936 7420 26942 7472
rect 27522 7420 27528 7472
rect 27580 7460 27586 7472
rect 28905 7463 28963 7469
rect 28905 7460 28917 7463
rect 27580 7432 28917 7460
rect 27580 7420 27586 7432
rect 28905 7429 28917 7432
rect 28951 7429 28963 7463
rect 28905 7423 28963 7429
rect 30098 7420 30104 7472
rect 30156 7420 30162 7472
rect 30466 7420 30472 7472
rect 30524 7460 30530 7472
rect 30524 7432 30880 7460
rect 30524 7420 30530 7432
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7392 4123 7395
rect 5718 7392 5724 7404
rect 4111 7364 5724 7392
rect 4111 7361 4123 7364
rect 4065 7355 4123 7361
rect 3436 7324 3464 7355
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 7926 7392 7932 7404
rect 7887 7364 7932 7392
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8202 7392 8208 7404
rect 8067 7364 8208 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 18800 7364 23213 7392
rect 4706 7324 4712 7336
rect 3436 7296 4712 7324
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5350 7324 5356 7336
rect 5307 7296 5356 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 5583 7296 6377 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 6365 7293 6377 7296
rect 6411 7324 6423 7327
rect 7650 7324 7656 7336
rect 6411 7296 7656 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 12406 7296 13737 7324
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 12406 7256 12434 7296
rect 13725 7293 13737 7296
rect 13771 7324 13783 7327
rect 13814 7324 13820 7336
rect 13771 7296 13820 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7324 14243 7327
rect 14366 7324 14372 7336
rect 14231 7296 14372 7324
rect 14231 7293 14243 7296
rect 14185 7287 14243 7293
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 17954 7324 17960 7336
rect 17451 7296 17960 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 17954 7284 17960 7296
rect 18012 7324 18018 7336
rect 18800 7324 18828 7364
rect 23201 7361 23213 7364
rect 23247 7361 23259 7395
rect 30116 7392 30144 7420
rect 30561 7395 30619 7401
rect 30561 7392 30573 7395
rect 30116 7364 30573 7392
rect 23201 7355 23259 7361
rect 30561 7361 30573 7364
rect 30607 7361 30619 7395
rect 30742 7392 30748 7404
rect 30703 7364 30748 7392
rect 30561 7355 30619 7361
rect 18012 7296 18828 7324
rect 18012 7284 18018 7296
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 23293 7327 23351 7333
rect 18932 7296 19025 7324
rect 18932 7284 18938 7296
rect 23293 7293 23305 7327
rect 23339 7293 23351 7327
rect 23293 7287 23351 7293
rect 3476 7228 12434 7256
rect 3476 7216 3482 7228
rect 18138 7216 18144 7268
rect 18196 7256 18202 7268
rect 18892 7256 18920 7284
rect 18196 7228 18920 7256
rect 23308 7256 23336 7287
rect 23382 7284 23388 7336
rect 23440 7324 23446 7336
rect 27246 7324 27252 7336
rect 23440 7296 23485 7324
rect 27207 7296 27252 7324
rect 23440 7284 23446 7296
rect 27246 7284 27252 7296
rect 27304 7284 27310 7336
rect 29089 7327 29147 7333
rect 29089 7293 29101 7327
rect 29135 7324 29147 7327
rect 30098 7324 30104 7336
rect 29135 7296 30104 7324
rect 29135 7293 29147 7296
rect 29089 7287 29147 7293
rect 30098 7284 30104 7296
rect 30156 7284 30162 7336
rect 30576 7324 30604 7355
rect 30742 7352 30748 7364
rect 30800 7352 30806 7404
rect 30852 7401 30880 7432
rect 30837 7395 30895 7401
rect 30837 7361 30849 7395
rect 30883 7361 30895 7395
rect 30837 7355 30895 7361
rect 30926 7352 30932 7404
rect 30984 7392 30990 7404
rect 31202 7392 31208 7404
rect 30984 7364 31208 7392
rect 30984 7352 30990 7364
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 34054 7352 34060 7404
rect 34112 7392 34118 7404
rect 34149 7395 34207 7401
rect 34149 7392 34161 7395
rect 34112 7364 34161 7392
rect 34112 7352 34118 7364
rect 34149 7361 34161 7364
rect 34195 7361 34207 7395
rect 34330 7392 34336 7404
rect 34291 7364 34336 7392
rect 34149 7355 34207 7361
rect 34330 7352 34336 7364
rect 34388 7352 34394 7404
rect 32674 7324 32680 7336
rect 30576 7296 32680 7324
rect 32674 7284 32680 7296
rect 32732 7284 32738 7336
rect 24121 7259 24179 7265
rect 24121 7256 24133 7259
rect 23308 7228 24133 7256
rect 18196 7216 18202 7228
rect 24121 7225 24133 7228
rect 24167 7256 24179 7259
rect 37918 7256 37924 7268
rect 24167 7228 37924 7256
rect 24167 7225 24179 7228
rect 24121 7219 24179 7225
rect 37918 7216 37924 7228
rect 37976 7216 37982 7268
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7188 4307 7191
rect 4614 7188 4620 7200
rect 4295 7160 4620 7188
rect 4295 7157 4307 7160
rect 4249 7151 4307 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 7834 7188 7840 7200
rect 7795 7160 7840 7188
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 8205 7191 8263 7197
rect 8205 7157 8217 7191
rect 8251 7188 8263 7191
rect 8662 7188 8668 7200
rect 8251 7160 8668 7188
rect 8251 7157 8263 7160
rect 8205 7151 8263 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 19426 7188 19432 7200
rect 9815 7160 19432 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 22833 7191 22891 7197
rect 22833 7157 22845 7191
rect 22879 7188 22891 7191
rect 23106 7188 23112 7200
rect 22879 7160 23112 7188
rect 22879 7157 22891 7160
rect 22833 7151 22891 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 27246 7148 27252 7200
rect 27304 7188 27310 7200
rect 30009 7191 30067 7197
rect 30009 7188 30021 7191
rect 27304 7160 30021 7188
rect 27304 7148 27310 7160
rect 30009 7157 30021 7160
rect 30055 7188 30067 7191
rect 30926 7188 30932 7200
rect 30055 7160 30932 7188
rect 30055 7157 30067 7160
rect 30009 7151 30067 7157
rect 30926 7148 30932 7160
rect 30984 7148 30990 7200
rect 31205 7191 31263 7197
rect 31205 7157 31217 7191
rect 31251 7188 31263 7191
rect 33042 7188 33048 7200
rect 31251 7160 33048 7188
rect 31251 7157 31263 7160
rect 31205 7151 31263 7157
rect 33042 7148 33048 7160
rect 33100 7148 33106 7200
rect 34241 7191 34299 7197
rect 34241 7157 34253 7191
rect 34287 7188 34299 7191
rect 34514 7188 34520 7200
rect 34287 7160 34520 7188
rect 34287 7157 34299 7160
rect 34241 7151 34299 7157
rect 34514 7148 34520 7160
rect 34572 7148 34578 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 4249 6987 4307 6993
rect 4249 6953 4261 6987
rect 4295 6953 4307 6987
rect 4706 6984 4712 6996
rect 4667 6956 4712 6984
rect 4249 6947 4307 6953
rect 4264 6916 4292 6947
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4856 6956 5181 6984
rect 4856 6944 4862 6956
rect 5169 6953 5181 6956
rect 5215 6984 5227 6987
rect 5350 6984 5356 6996
rect 5215 6956 5356 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 7834 6984 7840 6996
rect 7795 6956 7840 6984
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 30285 6987 30343 6993
rect 30285 6953 30297 6987
rect 30331 6984 30343 6987
rect 30742 6984 30748 6996
rect 30331 6956 30748 6984
rect 30331 6953 30343 6956
rect 30285 6947 30343 6953
rect 30742 6944 30748 6956
rect 30800 6944 30806 6996
rect 33873 6987 33931 6993
rect 33873 6953 33885 6987
rect 33919 6984 33931 6987
rect 34330 6984 34336 6996
rect 33919 6956 34336 6984
rect 33919 6953 33931 6956
rect 33873 6947 33931 6953
rect 34330 6944 34336 6956
rect 34388 6944 34394 6996
rect 4816 6916 4844 6944
rect 4264 6888 4844 6916
rect 34514 6876 34520 6928
rect 34572 6916 34578 6928
rect 35158 6916 35164 6928
rect 34572 6888 35164 6916
rect 34572 6876 34578 6888
rect 35158 6876 35164 6888
rect 35216 6876 35222 6928
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 4120 6820 4169 6848
rect 4120 6808 4126 6820
rect 4157 6817 4169 6820
rect 4203 6848 4215 6851
rect 4982 6848 4988 6860
rect 4203 6820 4988 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 10594 6848 10600 6860
rect 10555 6820 10600 6848
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 15102 6848 15108 6860
rect 13872 6820 15108 6848
rect 13872 6808 13878 6820
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6780 1458 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1452 6752 2053 6780
rect 1452 6740 1458 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 2041 6743 2099 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4522 6780 4528 6792
rect 4172 6752 4528 6780
rect 3988 6712 4016 6740
rect 4172 6712 4200 6752
rect 4522 6740 4528 6752
rect 4580 6780 4586 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4580 6752 4905 6780
rect 4580 6740 4586 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8202 6780 8208 6792
rect 8067 6752 8208 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8720 6752 8953 6780
rect 8720 6740 8726 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 12894 6780 12900 6792
rect 10919 6752 12900 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 14108 6789 14136 6820
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 16758 6848 16764 6860
rect 16719 6820 16764 6848
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6848 18475 6851
rect 19426 6848 19432 6860
rect 18463 6820 18552 6848
rect 19387 6820 19432 6848
rect 18463 6817 18475 6820
rect 18417 6811 18475 6817
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6749 14151 6783
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14093 6743 14151 6749
rect 14200 6752 14473 6780
rect 3988 6684 4200 6712
rect 4249 6715 4307 6721
rect 4249 6681 4261 6715
rect 4295 6712 4307 6715
rect 4614 6712 4620 6724
rect 4295 6684 4620 6712
rect 4295 6681 4307 6684
rect 4249 6675 4307 6681
rect 4614 6672 4620 6684
rect 4672 6712 4678 6724
rect 5166 6712 5172 6724
rect 4672 6684 5172 6712
rect 4672 6672 4678 6684
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 7742 6712 7748 6724
rect 7703 6684 7748 6712
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 14200 6712 14228 6752
rect 14461 6749 14473 6752
rect 14507 6780 14519 6783
rect 15930 6780 15936 6792
rect 14507 6752 15936 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 13320 6684 14228 6712
rect 14277 6715 14335 6721
rect 13320 6672 13326 6684
rect 14277 6681 14289 6715
rect 14323 6681 14335 6715
rect 14277 6675 14335 6681
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 8202 6644 8208 6656
rect 8163 6616 8208 6644
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 14292 6644 14320 6675
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 16592 6712 16620 6743
rect 16758 6712 16764 6724
rect 14424 6684 14469 6712
rect 14568 6684 16528 6712
rect 16592 6684 16764 6712
rect 14424 6672 14430 6684
rect 14568 6644 14596 6684
rect 14292 6616 14596 6644
rect 14645 6647 14703 6653
rect 14645 6613 14657 6647
rect 14691 6644 14703 6647
rect 14734 6644 14740 6656
rect 14691 6616 14740 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15102 6644 15108 6656
rect 15063 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 16500 6644 16528 6684
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 18524 6656 18552 6820
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 20714 6848 20720 6860
rect 20675 6820 20720 6848
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6848 23167 6851
rect 23382 6848 23388 6860
rect 23155 6820 23388 6848
rect 23155 6817 23167 6820
rect 23109 6811 23167 6817
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 24486 6848 24492 6860
rect 24447 6820 24492 6848
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 30466 6848 30472 6860
rect 30208 6820 30472 6848
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19260 6712 19288 6743
rect 22094 6740 22100 6792
rect 22152 6780 22158 6792
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 22152 6752 23213 6780
rect 22152 6740 22158 6752
rect 23201 6749 23213 6752
rect 23247 6780 23259 6783
rect 23934 6780 23940 6792
rect 23247 6752 23940 6780
rect 23247 6749 23259 6752
rect 23201 6743 23259 6749
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 20162 6712 20168 6724
rect 19260 6684 20168 6712
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 23293 6715 23351 6721
rect 23293 6681 23305 6715
rect 23339 6712 23351 6715
rect 23566 6712 23572 6724
rect 23339 6684 23572 6712
rect 23339 6681 23351 6684
rect 23293 6675 23351 6681
rect 23566 6672 23572 6684
rect 23624 6712 23630 6724
rect 24504 6712 24532 6808
rect 30208 6789 30236 6820
rect 30466 6808 30472 6820
rect 30524 6808 30530 6860
rect 34054 6808 34060 6860
rect 34112 6848 34118 6860
rect 34112 6820 34284 6848
rect 34112 6808 34118 6820
rect 30193 6783 30251 6789
rect 30193 6749 30205 6783
rect 30239 6749 30251 6783
rect 30374 6780 30380 6792
rect 30335 6752 30380 6780
rect 30193 6743 30251 6749
rect 30374 6740 30380 6752
rect 30432 6740 30438 6792
rect 33042 6740 33048 6792
rect 33100 6780 33106 6792
rect 34146 6780 34152 6792
rect 33100 6752 34008 6780
rect 34107 6752 34152 6780
rect 33100 6740 33106 6752
rect 33870 6712 33876 6724
rect 23624 6684 24532 6712
rect 33831 6684 33876 6712
rect 23624 6672 23630 6684
rect 33870 6672 33876 6684
rect 33928 6672 33934 6724
rect 33980 6712 34008 6752
rect 34146 6740 34152 6752
rect 34204 6740 34210 6792
rect 34256 6780 34284 6820
rect 34606 6808 34612 6860
rect 34664 6848 34670 6860
rect 35802 6848 35808 6860
rect 34664 6820 35808 6848
rect 34664 6808 34670 6820
rect 35802 6808 35808 6820
rect 35860 6848 35866 6860
rect 36357 6851 36415 6857
rect 36357 6848 36369 6851
rect 35860 6820 36369 6848
rect 35860 6808 35866 6820
rect 36357 6817 36369 6820
rect 36403 6817 36415 6851
rect 36357 6811 36415 6817
rect 34977 6783 35035 6789
rect 34977 6780 34989 6783
rect 34256 6752 34989 6780
rect 34977 6749 34989 6752
rect 35023 6749 35035 6783
rect 34977 6743 35035 6749
rect 35069 6783 35127 6789
rect 35069 6749 35081 6783
rect 35115 6749 35127 6783
rect 35069 6743 35127 6749
rect 33980 6684 34836 6712
rect 17034 6644 17040 6656
rect 16500 6616 17040 6644
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 23198 6644 23204 6656
rect 18564 6616 23204 6644
rect 18564 6604 18570 6616
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 23474 6604 23480 6656
rect 23532 6644 23538 6656
rect 23661 6647 23719 6653
rect 23661 6644 23673 6647
rect 23532 6616 23673 6644
rect 23532 6604 23538 6616
rect 23661 6613 23673 6616
rect 23707 6613 23719 6647
rect 34054 6644 34060 6656
rect 34015 6616 34060 6644
rect 23661 6607 23719 6613
rect 34054 6604 34060 6616
rect 34112 6604 34118 6656
rect 34698 6644 34704 6656
rect 34659 6616 34704 6644
rect 34698 6604 34704 6616
rect 34756 6604 34762 6656
rect 34808 6644 34836 6684
rect 34882 6672 34888 6724
rect 34940 6712 34946 6724
rect 35084 6712 35112 6743
rect 35158 6740 35164 6792
rect 35216 6780 35222 6792
rect 35216 6752 35261 6780
rect 35216 6740 35222 6752
rect 35342 6740 35348 6792
rect 35400 6780 35406 6792
rect 35400 6752 35445 6780
rect 35400 6740 35406 6752
rect 36602 6715 36660 6721
rect 36602 6712 36614 6715
rect 34940 6684 35112 6712
rect 35866 6684 36614 6712
rect 34940 6672 34946 6684
rect 35866 6644 35894 6684
rect 36602 6681 36614 6684
rect 36648 6681 36660 6715
rect 36602 6675 36660 6681
rect 37734 6644 37740 6656
rect 34808 6616 35894 6644
rect 37695 6616 37740 6644
rect 37734 6604 37740 6616
rect 37792 6604 37798 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 14274 6400 14280 6452
rect 14332 6440 14338 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 14332 6412 14565 6440
rect 14332 6400 14338 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16761 6443 16819 6449
rect 16761 6440 16773 6443
rect 16448 6412 16773 6440
rect 16448 6400 16454 6412
rect 16761 6409 16773 6412
rect 16807 6440 16819 6443
rect 18506 6440 18512 6452
rect 16807 6412 18512 6440
rect 16807 6409 16819 6412
rect 16761 6403 16819 6409
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 20625 6443 20683 6449
rect 20625 6409 20637 6443
rect 20671 6440 20683 6443
rect 20898 6440 20904 6452
rect 20671 6412 20904 6440
rect 20671 6409 20683 6412
rect 20625 6403 20683 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 22278 6400 22284 6452
rect 22336 6440 22342 6452
rect 22465 6443 22523 6449
rect 22465 6440 22477 6443
rect 22336 6412 22477 6440
rect 22336 6400 22342 6412
rect 22465 6409 22477 6412
rect 22511 6409 22523 6443
rect 23934 6440 23940 6452
rect 23895 6412 23940 6440
rect 22465 6403 22523 6409
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 33045 6443 33103 6449
rect 33045 6409 33057 6443
rect 33091 6440 33103 6443
rect 34882 6440 34888 6452
rect 33091 6412 34888 6440
rect 33091 6409 33103 6412
rect 33045 6403 33103 6409
rect 34882 6400 34888 6412
rect 34940 6400 34946 6452
rect 5629 6375 5687 6381
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 7742 6372 7748 6384
rect 5675 6344 7748 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 12980 6375 13038 6381
rect 12980 6341 12992 6375
rect 13026 6372 13038 6375
rect 14090 6372 14096 6384
rect 13026 6344 14096 6372
rect 13026 6341 13038 6344
rect 12980 6335 13038 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 20162 6332 20168 6384
rect 20220 6372 20226 6384
rect 22373 6375 22431 6381
rect 22373 6372 22385 6375
rect 20220 6344 22385 6372
rect 20220 6332 20226 6344
rect 22373 6341 22385 6344
rect 22419 6341 22431 6375
rect 22373 6335 22431 6341
rect 23198 6332 23204 6384
rect 23256 6372 23262 6384
rect 27338 6372 27344 6384
rect 23256 6344 27344 6372
rect 23256 6332 23262 6344
rect 27338 6332 27344 6344
rect 27396 6332 27402 6384
rect 27525 6375 27583 6381
rect 27525 6341 27537 6375
rect 27571 6372 27583 6375
rect 28074 6372 28080 6384
rect 27571 6344 28080 6372
rect 27571 6341 27583 6344
rect 27525 6335 27583 6341
rect 28074 6332 28080 6344
rect 28132 6332 28138 6384
rect 34698 6332 34704 6384
rect 34756 6372 34762 6384
rect 35630 6375 35688 6381
rect 35630 6372 35642 6375
rect 34756 6344 35642 6372
rect 34756 6332 34762 6344
rect 35630 6341 35642 6344
rect 35676 6341 35688 6375
rect 35630 6335 35688 6341
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4706 6304 4712 6316
rect 4580 6276 4712 6304
rect 4580 6264 4586 6276
rect 4706 6264 4712 6276
rect 4764 6304 4770 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 4764 6276 5365 6304
rect 4764 6264 4770 6276
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 8260 6276 8401 6304
rect 8260 6264 8266 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 14734 6304 14740 6316
rect 14695 6276 14740 6304
rect 8389 6267 8447 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 19058 6304 19064 6316
rect 19019 6276 19064 6304
rect 19058 6264 19064 6276
rect 19116 6264 19122 6316
rect 32953 6307 33011 6313
rect 32953 6273 32965 6307
rect 32999 6273 33011 6307
rect 33134 6304 33140 6316
rect 33095 6276 33140 6304
rect 32953 6267 33011 6273
rect 2682 6236 2688 6248
rect 2643 6208 2688 6236
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 2866 6236 2872 6248
rect 2827 6208 2872 6236
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3234 6236 3240 6248
rect 3195 6208 3240 6236
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 4948 6208 5457 6236
rect 4948 6196 4954 6208
rect 5445 6205 5457 6208
rect 5491 6236 5503 6239
rect 7834 6236 7840 6248
rect 5491 6208 7840 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6205 14979 6239
rect 14921 6199 14979 6205
rect 22281 6239 22339 6245
rect 22281 6205 22293 6239
rect 22327 6236 22339 6239
rect 23382 6236 23388 6248
rect 22327 6208 23388 6236
rect 22327 6205 22339 6208
rect 22281 6199 22339 6205
rect 4798 6128 4804 6180
rect 4856 6168 4862 6180
rect 4856 6140 5396 6168
rect 4856 6128 4862 6140
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5368 6109 5396 6140
rect 5353 6103 5411 6109
rect 5353 6069 5365 6103
rect 5399 6069 5411 6103
rect 5353 6063 5411 6069
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6100 8631 6103
rect 10318 6100 10324 6112
rect 8619 6072 10324 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 12728 6100 12756 6199
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6168 14151 6171
rect 14366 6168 14372 6180
rect 14139 6140 14372 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 13998 6100 14004 6112
rect 12728 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14936 6100 14964 6199
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 32968 6236 32996 6267
rect 33134 6264 33140 6276
rect 33192 6264 33198 6316
rect 34057 6307 34115 6313
rect 34057 6273 34069 6307
rect 34103 6304 34115 6307
rect 34146 6304 34152 6316
rect 34103 6276 34152 6304
rect 34103 6273 34115 6276
rect 34057 6267 34115 6273
rect 34146 6264 34152 6276
rect 34204 6264 34210 6316
rect 35802 6264 35808 6316
rect 35860 6304 35866 6316
rect 35897 6307 35955 6313
rect 35897 6304 35909 6307
rect 35860 6276 35909 6304
rect 35860 6264 35866 6276
rect 35897 6273 35909 6276
rect 35943 6273 35955 6307
rect 37826 6304 37832 6316
rect 37787 6276 37832 6304
rect 35897 6267 35955 6273
rect 37826 6264 37832 6276
rect 37884 6264 37890 6316
rect 33042 6236 33048 6248
rect 32968 6208 33048 6236
rect 33042 6196 33048 6208
rect 33100 6236 33106 6248
rect 33870 6236 33876 6248
rect 33100 6208 33876 6236
rect 33100 6196 33106 6208
rect 33870 6196 33876 6208
rect 33928 6196 33934 6248
rect 33962 6196 33968 6248
rect 34020 6236 34026 6248
rect 34020 6208 34065 6236
rect 34020 6196 34026 6208
rect 15102 6128 15108 6180
rect 15160 6168 15166 6180
rect 25682 6168 25688 6180
rect 15160 6140 25688 6168
rect 15160 6128 15166 6140
rect 25682 6128 25688 6140
rect 25740 6128 25746 6180
rect 25774 6128 25780 6180
rect 25832 6168 25838 6180
rect 27341 6171 27399 6177
rect 27341 6168 27353 6171
rect 25832 6140 27353 6168
rect 25832 6128 25838 6140
rect 27341 6137 27353 6140
rect 27387 6137 27399 6171
rect 33686 6168 33692 6180
rect 33647 6140 33692 6168
rect 27341 6131 27399 6137
rect 33686 6128 33692 6140
rect 33744 6128 33750 6180
rect 15473 6103 15531 6109
rect 15473 6100 15485 6103
rect 14936 6072 15485 6100
rect 15473 6069 15485 6072
rect 15519 6100 15531 6103
rect 16206 6100 16212 6112
rect 15519 6072 16212 6100
rect 15519 6069 15531 6072
rect 15473 6063 15531 6069
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 19150 6100 19156 6112
rect 19111 6072 19156 6100
rect 19150 6060 19156 6072
rect 19208 6060 19214 6112
rect 22833 6103 22891 6109
rect 22833 6069 22845 6103
rect 22879 6100 22891 6103
rect 23198 6100 23204 6112
rect 22879 6072 23204 6100
rect 22879 6069 22891 6072
rect 22833 6063 22891 6069
rect 23198 6060 23204 6072
rect 23256 6060 23262 6112
rect 33870 6100 33876 6112
rect 33831 6072 33876 6100
rect 33870 6060 33876 6072
rect 33928 6100 33934 6112
rect 34054 6100 34060 6112
rect 33928 6072 34060 6100
rect 33928 6060 33934 6072
rect 34054 6060 34060 6072
rect 34112 6100 34118 6112
rect 34517 6103 34575 6109
rect 34517 6100 34529 6103
rect 34112 6072 34529 6100
rect 34112 6060 34118 6072
rect 34517 6069 34529 6072
rect 34563 6069 34575 6103
rect 38010 6100 38016 6112
rect 37971 6072 38016 6100
rect 34517 6063 34575 6069
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2682 5896 2688 5908
rect 2643 5868 2688 5896
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 2924 5868 3801 5896
rect 2924 5856 2930 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 4798 5896 4804 5908
rect 4759 5868 4804 5896
rect 3789 5859 3847 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 14056 5868 14197 5896
rect 14056 5856 14062 5868
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 16850 5896 16856 5908
rect 15988 5868 16856 5896
rect 15988 5856 15994 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 21174 5856 21180 5908
rect 21232 5896 21238 5908
rect 21232 5868 31754 5896
rect 21232 5856 21238 5868
rect 3418 5788 3424 5840
rect 3476 5828 3482 5840
rect 16390 5828 16396 5840
rect 3476 5800 16396 5828
rect 3476 5788 3482 5800
rect 16390 5788 16396 5800
rect 16448 5788 16454 5840
rect 17681 5831 17739 5837
rect 17681 5828 17693 5831
rect 16776 5800 17693 5828
rect 4890 5760 4896 5772
rect 4851 5732 4896 5760
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 9122 5760 9128 5772
rect 9083 5732 9128 5760
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 13078 5760 13084 5772
rect 12032 5732 13084 5760
rect 12032 5720 12038 5732
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13412 5732 13553 5760
rect 13412 5720 13418 5732
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 16206 5720 16212 5772
rect 16264 5760 16270 5772
rect 16776 5769 16804 5800
rect 17681 5797 17693 5800
rect 17727 5828 17739 5831
rect 29730 5828 29736 5840
rect 17727 5800 29736 5828
rect 17727 5797 17739 5800
rect 17681 5791 17739 5797
rect 29730 5788 29736 5800
rect 29788 5788 29794 5840
rect 30193 5831 30251 5837
rect 30193 5797 30205 5831
rect 30239 5828 30251 5831
rect 30374 5828 30380 5840
rect 30239 5800 30380 5828
rect 30239 5797 30251 5800
rect 30193 5791 30251 5797
rect 30374 5788 30380 5800
rect 30432 5788 30438 5840
rect 31726 5828 31754 5868
rect 32858 5856 32864 5908
rect 32916 5896 32922 5908
rect 34606 5896 34612 5908
rect 32916 5868 34612 5896
rect 32916 5856 32922 5868
rect 34606 5856 34612 5868
rect 34664 5896 34670 5908
rect 34701 5899 34759 5905
rect 34701 5896 34713 5899
rect 34664 5868 34713 5896
rect 34664 5856 34670 5868
rect 34701 5865 34713 5868
rect 34747 5865 34759 5899
rect 34701 5859 34759 5865
rect 33134 5828 33140 5840
rect 31726 5800 33140 5828
rect 33134 5788 33140 5800
rect 33192 5788 33198 5840
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 16264 5732 16773 5760
rect 16264 5720 16270 5732
rect 16761 5729 16773 5732
rect 16807 5729 16819 5763
rect 22554 5760 22560 5772
rect 16761 5723 16819 5729
rect 20088 5732 22560 5760
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3844 5664 3985 5692
rect 3844 5652 3850 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4614 5652 4620 5704
rect 4672 5652 4678 5704
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 4764 5664 4809 5692
rect 4764 5652 4770 5664
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8352 5664 8953 5692
rect 8352 5652 8358 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 15930 5692 15936 5704
rect 15891 5664 15936 5692
rect 8941 5655 8999 5661
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4632 5624 4660 5652
rect 4985 5627 5043 5633
rect 4985 5624 4997 5627
rect 4212 5596 4997 5624
rect 4212 5584 4218 5596
rect 4985 5593 4997 5596
rect 5031 5593 5043 5627
rect 8956 5624 8984 5655
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16390 5692 16396 5704
rect 16347 5664 16396 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16942 5692 16948 5704
rect 16903 5664 16948 5692
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 20088 5701 20116 5732
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 22738 5720 22744 5772
rect 22796 5760 22802 5772
rect 22925 5763 22983 5769
rect 22925 5760 22937 5763
rect 22796 5732 22937 5760
rect 22796 5720 22802 5732
rect 22925 5729 22937 5732
rect 22971 5729 22983 5763
rect 23106 5760 23112 5772
rect 23067 5732 23112 5760
rect 22925 5723 22983 5729
rect 23106 5720 23112 5732
rect 23164 5720 23170 5772
rect 33045 5763 33103 5769
rect 33045 5729 33057 5763
rect 33091 5760 33103 5763
rect 33870 5760 33876 5772
rect 33091 5732 33876 5760
rect 33091 5729 33103 5732
rect 33045 5723 33103 5729
rect 33870 5720 33876 5732
rect 33928 5720 33934 5772
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 19484 5664 20085 5692
rect 19484 5652 19490 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 20162 5652 20168 5704
rect 20220 5692 20226 5704
rect 20441 5695 20499 5701
rect 20220 5664 20265 5692
rect 20220 5652 20226 5664
rect 20441 5661 20453 5695
rect 20487 5692 20499 5695
rect 20898 5692 20904 5704
rect 20487 5664 20904 5692
rect 20487 5661 20499 5664
rect 20441 5655 20499 5661
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 23198 5692 23204 5704
rect 23159 5664 23204 5692
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 23566 5692 23572 5704
rect 23400 5664 23572 5692
rect 10594 5624 10600 5636
rect 8956 5596 10600 5624
rect 4985 5587 5043 5593
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 10778 5624 10784 5636
rect 10739 5596 10784 5624
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 13357 5627 13415 5633
rect 13357 5624 13369 5627
rect 12952 5596 13369 5624
rect 12952 5584 12958 5596
rect 13357 5593 13369 5596
rect 13403 5593 13415 5627
rect 13357 5587 13415 5593
rect 16025 5627 16083 5633
rect 16025 5593 16037 5627
rect 16071 5593 16083 5627
rect 16025 5587 16083 5593
rect 16117 5627 16175 5633
rect 16117 5593 16129 5627
rect 16163 5624 16175 5627
rect 17034 5624 17040 5636
rect 16163 5596 17040 5624
rect 16163 5593 16175 5596
rect 16117 5587 16175 5593
rect 4525 5559 4583 5565
rect 4525 5525 4537 5559
rect 4571 5556 4583 5559
rect 4614 5556 4620 5568
rect 4571 5528 4620 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13630 5556 13636 5568
rect 13136 5528 13636 5556
rect 13136 5516 13142 5528
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 15930 5556 15936 5568
rect 15795 5528 15936 5556
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 16040 5556 16068 5587
rect 17034 5584 17040 5596
rect 17092 5584 17098 5636
rect 19058 5584 19064 5636
rect 19116 5624 19122 5636
rect 20257 5627 20315 5633
rect 20257 5624 20269 5627
rect 19116 5596 20269 5624
rect 19116 5584 19122 5596
rect 20257 5593 20269 5596
rect 20303 5624 20315 5627
rect 23290 5624 23296 5636
rect 20303 5596 23296 5624
rect 20303 5593 20315 5596
rect 20257 5587 20315 5593
rect 23290 5584 23296 5596
rect 23348 5584 23354 5636
rect 16758 5556 16764 5568
rect 16040 5528 16764 5556
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 17129 5559 17187 5565
rect 17129 5525 17141 5559
rect 17175 5556 17187 5559
rect 17402 5556 17408 5568
rect 17175 5528 17408 5556
rect 17175 5525 17187 5528
rect 17129 5519 17187 5525
rect 17402 5516 17408 5528
rect 17460 5516 17466 5568
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 19978 5556 19984 5568
rect 19935 5528 19984 5556
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 20772 5528 21097 5556
rect 20772 5516 20778 5528
rect 21085 5525 21097 5528
rect 21131 5556 21143 5559
rect 23400 5556 23428 5664
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 30098 5692 30104 5704
rect 30059 5664 30104 5692
rect 30098 5652 30104 5664
rect 30156 5692 30162 5704
rect 32953 5695 33011 5701
rect 30156 5664 31754 5692
rect 30156 5652 30162 5664
rect 31726 5624 31754 5664
rect 32953 5661 32965 5695
rect 32999 5692 33011 5695
rect 33134 5692 33140 5704
rect 32999 5664 33140 5692
rect 32999 5661 33011 5664
rect 32953 5655 33011 5661
rect 33134 5652 33140 5664
rect 33192 5652 33198 5704
rect 33226 5652 33232 5704
rect 33284 5692 33290 5704
rect 33284 5664 33329 5692
rect 33284 5652 33290 5664
rect 37734 5624 37740 5636
rect 31726 5596 37740 5624
rect 37734 5584 37740 5596
rect 37792 5584 37798 5636
rect 21131 5528 23428 5556
rect 23569 5559 23627 5565
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 23569 5525 23581 5559
rect 23615 5556 23627 5559
rect 25130 5556 25136 5568
rect 23615 5528 25136 5556
rect 23615 5525 23627 5528
rect 23569 5519 23627 5525
rect 25130 5516 25136 5528
rect 25188 5516 25194 5568
rect 32214 5516 32220 5568
rect 32272 5556 32278 5568
rect 32769 5559 32827 5565
rect 32769 5556 32781 5559
rect 32272 5528 32781 5556
rect 32272 5516 32278 5528
rect 32769 5525 32781 5528
rect 32815 5525 32827 5559
rect 32769 5519 32827 5525
rect 33318 5516 33324 5568
rect 33376 5556 33382 5568
rect 33781 5559 33839 5565
rect 33781 5556 33793 5559
rect 33376 5528 33793 5556
rect 33376 5516 33382 5528
rect 33781 5525 33793 5528
rect 33827 5525 33839 5559
rect 33781 5519 33839 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 2222 5352 2228 5364
rect 1627 5324 2228 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 15289 5355 15347 5361
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 16206 5352 16212 5364
rect 15335 5324 16212 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5216 1458 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1452 5188 2053 5216
rect 1452 5176 1458 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3712 5216 3740 5315
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 16942 5352 16948 5364
rect 16715 5324 16948 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17954 5352 17960 5364
rect 17184 5324 17960 5352
rect 17184 5312 17190 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 22097 5355 22155 5361
rect 22097 5321 22109 5355
rect 22143 5321 22155 5355
rect 22097 5315 22155 5321
rect 4154 5284 4160 5296
rect 4115 5256 4160 5284
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 10318 5284 10324 5296
rect 10279 5256 10324 5284
rect 10318 5244 10324 5256
rect 10376 5244 10382 5296
rect 12342 5284 12348 5296
rect 11716 5256 12348 5284
rect 3283 5188 3740 5216
rect 3881 5219 3939 5225
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 3970 5216 3976 5228
rect 3927 5188 3976 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 11716 5225 11744 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 13449 5287 13507 5293
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 17034 5284 17040 5296
rect 13495 5256 17040 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 17034 5244 17040 5256
rect 17092 5284 17098 5296
rect 19150 5284 19156 5296
rect 17092 5256 19156 5284
rect 17092 5244 17098 5256
rect 19150 5244 19156 5256
rect 19208 5284 19214 5296
rect 20806 5284 20812 5296
rect 19208 5256 20668 5284
rect 20767 5256 20812 5284
rect 19208 5244 19214 5256
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5224 5188 5457 5216
rect 5224 5176 5230 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 4062 5148 4068 5160
rect 4023 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 8754 5108 8760 5160
rect 8812 5148 8818 5160
rect 10045 5151 10103 5157
rect 10045 5148 10057 5151
rect 8812 5120 10057 5148
rect 8812 5108 8818 5120
rect 10045 5117 10057 5120
rect 10091 5117 10103 5151
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 10045 5111 10103 5117
rect 4798 5080 4804 5092
rect 4172 5052 4804 5080
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 4172 5021 4200 5052
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 10060 5080 10088 5111
rect 10502 5108 10508 5120
rect 10560 5148 10566 5160
rect 11808 5148 11836 5179
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 12069 5219 12127 5225
rect 11940 5188 11985 5216
rect 11940 5176 11946 5188
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 13262 5216 13268 5228
rect 12115 5188 12296 5216
rect 13223 5188 13268 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 10560 5120 11836 5148
rect 10560 5108 10566 5120
rect 12268 5080 12296 5188
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 13630 5216 13636 5228
rect 13412 5188 13457 5216
rect 13543 5188 13636 5216
rect 13412 5176 13418 5188
rect 13630 5176 13636 5188
rect 13688 5216 13694 5228
rect 14182 5216 14188 5228
rect 13688 5188 14188 5216
rect 13688 5176 13694 5188
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16850 5216 16856 5228
rect 16811 5188 16856 5216
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17126 5216 17132 5228
rect 16991 5188 17132 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 17681 5219 17739 5225
rect 17681 5216 17693 5219
rect 17276 5188 17693 5216
rect 17276 5176 17282 5188
rect 17681 5185 17693 5188
rect 17727 5216 17739 5219
rect 18138 5216 18144 5228
rect 17727 5188 18144 5216
rect 17727 5185 17739 5188
rect 17681 5179 17739 5185
rect 18138 5176 18144 5188
rect 18196 5176 18202 5228
rect 18966 5216 18972 5228
rect 18879 5188 18972 5216
rect 18966 5176 18972 5188
rect 19024 5216 19030 5228
rect 19613 5219 19671 5225
rect 19024 5188 19564 5216
rect 19024 5176 19030 5188
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 16206 5148 16212 5160
rect 16163 5120 16212 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 19426 5148 19432 5160
rect 17092 5120 19432 5148
rect 17092 5108 17098 5120
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19536 5148 19564 5188
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 19978 5216 19984 5228
rect 19659 5188 19984 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 20530 5216 20536 5228
rect 20491 5188 20536 5216
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 20640 5216 20668 5256
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 20640 5188 20729 5216
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 19797 5151 19855 5157
rect 19797 5148 19809 5151
rect 19536 5120 19809 5148
rect 19797 5117 19809 5120
rect 19843 5148 19855 5151
rect 20254 5148 20260 5160
rect 19843 5120 20260 5148
rect 19843 5117 19855 5120
rect 19797 5111 19855 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 20824 5148 20852 5244
rect 20937 5219 20995 5225
rect 20937 5185 20949 5219
rect 20983 5216 20995 5219
rect 22112 5216 22140 5315
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22336 5324 22477 5352
rect 22336 5312 22342 5324
rect 22465 5321 22477 5324
rect 22511 5321 22523 5355
rect 22465 5315 22523 5321
rect 22557 5355 22615 5361
rect 22557 5321 22569 5355
rect 22603 5352 22615 5355
rect 23106 5352 23112 5364
rect 22603 5324 23112 5352
rect 22603 5321 22615 5324
rect 22557 5315 22615 5321
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 24673 5355 24731 5361
rect 23308 5324 23612 5352
rect 23308 5284 23336 5324
rect 23474 5284 23480 5296
rect 20983 5188 22140 5216
rect 22664 5256 23336 5284
rect 23435 5256 23480 5284
rect 20983 5185 20995 5188
rect 20937 5179 20995 5185
rect 22664 5148 22692 5256
rect 23474 5244 23480 5256
rect 23532 5244 23538 5296
rect 23584 5228 23612 5324
rect 24673 5321 24685 5355
rect 24719 5321 24731 5355
rect 25130 5352 25136 5364
rect 25091 5324 25136 5352
rect 24673 5315 24731 5321
rect 23290 5216 23296 5228
rect 23251 5188 23296 5216
rect 23290 5176 23296 5188
rect 23348 5176 23354 5228
rect 23566 5216 23572 5228
rect 23479 5188 23572 5216
rect 23566 5176 23572 5188
rect 23624 5176 23630 5228
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5216 23719 5219
rect 24688 5216 24716 5315
rect 25130 5312 25136 5324
rect 25188 5312 25194 5364
rect 27433 5355 27491 5361
rect 27433 5321 27445 5355
rect 27479 5352 27491 5355
rect 27614 5352 27620 5364
rect 27479 5324 27620 5352
rect 27479 5321 27491 5324
rect 27433 5315 27491 5321
rect 27614 5312 27620 5324
rect 27672 5352 27678 5364
rect 29181 5355 29239 5361
rect 29181 5352 29193 5355
rect 27672 5324 29193 5352
rect 27672 5312 27678 5324
rect 29181 5321 29193 5324
rect 29227 5321 29239 5355
rect 29181 5315 29239 5321
rect 30285 5355 30343 5361
rect 30285 5321 30297 5355
rect 30331 5352 30343 5355
rect 30834 5352 30840 5364
rect 30331 5324 30840 5352
rect 30331 5321 30343 5324
rect 30285 5315 30343 5321
rect 27338 5284 27344 5296
rect 27251 5256 27344 5284
rect 27338 5244 27344 5256
rect 27396 5284 27402 5296
rect 30300 5284 30328 5315
rect 30834 5312 30840 5324
rect 30892 5312 30898 5364
rect 32861 5355 32919 5361
rect 32861 5321 32873 5355
rect 32907 5352 32919 5355
rect 33226 5352 33232 5364
rect 32907 5324 33232 5352
rect 32907 5321 32919 5324
rect 32861 5315 32919 5321
rect 33226 5312 33232 5324
rect 33284 5312 33290 5364
rect 33962 5352 33968 5364
rect 33612 5324 33968 5352
rect 33612 5293 33640 5324
rect 33962 5312 33968 5324
rect 34020 5352 34026 5364
rect 34241 5355 34299 5361
rect 34241 5352 34253 5355
rect 34020 5324 34253 5352
rect 34020 5312 34026 5324
rect 34241 5321 34253 5324
rect 34287 5321 34299 5355
rect 34241 5315 34299 5321
rect 33597 5287 33655 5293
rect 33597 5284 33609 5287
rect 27396 5256 30328 5284
rect 31864 5256 33609 5284
rect 27396 5244 27402 5256
rect 23707 5188 24716 5216
rect 25041 5219 25099 5225
rect 23707 5185 23719 5188
rect 23661 5179 23719 5185
rect 25041 5185 25053 5219
rect 25087 5216 25099 5219
rect 25958 5216 25964 5228
rect 25087 5188 25964 5216
rect 25087 5185 25099 5188
rect 25041 5179 25099 5185
rect 25958 5176 25964 5188
rect 26016 5176 26022 5228
rect 29178 5219 29236 5225
rect 29178 5185 29190 5219
rect 29224 5216 29236 5219
rect 30282 5219 30340 5225
rect 30282 5216 30294 5219
rect 29224 5188 30294 5216
rect 29224 5185 29236 5188
rect 29178 5179 29236 5185
rect 30282 5185 30294 5188
rect 30328 5216 30340 5219
rect 30328 5188 31754 5216
rect 30328 5185 30340 5188
rect 30282 5179 30340 5185
rect 20824 5120 22692 5148
rect 22738 5108 22744 5160
rect 22796 5148 22802 5160
rect 25317 5151 25375 5157
rect 22796 5120 24808 5148
rect 22796 5108 22802 5120
rect 10060 5052 12296 5080
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2924 4984 3065 5012
rect 2924 4972 2930 4984
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 3053 4975 3111 4981
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 4981 4215 5015
rect 4157 4975 4215 4981
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 4706 5012 4712 5024
rect 4663 4984 4712 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5074 4972 5080 5024
rect 5132 5012 5138 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 5132 4984 5273 5012
rect 5132 4972 5138 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5261 4975 5319 4981
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 9732 4984 11529 5012
rect 9732 4972 9738 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 12268 5012 12296 5052
rect 12621 5083 12679 5089
rect 12621 5049 12633 5083
rect 12667 5080 12679 5083
rect 24780 5080 24808 5120
rect 25317 5117 25329 5151
rect 25363 5148 25375 5151
rect 26878 5148 26884 5160
rect 25363 5120 26884 5148
rect 25363 5117 25375 5120
rect 25317 5111 25375 5117
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 27522 5148 27528 5160
rect 27483 5120 27528 5148
rect 27522 5108 27528 5120
rect 27580 5108 27586 5160
rect 29641 5151 29699 5157
rect 29641 5117 29653 5151
rect 29687 5148 29699 5151
rect 30098 5148 30104 5160
rect 29687 5120 30104 5148
rect 29687 5117 29699 5120
rect 29641 5111 29699 5117
rect 30098 5108 30104 5120
rect 30156 5108 30162 5160
rect 30374 5108 30380 5160
rect 30432 5148 30438 5160
rect 30745 5151 30803 5157
rect 30745 5148 30757 5151
rect 30432 5120 30757 5148
rect 30432 5108 30438 5120
rect 30745 5117 30757 5120
rect 30791 5117 30803 5151
rect 31726 5148 31754 5188
rect 31864 5148 31892 5256
rect 33597 5253 33609 5256
rect 33643 5253 33655 5287
rect 34514 5284 34520 5296
rect 33597 5247 33655 5253
rect 33704 5256 34520 5284
rect 31938 5176 31944 5228
rect 31996 5216 32002 5228
rect 32769 5219 32827 5225
rect 32769 5216 32781 5219
rect 31996 5188 32781 5216
rect 31996 5176 32002 5188
rect 32769 5185 32781 5188
rect 32815 5185 32827 5219
rect 32769 5179 32827 5185
rect 32953 5219 33011 5225
rect 32953 5185 32965 5219
rect 32999 5185 33011 5219
rect 32953 5179 33011 5185
rect 31726 5120 31892 5148
rect 32968 5148 32996 5179
rect 33318 5176 33324 5228
rect 33376 5216 33382 5228
rect 33704 5225 33732 5256
rect 34514 5244 34520 5256
rect 34572 5244 34578 5296
rect 33413 5219 33471 5225
rect 33413 5216 33425 5219
rect 33376 5188 33425 5216
rect 33376 5176 33382 5188
rect 33413 5185 33425 5188
rect 33459 5185 33471 5219
rect 33413 5179 33471 5185
rect 33689 5219 33747 5225
rect 33689 5185 33701 5219
rect 33735 5185 33747 5219
rect 34146 5216 34152 5228
rect 34107 5188 34152 5216
rect 33689 5179 33747 5185
rect 34146 5176 34152 5188
rect 34204 5176 34210 5228
rect 33134 5148 33140 5160
rect 32968 5120 33140 5148
rect 30745 5111 30803 5117
rect 33134 5108 33140 5120
rect 33192 5148 33198 5160
rect 34164 5148 34192 5176
rect 33192 5120 34192 5148
rect 33192 5108 33198 5120
rect 26973 5083 27031 5089
rect 26973 5080 26985 5083
rect 12667 5052 22094 5080
rect 12667 5049 12679 5052
rect 12621 5043 12679 5049
rect 12636 5012 12664 5043
rect 12268 4984 12664 5012
rect 13081 5015 13139 5021
rect 11517 4975 11575 4981
rect 13081 4981 13093 5015
rect 13127 5012 13139 5015
rect 13170 5012 13176 5024
rect 13127 4984 13176 5012
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 13170 4972 13176 4984
rect 13228 4972 13234 5024
rect 15749 5015 15807 5021
rect 15749 4981 15761 5015
rect 15795 5012 15807 5015
rect 15930 5012 15936 5024
rect 15795 4984 15936 5012
rect 15795 4981 15807 4984
rect 15749 4975 15807 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 19426 5012 19432 5024
rect 19387 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20533 5015 20591 5021
rect 20533 4981 20545 5015
rect 20579 5012 20591 5015
rect 21266 5012 21272 5024
rect 20579 4984 21272 5012
rect 20579 4981 20591 4984
rect 20533 4975 20591 4981
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 22066 5012 22094 5052
rect 23768 5052 24716 5080
rect 24780 5052 26985 5080
rect 23768 5012 23796 5052
rect 22066 4984 23796 5012
rect 23845 5015 23903 5021
rect 23845 4981 23857 5015
rect 23891 5012 23903 5015
rect 24578 5012 24584 5024
rect 23891 4984 24584 5012
rect 23891 4981 23903 4984
rect 23845 4975 23903 4981
rect 24578 4972 24584 4984
rect 24636 4972 24642 5024
rect 24688 5012 24716 5052
rect 26973 5049 26985 5052
rect 27019 5049 27031 5083
rect 26973 5043 27031 5049
rect 29549 5083 29607 5089
rect 29549 5049 29561 5083
rect 29595 5080 29607 5083
rect 30653 5083 30711 5089
rect 30653 5080 30665 5083
rect 29595 5052 30665 5080
rect 29595 5049 29607 5052
rect 29549 5043 29607 5049
rect 30653 5049 30665 5052
rect 30699 5080 30711 5083
rect 33686 5080 33692 5092
rect 30699 5052 33692 5080
rect 30699 5049 30711 5052
rect 30653 5043 30711 5049
rect 33686 5040 33692 5052
rect 33744 5040 33750 5092
rect 28350 5012 28356 5024
rect 24688 4984 28356 5012
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 28442 4972 28448 5024
rect 28500 5012 28506 5024
rect 28997 5015 29055 5021
rect 28997 5012 29009 5015
rect 28500 4984 29009 5012
rect 28500 4972 28506 4984
rect 28997 4981 29009 4984
rect 29043 4981 29055 5015
rect 28997 4975 29055 4981
rect 29730 4972 29736 5024
rect 29788 5012 29794 5024
rect 30101 5015 30159 5021
rect 30101 5012 30113 5015
rect 29788 4984 30113 5012
rect 29788 4972 29794 4984
rect 30101 4981 30113 4984
rect 30147 4981 30159 5015
rect 33410 5012 33416 5024
rect 33371 4984 33416 5012
rect 30101 4975 30159 4981
rect 33410 4972 33416 4984
rect 33468 4972 33474 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 16758 4808 16764 4820
rect 11940 4780 16620 4808
rect 16719 4780 16764 4808
rect 11940 4768 11946 4780
rect 16592 4740 16620 4780
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 20162 4768 20168 4820
rect 20220 4808 20226 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20220 4780 20637 4808
rect 20220 4768 20226 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 23477 4811 23535 4817
rect 23477 4777 23489 4811
rect 23523 4808 23535 4811
rect 23566 4808 23572 4820
rect 23523 4780 23572 4808
rect 23523 4777 23535 4780
rect 23477 4771 23535 4777
rect 23566 4768 23572 4780
rect 23624 4768 23630 4820
rect 25317 4811 25375 4817
rect 25317 4808 25329 4811
rect 24780 4780 25329 4808
rect 19058 4740 19064 4752
rect 16592 4712 19064 4740
rect 19058 4700 19064 4712
rect 19116 4700 19122 4752
rect 20254 4700 20260 4752
rect 20312 4740 20318 4752
rect 24780 4740 24808 4780
rect 25317 4777 25329 4780
rect 25363 4808 25375 4811
rect 25774 4808 25780 4820
rect 25363 4780 25780 4808
rect 25363 4777 25375 4780
rect 25317 4771 25375 4777
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26878 4808 26884 4820
rect 26839 4780 26884 4808
rect 26878 4768 26884 4780
rect 26936 4768 26942 4820
rect 28905 4811 28963 4817
rect 28905 4808 28917 4811
rect 28276 4780 28917 4808
rect 28276 4740 28304 4780
rect 28905 4777 28917 4780
rect 28951 4808 28963 4811
rect 34146 4808 34152 4820
rect 28951 4780 33732 4808
rect 34107 4780 34152 4808
rect 28951 4777 28963 4780
rect 28905 4771 28963 4777
rect 20312 4712 24808 4740
rect 20312 4700 20318 4712
rect 5074 4672 5080 4684
rect 5035 4644 5080 4672
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 6733 4675 6791 4681
rect 6733 4641 6745 4675
rect 6779 4672 6791 4675
rect 9582 4672 9588 4684
rect 6779 4644 9588 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 10520 4644 12541 4672
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4614 4604 4620 4616
rect 4295 4576 4620 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 9674 4604 9680 4616
rect 9635 4576 9680 4604
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10520 4613 10548 4644
rect 12529 4641 12541 4644
rect 12575 4672 12587 4675
rect 13262 4672 13268 4684
rect 12575 4644 13268 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 22554 4672 22560 4684
rect 13924 4644 15516 4672
rect 22515 4644 22560 4672
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 10652 4576 10697 4604
rect 10652 4564 10658 4576
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 10873 4607 10931 4613
rect 10873 4604 10885 4607
rect 10836 4576 10885 4604
rect 10836 4564 10842 4576
rect 10873 4573 10885 4576
rect 10919 4604 10931 4607
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 10919 4576 11437 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 11425 4573 11437 4576
rect 11471 4604 11483 4607
rect 12342 4604 12348 4616
rect 11471 4576 12020 4604
rect 12255 4576 12348 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 9033 4539 9091 4545
rect 9033 4505 9045 4539
rect 9079 4536 9091 4539
rect 9876 4536 9904 4564
rect 9079 4508 9904 4536
rect 10689 4539 10747 4545
rect 9079 4505 9091 4508
rect 9033 4499 9091 4505
rect 10689 4505 10701 4539
rect 10735 4536 10747 4539
rect 11882 4536 11888 4548
rect 10735 4508 11888 4536
rect 10735 4505 10747 4508
rect 10689 4499 10747 4505
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 11992 4536 12020 4576
rect 12342 4564 12348 4576
rect 12400 4604 12406 4616
rect 13924 4604 13952 4644
rect 12400 4576 13952 4604
rect 12400 4564 12406 4576
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 15102 4604 15108 4616
rect 14056 4576 15108 4604
rect 14056 4564 14062 4576
rect 15102 4564 15108 4576
rect 15160 4604 15166 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 15160 4576 15393 4604
rect 15160 4564 15166 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15488 4604 15516 4644
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 24780 4681 24808 4712
rect 27172 4712 28304 4740
rect 33704 4740 33732 4780
rect 34146 4768 34152 4780
rect 34204 4768 34210 4820
rect 34790 4740 34796 4752
rect 33704 4712 34796 4740
rect 24765 4675 24823 4681
rect 22848 4644 24716 4672
rect 17034 4604 17040 4616
rect 15488 4576 17040 4604
rect 15381 4567 15439 4573
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 19242 4604 19248 4616
rect 17972 4576 19248 4604
rect 15648 4539 15706 4545
rect 11992 4508 15608 4536
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 4614 4468 4620 4480
rect 4479 4440 4620 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 9493 4471 9551 4477
rect 9493 4468 9505 4471
rect 8444 4440 9505 4468
rect 8444 4428 8450 4440
rect 9493 4437 9505 4440
rect 9539 4437 9551 4471
rect 10318 4468 10324 4480
rect 10279 4440 10324 4468
rect 9493 4431 9551 4437
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 15580 4468 15608 4508
rect 15648 4505 15660 4539
rect 15694 4536 15706 4539
rect 15746 4536 15752 4548
rect 15694 4508 15752 4536
rect 15694 4505 15706 4508
rect 15648 4499 15706 4505
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 17972 4480 18000 4576
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 21266 4604 21272 4616
rect 21227 4576 21272 4604
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4604 21511 4607
rect 21913 4607 21971 4613
rect 21913 4604 21925 4607
rect 21499 4576 21925 4604
rect 21499 4573 21511 4576
rect 21453 4567 21511 4573
rect 21913 4573 21925 4576
rect 21959 4604 21971 4607
rect 22738 4604 22744 4616
rect 21959 4576 22600 4604
rect 22699 4576 22744 4604
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 19490 4539 19548 4545
rect 19490 4536 19502 4539
rect 19392 4508 19502 4536
rect 19392 4496 19398 4508
rect 19490 4505 19502 4508
rect 19536 4505 19548 4539
rect 19490 4499 19548 4505
rect 21361 4539 21419 4545
rect 21361 4505 21373 4539
rect 21407 4536 21419 4539
rect 22094 4536 22100 4548
rect 21407 4508 22100 4536
rect 21407 4505 21419 4508
rect 21361 4499 21419 4505
rect 22094 4496 22100 4508
rect 22152 4496 22158 4548
rect 22572 4536 22600 4576
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 22848 4536 22876 4644
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4604 22983 4607
rect 23569 4607 23627 4613
rect 23569 4604 23581 4607
rect 22971 4576 23581 4604
rect 22971 4573 22983 4576
rect 22925 4567 22983 4573
rect 23569 4573 23581 4576
rect 23615 4573 23627 4607
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 23569 4567 23627 4573
rect 22572 4508 22876 4536
rect 23584 4536 23612 4567
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 24688 4604 24716 4644
rect 24765 4641 24777 4675
rect 24811 4641 24823 4675
rect 24765 4635 24823 4641
rect 27172 4604 27200 4712
rect 27338 4672 27344 4684
rect 27299 4644 27344 4672
rect 27338 4632 27344 4644
rect 27396 4632 27402 4684
rect 27522 4672 27528 4684
rect 27483 4644 27528 4672
rect 27522 4632 27528 4644
rect 27580 4632 27586 4684
rect 24688 4576 27200 4604
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4604 27307 4607
rect 27614 4604 27620 4616
rect 27295 4576 27620 4604
rect 27295 4573 27307 4576
rect 27249 4567 27307 4573
rect 27614 4564 27620 4576
rect 27672 4564 27678 4616
rect 28276 4613 28304 4712
rect 34790 4700 34796 4712
rect 34848 4700 34854 4752
rect 30193 4675 30251 4681
rect 30193 4672 30205 4675
rect 29564 4644 30205 4672
rect 28261 4607 28319 4613
rect 28261 4573 28273 4607
rect 28307 4573 28319 4607
rect 28442 4604 28448 4616
rect 28403 4576 28448 4604
rect 28261 4567 28319 4573
rect 28442 4564 28448 4576
rect 28500 4564 28506 4616
rect 29178 4564 29184 4616
rect 29236 4604 29242 4616
rect 29564 4613 29592 4644
rect 30193 4641 30205 4644
rect 30239 4672 30251 4675
rect 31481 4675 31539 4681
rect 31481 4672 31493 4675
rect 30239 4644 31493 4672
rect 30239 4641 30251 4644
rect 30193 4635 30251 4641
rect 31481 4641 31493 4644
rect 31527 4672 31539 4675
rect 31527 4644 32076 4672
rect 31527 4641 31539 4644
rect 31481 4635 31539 4641
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29236 4576 29561 4604
rect 29236 4564 29242 4576
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29730 4604 29736 4616
rect 29691 4576 29736 4604
rect 29549 4567 29607 4573
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 32048 4613 32076 4644
rect 32033 4607 32091 4613
rect 32033 4573 32045 4607
rect 32079 4573 32091 4607
rect 32214 4604 32220 4616
rect 32175 4576 32220 4604
rect 32033 4567 32091 4573
rect 31938 4536 31944 4548
rect 23584 4508 31944 4536
rect 31938 4496 31944 4508
rect 31996 4496 32002 4548
rect 32048 4536 32076 4567
rect 32214 4564 32220 4576
rect 32272 4564 32278 4616
rect 32769 4607 32827 4613
rect 32769 4573 32781 4607
rect 32815 4604 32827 4607
rect 32858 4604 32864 4616
rect 32815 4576 32864 4604
rect 32815 4573 32827 4576
rect 32769 4567 32827 4573
rect 32858 4564 32864 4576
rect 32916 4564 32922 4616
rect 33036 4607 33094 4613
rect 33036 4573 33048 4607
rect 33082 4604 33094 4607
rect 33410 4604 33416 4616
rect 33082 4576 33416 4604
rect 33082 4573 33094 4576
rect 33036 4567 33094 4573
rect 33410 4564 33416 4576
rect 33468 4564 33474 4616
rect 33318 4536 33324 4548
rect 32048 4508 33324 4536
rect 33318 4496 33324 4508
rect 33376 4496 33382 4548
rect 17034 4468 17040 4480
rect 15580 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 17218 4468 17224 4480
rect 17179 4440 17224 4468
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17954 4468 17960 4480
rect 17915 4440 17960 4468
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 24394 4468 24400 4480
rect 24355 4440 24400 4468
rect 24394 4428 24400 4440
rect 24452 4428 24458 4480
rect 28350 4468 28356 4480
rect 28311 4440 28356 4468
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 29641 4471 29699 4477
rect 29641 4437 29653 4471
rect 29687 4468 29699 4471
rect 29730 4468 29736 4480
rect 29687 4440 29736 4468
rect 29687 4437 29699 4440
rect 29641 4431 29699 4437
rect 29730 4428 29736 4440
rect 29788 4428 29794 4480
rect 32122 4468 32128 4480
rect 32083 4440 32128 4468
rect 32122 4428 32128 4440
rect 32180 4428 32186 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 8294 4264 8300 4276
rect 8255 4236 8300 4264
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 15746 4264 15752 4276
rect 15707 4236 15752 4264
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 17034 4224 17040 4276
rect 17092 4264 17098 4276
rect 17092 4236 17356 4264
rect 17092 4224 17098 4236
rect 2866 4196 2872 4208
rect 2827 4168 2872 4196
rect 2866 4156 2872 4168
rect 2924 4156 2930 4208
rect 17120 4199 17178 4205
rect 15764 4168 16068 4196
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4128 1458 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1452 4100 2053 4128
rect 1452 4088 1458 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2682 4128 2688 4140
rect 2643 4100 2688 4128
rect 2041 4091 2099 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4948 4100 4997 4128
rect 4948 4088 4954 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 9398 4128 9404 4140
rect 9456 4137 9462 4140
rect 9368 4100 9404 4128
rect 4985 4091 5043 4097
rect 9398 4088 9404 4100
rect 9456 4091 9468 4137
rect 10318 4128 10324 4140
rect 10279 4100 10324 4128
rect 9456 4088 9462 4091
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12575 4100 13001 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 12989 4091 13047 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13403 4100 13921 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13909 4097 13921 4100
rect 13955 4128 13967 4131
rect 15764 4128 15792 4168
rect 15930 4128 15936 4140
rect 13955 4100 15792 4128
rect 15891 4100 15936 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 3878 4060 3884 4072
rect 3839 4032 3884 4060
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 9692 3992 9720 4023
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 9916 4032 10517 4060
rect 9916 4020 9922 4032
rect 10505 4029 10517 4032
rect 10551 4060 10563 4063
rect 10870 4060 10876 4072
rect 10551 4032 10876 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 10870 4020 10876 4032
rect 10928 4060 10934 4072
rect 13372 4060 13400 4091
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16040 4128 16068 4168
rect 17120 4165 17132 4199
rect 17166 4196 17178 4199
rect 17218 4196 17224 4208
rect 17166 4168 17224 4196
rect 17166 4165 17178 4168
rect 17120 4159 17178 4165
rect 17218 4156 17224 4168
rect 17276 4156 17282 4208
rect 17328 4196 17356 4236
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 18233 4267 18291 4273
rect 18233 4264 18245 4267
rect 18104 4236 18245 4264
rect 18104 4224 18110 4236
rect 18233 4233 18245 4236
rect 18279 4233 18291 4267
rect 19334 4264 19340 4276
rect 19295 4236 19340 4264
rect 18233 4227 18291 4233
rect 19334 4224 19340 4236
rect 19392 4224 19398 4276
rect 22278 4224 22284 4276
rect 22336 4264 22342 4276
rect 23201 4267 23259 4273
rect 23201 4264 23213 4267
rect 22336 4236 23213 4264
rect 22336 4224 22342 4236
rect 23201 4233 23213 4236
rect 23247 4233 23259 4267
rect 27614 4264 27620 4276
rect 27575 4236 27620 4264
rect 23201 4227 23259 4233
rect 27614 4224 27620 4236
rect 27672 4224 27678 4276
rect 30834 4264 30840 4276
rect 30795 4236 30840 4264
rect 30834 4224 30840 4236
rect 30892 4224 30898 4276
rect 32677 4267 32735 4273
rect 32677 4233 32689 4267
rect 32723 4264 32735 4267
rect 32858 4264 32864 4276
rect 32723 4236 32864 4264
rect 32723 4233 32735 4236
rect 32677 4227 32735 4233
rect 32858 4224 32864 4236
rect 32916 4224 32922 4276
rect 23658 4196 23664 4208
rect 17328 4168 23664 4196
rect 23658 4156 23664 4168
rect 23716 4156 23722 4208
rect 28350 4156 28356 4208
rect 28408 4196 28414 4208
rect 28730 4199 28788 4205
rect 28730 4196 28742 4199
rect 28408 4168 28742 4196
rect 28408 4156 28414 4168
rect 28730 4165 28742 4168
rect 28776 4165 28788 4199
rect 28730 4159 28788 4165
rect 18966 4128 18972 4140
rect 16040 4100 18972 4128
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4097 19211 4131
rect 19153 4091 19211 4097
rect 10928 4032 13400 4060
rect 10928 4020 10934 4032
rect 15102 4020 15108 4072
rect 15160 4060 15166 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 15160 4032 16865 4060
rect 15160 4020 15166 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 19168 4060 19196 4091
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 22094 4137 22100 4140
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 19300 4100 20729 4128
rect 19300 4088 19306 4100
rect 20717 4097 20729 4100
rect 20763 4128 20775 4131
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 20763 4100 21833 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 22088 4091 22100 4137
rect 22152 4128 22158 4140
rect 24394 4128 24400 4140
rect 22152 4100 22188 4128
rect 24355 4100 24400 4128
rect 19426 4060 19432 4072
rect 19168 4032 19432 4060
rect 16853 4023 16911 4029
rect 9692 3964 11652 3992
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2590 3924 2596 3936
rect 1627 3896 2596 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9692 3924 9720 3964
rect 11624 3936 11652 3964
rect 10134 3924 10140 3936
rect 8996 3896 9720 3924
rect 10095 3896 10140 3924
rect 8996 3884 9002 3896
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 11606 3924 11612 3936
rect 11567 3896 11612 3924
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 12345 3927 12403 3933
rect 12345 3893 12357 3927
rect 12391 3924 12403 3927
rect 12434 3924 12440 3936
rect 12391 3896 12440 3924
rect 12391 3893 12403 3896
rect 12345 3887 12403 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 16868 3924 16896 4023
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 17954 3924 17960 3936
rect 16868 3896 17960 3924
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 21836 3924 21864 4091
rect 22094 4088 22100 4091
rect 22152 4088 22158 4100
rect 24394 4088 24400 4100
rect 24452 4088 24458 4140
rect 29730 4137 29736 4140
rect 29724 4128 29736 4137
rect 29691 4100 29736 4128
rect 29724 4091 29736 4100
rect 29730 4088 29736 4091
rect 29788 4088 29794 4140
rect 23753 4063 23811 4069
rect 23753 4029 23765 4063
rect 23799 4060 23811 4063
rect 24854 4060 24860 4072
rect 23799 4032 24860 4060
rect 23799 4029 23811 4032
rect 23753 4023 23811 4029
rect 23768 3992 23796 4023
rect 24854 4020 24860 4032
rect 24912 4020 24918 4072
rect 28997 4063 29055 4069
rect 28997 4029 29009 4063
rect 29043 4060 29055 4063
rect 29454 4060 29460 4072
rect 29043 4032 29460 4060
rect 29043 4029 29055 4032
rect 28997 4023 29055 4029
rect 29454 4020 29460 4032
rect 29512 4020 29518 4072
rect 23124 3964 23796 3992
rect 23124 3924 23152 3964
rect 21836 3896 23152 3924
rect 24581 3927 24639 3933
rect 24581 3893 24593 3927
rect 24627 3924 24639 3927
rect 24670 3924 24676 3936
rect 24627 3896 24676 3924
rect 24627 3893 24639 3896
rect 24581 3887 24639 3893
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2498 3720 2504 3732
rect 2459 3692 2504 3720
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3476 3692 11008 3720
rect 3476 3680 3482 3692
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 4982 3652 4988 3664
rect 2915 3624 4988 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 8389 3655 8447 3661
rect 8389 3621 8401 3655
rect 8435 3652 8447 3655
rect 10321 3655 10379 3661
rect 8435 3624 8800 3652
rect 8435 3621 8447 3624
rect 8389 3615 8447 3621
rect 2590 3584 2596 3596
rect 2551 3556 2596 3584
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4706 3584 4712 3596
rect 4571 3556 4712 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 1636 3488 2513 3516
rect 1636 3476 1642 3488
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8386 3516 8392 3528
rect 8251 3488 8392 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 4706 3448 4712 3460
rect 4667 3420 4712 3448
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 6365 3451 6423 3457
rect 6365 3417 6377 3451
rect 6411 3448 6423 3451
rect 8772 3448 8800 3624
rect 10321 3621 10333 3655
rect 10367 3652 10379 3655
rect 10502 3652 10508 3664
rect 10367 3624 10508 3652
rect 10367 3621 10379 3624
rect 10321 3615 10379 3621
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 10870 3652 10876 3664
rect 10831 3624 10876 3652
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 8938 3584 8944 3596
rect 8899 3556 8944 3584
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9186 3451 9244 3457
rect 9186 3448 9198 3451
rect 6411 3420 6914 3448
rect 8772 3420 9198 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 6886 3380 6914 3420
rect 9186 3417 9198 3420
rect 9232 3417 9244 3451
rect 10980 3448 11008 3692
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 13998 3720 14004 3732
rect 11664 3692 14004 3720
rect 11664 3680 11670 3692
rect 12176 3593 12204 3692
rect 13998 3680 14004 3692
rect 14056 3720 14062 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 14056 3692 14105 3720
rect 14056 3680 14062 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 18012 3692 18337 3720
rect 18012 3680 18018 3692
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 24854 3720 24860 3732
rect 18325 3683 18383 3689
rect 24596 3692 24860 3720
rect 13354 3612 13360 3664
rect 13412 3652 13418 3664
rect 13541 3655 13599 3661
rect 13541 3652 13553 3655
rect 13412 3624 13553 3652
rect 13412 3612 13418 3624
rect 13541 3621 13553 3624
rect 13587 3621 13599 3655
rect 13541 3615 13599 3621
rect 24596 3593 24624 3692
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 25958 3720 25964 3732
rect 25919 3692 25964 3720
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 29454 3680 29460 3732
rect 29512 3720 29518 3732
rect 29549 3723 29607 3729
rect 29549 3720 29561 3723
rect 29512 3692 29561 3720
rect 29512 3680 29518 3692
rect 29549 3689 29561 3692
rect 29595 3720 29607 3723
rect 30101 3723 30159 3729
rect 30101 3720 30113 3723
rect 29595 3692 30113 3720
rect 29595 3689 29607 3692
rect 29549 3683 29607 3689
rect 30101 3689 30113 3692
rect 30147 3720 30159 3723
rect 31021 3723 31079 3729
rect 31021 3720 31033 3723
rect 30147 3692 31033 3720
rect 30147 3689 30159 3692
rect 30101 3683 30159 3689
rect 31021 3689 31033 3692
rect 31067 3689 31079 3723
rect 31021 3683 31079 3689
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 24581 3587 24639 3593
rect 24581 3553 24593 3587
rect 24627 3553 24639 3587
rect 31036 3584 31064 3683
rect 31938 3680 31944 3732
rect 31996 3720 32002 3732
rect 32953 3723 33011 3729
rect 32953 3720 32965 3723
rect 31996 3692 32965 3720
rect 31996 3680 32002 3692
rect 32953 3689 32965 3692
rect 32999 3689 33011 3723
rect 32953 3683 33011 3689
rect 31573 3587 31631 3593
rect 31573 3584 31585 3587
rect 31036 3556 31585 3584
rect 24581 3547 24639 3553
rect 31573 3553 31585 3556
rect 31619 3553 31631 3587
rect 31573 3547 31631 3553
rect 12434 3525 12440 3528
rect 12428 3479 12440 3525
rect 12492 3516 12498 3528
rect 12492 3488 12528 3516
rect 12434 3476 12440 3479
rect 12492 3476 12498 3488
rect 24670 3476 24676 3528
rect 24728 3516 24734 3528
rect 24837 3519 24895 3525
rect 24837 3516 24849 3519
rect 24728 3488 24849 3516
rect 24728 3476 24734 3488
rect 24837 3485 24849 3488
rect 24883 3485 24895 3519
rect 31588 3516 31616 3547
rect 32858 3516 32864 3528
rect 31588 3488 32864 3516
rect 24837 3479 24895 3485
rect 32858 3476 32864 3488
rect 32916 3476 32922 3528
rect 20530 3448 20536 3460
rect 10980 3420 20536 3448
rect 9186 3411 9244 3417
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 31840 3451 31898 3457
rect 31840 3417 31852 3451
rect 31886 3448 31898 3451
rect 32122 3448 32128 3460
rect 31886 3420 32128 3448
rect 31886 3417 31898 3420
rect 31840 3411 31898 3417
rect 32122 3408 32128 3420
rect 32180 3408 32186 3460
rect 10226 3380 10232 3392
rect 6886 3352 10232 3380
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 5166 3176 5172 3188
rect 2823 3148 5172 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 9309 3179 9367 3185
rect 9309 3145 9321 3179
rect 9355 3176 9367 3179
rect 9398 3176 9404 3188
rect 9355 3148 9404 3176
rect 9355 3145 9367 3148
rect 9309 3139 9367 3145
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 11606 3176 11612 3188
rect 10551 3148 11612 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 24489 3179 24547 3185
rect 24489 3145 24501 3179
rect 24535 3176 24547 3179
rect 24854 3176 24860 3188
rect 24535 3148 24860 3176
rect 24535 3145 24547 3148
rect 24489 3139 24547 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 10134 3040 10140 3052
rect 9539 3012 10140 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 1394 2836 1400 2848
rect 1355 2808 1400 2836
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 1854 2796 1860 2848
rect 1912 2836 1918 2848
rect 2041 2839 2099 2845
rect 2041 2836 2053 2839
rect 1912 2808 2053 2836
rect 1912 2796 1918 2808
rect 2041 2805 2053 2808
rect 2087 2805 2099 2839
rect 2041 2799 2099 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2498 2632 2504 2644
rect 2459 2604 2504 2632
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 2924 2604 3801 2632
rect 2924 2592 2930 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 5258 2564 5264 2576
rect 2087 2536 5264 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2774 2428 2780 2440
rect 2731 2400 2780 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2774 2388 2780 2400
rect 2832 2428 2838 2440
rect 3145 2431 3203 2437
rect 3145 2428 3157 2431
rect 2832 2400 3157 2428
rect 2832 2388 2838 2400
rect 3145 2397 3157 2400
rect 3191 2397 3203 2431
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 3145 2391 3203 2397
rect 3970 2388 3976 2400
rect 4028 2428 4034 2440
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 4028 2400 4445 2428
rect 4028 2388 4034 2400
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 37734 2388 37740 2440
rect 37792 2428 37798 2440
rect 37829 2431 37887 2437
rect 37829 2428 37841 2431
rect 37792 2400 37841 2428
rect 37792 2388 37798 2400
rect 37829 2397 37841 2400
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 38010 2292 38016 2304
rect 37971 2264 38016 2292
rect 38010 2252 38016 2264
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 3424 37408 3476 37460
rect 23940 37408 23992 37460
rect 38016 37451 38068 37460
rect 38016 37417 38025 37451
rect 38025 37417 38059 37451
rect 38059 37417 38068 37451
rect 38016 37408 38068 37417
rect 3240 37340 3292 37392
rect 13360 37340 13412 37392
rect 16764 37315 16816 37324
rect 16764 37281 16773 37315
rect 16773 37281 16807 37315
rect 16807 37281 16816 37315
rect 16764 37272 16816 37281
rect 22192 37204 22244 37256
rect 29920 37204 29972 37256
rect 29184 37068 29236 37120
rect 37648 37068 37700 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 29920 36907 29972 36916
rect 29920 36873 29929 36907
rect 29929 36873 29963 36907
rect 29963 36873 29972 36907
rect 29920 36864 29972 36873
rect 14372 36796 14424 36848
rect 22192 36771 22244 36780
rect 22192 36737 22201 36771
rect 22201 36737 22235 36771
rect 22235 36737 22244 36771
rect 22192 36728 22244 36737
rect 2320 36660 2372 36712
rect 2872 36703 2924 36712
rect 2872 36669 2881 36703
rect 2881 36669 2915 36703
rect 2915 36669 2924 36703
rect 2872 36660 2924 36669
rect 4160 36703 4212 36712
rect 4160 36669 4169 36703
rect 4169 36669 4203 36703
rect 4203 36669 4212 36703
rect 4160 36660 4212 36669
rect 4712 36660 4764 36712
rect 12900 36660 12952 36712
rect 13820 36703 13872 36712
rect 13820 36669 13829 36703
rect 13829 36669 13863 36703
rect 13863 36669 13872 36703
rect 13820 36660 13872 36669
rect 22376 36703 22428 36712
rect 22376 36669 22385 36703
rect 22385 36669 22419 36703
rect 22419 36669 22428 36703
rect 22376 36660 22428 36669
rect 22100 36592 22152 36644
rect 4620 36524 4672 36576
rect 8944 36524 8996 36576
rect 18696 36524 18748 36576
rect 25412 36524 25464 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2320 36363 2372 36372
rect 2320 36329 2329 36363
rect 2329 36329 2363 36363
rect 2363 36329 2372 36363
rect 2320 36320 2372 36329
rect 12900 36363 12952 36372
rect 12900 36329 12909 36363
rect 12909 36329 12943 36363
rect 12943 36329 12952 36363
rect 12900 36320 12952 36329
rect 3976 36252 4028 36304
rect 5540 36252 5592 36304
rect 4068 36184 4120 36236
rect 6920 36184 6972 36236
rect 2780 36159 2832 36168
rect 2780 36125 2789 36159
rect 2789 36125 2823 36159
rect 2823 36125 2832 36159
rect 2780 36116 2832 36125
rect 4988 36091 5040 36100
rect 4988 36057 4997 36091
rect 4997 36057 5031 36091
rect 5031 36057 5040 36091
rect 4988 36048 5040 36057
rect 5540 35980 5592 36032
rect 9588 36048 9640 36100
rect 18696 36227 18748 36236
rect 18696 36193 18705 36227
rect 18705 36193 18739 36227
rect 18739 36193 18748 36227
rect 18696 36184 18748 36193
rect 22100 36227 22152 36236
rect 22100 36193 22109 36227
rect 22109 36193 22143 36227
rect 22143 36193 22152 36227
rect 22100 36184 22152 36193
rect 23480 36184 23532 36236
rect 25412 36227 25464 36236
rect 25412 36193 25421 36227
rect 25421 36193 25455 36227
rect 25455 36193 25464 36227
rect 25412 36184 25464 36193
rect 13636 36116 13688 36168
rect 30932 36159 30984 36168
rect 30932 36125 30941 36159
rect 30941 36125 30975 36159
rect 30975 36125 30984 36159
rect 30932 36116 30984 36125
rect 13820 36048 13872 36100
rect 16856 36091 16908 36100
rect 16856 36057 16865 36091
rect 16865 36057 16899 36091
rect 16899 36057 16908 36091
rect 16856 36048 16908 36057
rect 19340 36048 19392 36100
rect 21824 36091 21876 36100
rect 21824 36057 21833 36091
rect 21833 36057 21867 36091
rect 21867 36057 21876 36091
rect 21824 36048 21876 36057
rect 25596 36091 25648 36100
rect 25596 36057 25605 36091
rect 25605 36057 25639 36091
rect 25639 36057 25648 36091
rect 25596 36048 25648 36057
rect 27252 36091 27304 36100
rect 27252 36057 27261 36091
rect 27261 36057 27295 36091
rect 27295 36057 27304 36091
rect 27252 36048 27304 36057
rect 30380 36048 30432 36100
rect 18420 35980 18472 36032
rect 29552 36023 29604 36032
rect 29552 35989 29561 36023
rect 29561 35989 29595 36023
rect 29595 35989 29604 36023
rect 29552 35980 29604 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 2780 35776 2832 35828
rect 4988 35819 5040 35828
rect 4988 35785 4997 35819
rect 4997 35785 5031 35819
rect 5031 35785 5040 35819
rect 4988 35776 5040 35785
rect 21824 35819 21876 35828
rect 21824 35785 21833 35819
rect 21833 35785 21867 35819
rect 21867 35785 21876 35819
rect 21824 35776 21876 35785
rect 30380 35776 30432 35828
rect 4712 35708 4764 35760
rect 5172 35683 5224 35692
rect 5172 35649 5181 35683
rect 5181 35649 5215 35683
rect 5215 35649 5224 35683
rect 5172 35640 5224 35649
rect 13636 35683 13688 35692
rect 13636 35649 13645 35683
rect 13645 35649 13679 35683
rect 13679 35649 13688 35683
rect 13636 35640 13688 35649
rect 2964 35572 3016 35624
rect 3148 35615 3200 35624
rect 3148 35581 3157 35615
rect 3157 35581 3191 35615
rect 3191 35581 3200 35615
rect 7288 35615 7340 35624
rect 3148 35572 3200 35581
rect 7288 35581 7297 35615
rect 7297 35581 7331 35615
rect 7331 35581 7340 35615
rect 7288 35572 7340 35581
rect 7564 35572 7616 35624
rect 11796 35615 11848 35624
rect 11796 35581 11805 35615
rect 11805 35581 11839 35615
rect 11839 35581 11848 35615
rect 11796 35572 11848 35581
rect 13452 35615 13504 35624
rect 13452 35581 13461 35615
rect 13461 35581 13495 35615
rect 13495 35581 13504 35615
rect 13452 35572 13504 35581
rect 16764 35683 16816 35692
rect 16764 35649 16773 35683
rect 16773 35649 16807 35683
rect 16807 35649 16816 35683
rect 16764 35640 16816 35649
rect 17132 35572 17184 35624
rect 22100 35708 22152 35760
rect 19340 35683 19392 35692
rect 19340 35649 19349 35683
rect 19349 35649 19383 35683
rect 19383 35649 19392 35683
rect 19340 35640 19392 35649
rect 21732 35640 21784 35692
rect 22468 35683 22520 35692
rect 22468 35649 22477 35683
rect 22477 35649 22511 35683
rect 22511 35649 22520 35683
rect 22468 35640 22520 35649
rect 23480 35683 23532 35692
rect 23480 35649 23489 35683
rect 23489 35649 23523 35683
rect 23523 35649 23532 35683
rect 23480 35640 23532 35649
rect 28448 35640 28500 35692
rect 29644 35640 29696 35692
rect 19064 35615 19116 35624
rect 19064 35581 19073 35615
rect 19073 35581 19107 35615
rect 19107 35581 19116 35615
rect 19064 35572 19116 35581
rect 23848 35572 23900 35624
rect 30932 35572 30984 35624
rect 32588 35572 32640 35624
rect 13544 35436 13596 35488
rect 15476 35479 15528 35488
rect 15476 35445 15485 35479
rect 15485 35445 15519 35479
rect 15519 35445 15528 35479
rect 15476 35436 15528 35445
rect 26240 35436 26292 35488
rect 27712 35479 27764 35488
rect 27712 35445 27721 35479
rect 27721 35445 27755 35479
rect 27755 35445 27764 35479
rect 27712 35436 27764 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 7288 35232 7340 35284
rect 19064 35232 19116 35284
rect 19524 35232 19576 35284
rect 21732 35275 21784 35284
rect 21732 35241 21741 35275
rect 21741 35241 21775 35275
rect 21775 35241 21784 35275
rect 21732 35232 21784 35241
rect 22376 35275 22428 35284
rect 22376 35241 22385 35275
rect 22385 35241 22419 35275
rect 22419 35241 22428 35275
rect 22376 35232 22428 35241
rect 28448 35275 28500 35284
rect 28448 35241 28457 35275
rect 28457 35241 28491 35275
rect 28491 35241 28500 35275
rect 28448 35232 28500 35241
rect 6920 35164 6972 35216
rect 2872 35096 2924 35148
rect 4620 35139 4672 35148
rect 4620 35105 4629 35139
rect 4629 35105 4663 35139
rect 4663 35105 4672 35139
rect 4620 35096 4672 35105
rect 5540 35139 5592 35148
rect 5540 35105 5549 35139
rect 5549 35105 5583 35139
rect 5583 35105 5592 35139
rect 5540 35096 5592 35105
rect 8944 35139 8996 35148
rect 8944 35105 8953 35139
rect 8953 35105 8987 35139
rect 8987 35105 8996 35139
rect 8944 35096 8996 35105
rect 11796 35139 11848 35148
rect 11796 35105 11805 35139
rect 11805 35105 11839 35139
rect 11839 35105 11848 35139
rect 11796 35096 11848 35105
rect 13544 35139 13596 35148
rect 13544 35105 13553 35139
rect 13553 35105 13587 35139
rect 13587 35105 13596 35139
rect 13544 35096 13596 35105
rect 14372 35139 14424 35148
rect 14372 35105 14381 35139
rect 14381 35105 14415 35139
rect 14415 35105 14424 35139
rect 14372 35096 14424 35105
rect 15476 35139 15528 35148
rect 15476 35105 15485 35139
rect 15485 35105 15519 35139
rect 15519 35105 15528 35139
rect 15476 35096 15528 35105
rect 16856 35139 16908 35148
rect 16856 35105 16865 35139
rect 16865 35105 16899 35139
rect 16899 35105 16908 35139
rect 16856 35096 16908 35105
rect 18420 35139 18472 35148
rect 18420 35105 18429 35139
rect 18429 35105 18463 35139
rect 18463 35105 18472 35139
rect 18420 35096 18472 35105
rect 20812 35164 20864 35216
rect 26240 35139 26292 35148
rect 26240 35105 26249 35139
rect 26249 35105 26283 35139
rect 26283 35105 26292 35139
rect 26240 35096 26292 35105
rect 3976 35071 4028 35080
rect 3976 35037 3985 35071
rect 3985 35037 4019 35071
rect 4019 35037 4028 35071
rect 3976 35028 4028 35037
rect 14188 35028 14240 35080
rect 19984 35028 20036 35080
rect 22192 35071 22244 35080
rect 22192 35037 22201 35071
rect 22201 35037 22235 35071
rect 22235 35037 22244 35071
rect 22192 35028 22244 35037
rect 28356 35028 28408 35080
rect 4620 34960 4672 35012
rect 8576 34960 8628 35012
rect 13268 34960 13320 35012
rect 15660 35003 15712 35012
rect 15660 34969 15669 35003
rect 15669 34969 15703 35003
rect 15703 34969 15712 35003
rect 15660 34960 15712 34969
rect 20720 34960 20772 35012
rect 23848 34960 23900 35012
rect 25044 34960 25096 35012
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 3976 34688 4028 34740
rect 7564 34731 7616 34740
rect 7564 34697 7573 34731
rect 7573 34697 7607 34731
rect 7607 34697 7616 34731
rect 7564 34688 7616 34697
rect 8576 34731 8628 34740
rect 8576 34697 8585 34731
rect 8585 34697 8619 34731
rect 8619 34697 8628 34731
rect 8576 34688 8628 34697
rect 15660 34688 15712 34740
rect 3424 34620 3476 34672
rect 22468 34688 22520 34740
rect 28356 34731 28408 34740
rect 28356 34697 28365 34731
rect 28365 34697 28399 34731
rect 28399 34697 28408 34731
rect 28356 34688 28408 34697
rect 29644 34731 29696 34740
rect 29644 34697 29653 34731
rect 29653 34697 29687 34731
rect 29687 34697 29696 34731
rect 29644 34688 29696 34697
rect 2964 34552 3016 34604
rect 4896 34595 4948 34604
rect 4896 34561 4905 34595
rect 4905 34561 4939 34595
rect 4939 34561 4948 34595
rect 4896 34552 4948 34561
rect 5724 34552 5776 34604
rect 7380 34595 7432 34604
rect 7380 34561 7389 34595
rect 7389 34561 7423 34595
rect 7423 34561 7432 34595
rect 7380 34552 7432 34561
rect 8392 34595 8444 34604
rect 8392 34561 8401 34595
rect 8401 34561 8435 34595
rect 8435 34561 8444 34595
rect 8392 34552 8444 34561
rect 13268 34595 13320 34604
rect 13268 34561 13277 34595
rect 13277 34561 13311 34595
rect 13311 34561 13320 34595
rect 13268 34552 13320 34561
rect 13452 34552 13504 34604
rect 4068 34484 4120 34536
rect 4988 34527 5040 34536
rect 4988 34493 4997 34527
rect 4997 34493 5031 34527
rect 5031 34493 5040 34527
rect 4988 34484 5040 34493
rect 9036 34527 9088 34536
rect 9036 34493 9045 34527
rect 9045 34493 9079 34527
rect 9079 34493 9088 34527
rect 9036 34484 9088 34493
rect 9220 34527 9272 34536
rect 9220 34493 9229 34527
rect 9229 34493 9263 34527
rect 9263 34493 9272 34527
rect 9220 34484 9272 34493
rect 15200 34552 15252 34604
rect 15384 34595 15436 34604
rect 15384 34561 15393 34595
rect 15393 34561 15427 34595
rect 15427 34561 15436 34595
rect 15384 34552 15436 34561
rect 15660 34484 15712 34536
rect 19984 34620 20036 34672
rect 17960 34552 18012 34604
rect 20720 34595 20772 34604
rect 20720 34561 20729 34595
rect 20729 34561 20763 34595
rect 20763 34561 20772 34595
rect 20720 34552 20772 34561
rect 25044 34552 25096 34604
rect 25596 34552 25648 34604
rect 28540 34595 28592 34604
rect 28540 34561 28549 34595
rect 28549 34561 28583 34595
rect 28583 34561 28592 34595
rect 28540 34552 28592 34561
rect 29460 34595 29512 34604
rect 29460 34561 29469 34595
rect 29469 34561 29503 34595
rect 29503 34561 29512 34595
rect 29460 34552 29512 34561
rect 31300 34595 31352 34604
rect 31300 34561 31309 34595
rect 31309 34561 31343 34595
rect 31343 34561 31352 34595
rect 31300 34552 31352 34561
rect 18052 34527 18104 34536
rect 18052 34493 18061 34527
rect 18061 34493 18095 34527
rect 18095 34493 18104 34527
rect 18052 34484 18104 34493
rect 19248 34484 19300 34536
rect 20812 34527 20864 34536
rect 20812 34493 20821 34527
rect 20821 34493 20855 34527
rect 20855 34493 20864 34527
rect 20812 34484 20864 34493
rect 23020 34484 23072 34536
rect 24032 34484 24084 34536
rect 32036 34484 32088 34536
rect 4712 34348 4764 34400
rect 5540 34348 5592 34400
rect 5724 34391 5776 34400
rect 5724 34357 5733 34391
rect 5733 34357 5767 34391
rect 5767 34357 5776 34391
rect 5724 34348 5776 34357
rect 19340 34348 19392 34400
rect 20352 34348 20404 34400
rect 32312 34391 32364 34400
rect 32312 34357 32321 34391
rect 32321 34357 32355 34391
rect 32355 34357 32364 34391
rect 32312 34348 32364 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4712 34187 4764 34196
rect 4712 34153 4721 34187
rect 4721 34153 4755 34187
rect 4755 34153 4764 34187
rect 4712 34144 4764 34153
rect 5172 34144 5224 34196
rect 5540 34187 5592 34196
rect 5540 34153 5549 34187
rect 5549 34153 5583 34187
rect 5583 34153 5592 34187
rect 5540 34144 5592 34153
rect 9220 34144 9272 34196
rect 9588 34187 9640 34196
rect 9588 34153 9597 34187
rect 9597 34153 9631 34187
rect 9631 34153 9640 34187
rect 9588 34144 9640 34153
rect 15660 34187 15712 34196
rect 15660 34153 15669 34187
rect 15669 34153 15703 34187
rect 15703 34153 15712 34187
rect 15660 34144 15712 34153
rect 16396 34144 16448 34196
rect 19340 34144 19392 34196
rect 4620 34076 4672 34128
rect 17960 34076 18012 34128
rect 4988 34008 5040 34060
rect 16028 34051 16080 34060
rect 16028 34017 16037 34051
rect 16037 34017 16071 34051
rect 16071 34017 16080 34051
rect 16028 34008 16080 34017
rect 26332 34051 26384 34060
rect 26332 34017 26341 34051
rect 26341 34017 26375 34051
rect 26375 34017 26384 34051
rect 26332 34008 26384 34017
rect 27252 34008 27304 34060
rect 32588 34051 32640 34060
rect 32588 34017 32597 34051
rect 32597 34017 32631 34051
rect 32631 34017 32640 34051
rect 32588 34008 32640 34017
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 2412 33940 2464 33992
rect 3976 33983 4028 33992
rect 3976 33949 3985 33983
rect 3985 33949 4019 33983
rect 4019 33949 4028 33983
rect 3976 33940 4028 33949
rect 4620 33983 4672 33992
rect 4620 33949 4629 33983
rect 4629 33949 4663 33983
rect 4663 33949 4672 33983
rect 4620 33940 4672 33949
rect 4896 33940 4948 33992
rect 8944 33983 8996 33992
rect 8944 33949 8953 33983
rect 8953 33949 8987 33983
rect 8987 33949 8996 33983
rect 8944 33940 8996 33949
rect 9772 33983 9824 33992
rect 9772 33949 9781 33983
rect 9781 33949 9815 33983
rect 9815 33949 9824 33983
rect 9772 33940 9824 33949
rect 14280 33940 14332 33992
rect 15844 33983 15896 33992
rect 15844 33949 15853 33983
rect 15853 33949 15887 33983
rect 15887 33949 15896 33983
rect 15844 33940 15896 33949
rect 18328 33983 18380 33992
rect 18328 33949 18337 33983
rect 18337 33949 18371 33983
rect 18371 33949 18380 33983
rect 18328 33940 18380 33949
rect 19984 33940 20036 33992
rect 25412 33983 25464 33992
rect 25412 33949 25421 33983
rect 25421 33949 25455 33983
rect 25455 33949 25464 33983
rect 25412 33940 25464 33949
rect 32312 33983 32364 33992
rect 32312 33949 32330 33983
rect 32330 33949 32364 33983
rect 32312 33940 32364 33949
rect 38108 33983 38160 33992
rect 38108 33949 38117 33983
rect 38117 33949 38151 33983
rect 38151 33949 38160 33983
rect 38108 33940 38160 33949
rect 16120 33915 16172 33924
rect 2504 33804 2556 33856
rect 2596 33804 2648 33856
rect 5724 33804 5776 33856
rect 16120 33881 16129 33915
rect 16129 33881 16163 33915
rect 16163 33881 16172 33915
rect 16120 33872 16172 33881
rect 25596 33915 25648 33924
rect 25596 33881 25605 33915
rect 25605 33881 25639 33915
rect 25639 33881 25648 33915
rect 25596 33872 25648 33881
rect 28632 33872 28684 33924
rect 8760 33804 8812 33856
rect 29736 33804 29788 33856
rect 35348 33872 35400 33924
rect 30932 33804 30984 33856
rect 31208 33847 31260 33856
rect 31208 33813 31217 33847
rect 31217 33813 31251 33847
rect 31251 33813 31260 33847
rect 31208 33804 31260 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 3976 33600 4028 33652
rect 5724 33643 5776 33652
rect 5724 33609 5733 33643
rect 5733 33609 5767 33643
rect 5767 33609 5776 33643
rect 5724 33600 5776 33609
rect 24032 33600 24084 33652
rect 28540 33600 28592 33652
rect 29460 33600 29512 33652
rect 1400 33575 1452 33584
rect 1400 33541 1409 33575
rect 1409 33541 1443 33575
rect 1443 33541 1452 33575
rect 1400 33532 1452 33541
rect 2596 33575 2648 33584
rect 2596 33541 2605 33575
rect 2605 33541 2639 33575
rect 2639 33541 2648 33575
rect 2596 33532 2648 33541
rect 2412 33507 2464 33516
rect 2412 33473 2421 33507
rect 2421 33473 2455 33507
rect 2455 33473 2464 33507
rect 2412 33464 2464 33473
rect 4988 33464 5040 33516
rect 5264 33464 5316 33516
rect 9036 33507 9088 33516
rect 9036 33473 9045 33507
rect 9045 33473 9079 33507
rect 9079 33473 9088 33507
rect 9036 33464 9088 33473
rect 14280 33507 14332 33516
rect 14280 33473 14289 33507
rect 14289 33473 14323 33507
rect 14323 33473 14332 33507
rect 20720 33532 20772 33584
rect 27712 33532 27764 33584
rect 14280 33464 14332 33473
rect 18052 33464 18104 33516
rect 20352 33507 20404 33516
rect 20352 33473 20361 33507
rect 20361 33473 20395 33507
rect 20395 33473 20404 33507
rect 20352 33464 20404 33473
rect 22928 33507 22980 33516
rect 22928 33473 22937 33507
rect 22937 33473 22971 33507
rect 22971 33473 22980 33507
rect 22928 33464 22980 33473
rect 25412 33507 25464 33516
rect 25412 33473 25421 33507
rect 25421 33473 25455 33507
rect 25455 33473 25464 33507
rect 25412 33464 25464 33473
rect 28632 33575 28684 33584
rect 28632 33541 28641 33575
rect 28641 33541 28675 33575
rect 28675 33541 28684 33575
rect 29552 33575 29604 33584
rect 28632 33532 28684 33541
rect 29552 33541 29561 33575
rect 29561 33541 29595 33575
rect 29595 33541 29604 33575
rect 29552 33532 29604 33541
rect 30932 33575 30984 33584
rect 30932 33541 30941 33575
rect 30941 33541 30975 33575
rect 30975 33541 30984 33575
rect 30932 33532 30984 33541
rect 31116 33600 31168 33652
rect 31300 33643 31352 33652
rect 31300 33609 31309 33643
rect 31309 33609 31343 33643
rect 31343 33609 31352 33643
rect 31300 33600 31352 33609
rect 28816 33507 28868 33516
rect 2872 33439 2924 33448
rect 2872 33405 2881 33439
rect 2881 33405 2915 33439
rect 2915 33405 2924 33439
rect 2872 33396 2924 33405
rect 4620 33396 4672 33448
rect 5356 33396 5408 33448
rect 12440 33439 12492 33448
rect 12440 33405 12449 33439
rect 12449 33405 12483 33439
rect 12483 33405 12492 33439
rect 12440 33396 12492 33405
rect 16580 33396 16632 33448
rect 6092 33328 6144 33380
rect 20352 33328 20404 33380
rect 20812 33396 20864 33448
rect 28816 33473 28825 33507
rect 28825 33473 28859 33507
rect 28859 33473 28868 33507
rect 28816 33464 28868 33473
rect 29460 33507 29512 33516
rect 29460 33473 29469 33507
rect 29469 33473 29503 33507
rect 29503 33473 29512 33507
rect 29460 33464 29512 33473
rect 30748 33507 30800 33516
rect 29000 33396 29052 33448
rect 29736 33396 29788 33448
rect 30748 33473 30757 33507
rect 30757 33473 30791 33507
rect 30791 33473 30800 33507
rect 30748 33464 30800 33473
rect 29460 33328 29512 33380
rect 32496 33328 32548 33380
rect 5540 33260 5592 33312
rect 22836 33303 22888 33312
rect 22836 33269 22845 33303
rect 22845 33269 22879 33303
rect 22879 33269 22888 33303
rect 22836 33260 22888 33269
rect 28356 33260 28408 33312
rect 28816 33260 28868 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4068 33099 4120 33108
rect 4068 33065 4077 33099
rect 4077 33065 4111 33099
rect 4111 33065 4120 33099
rect 4068 33056 4120 33065
rect 5540 33056 5592 33108
rect 8392 33099 8444 33108
rect 8392 33065 8401 33099
rect 8401 33065 8435 33099
rect 8435 33065 8444 33099
rect 8392 33056 8444 33065
rect 8944 33099 8996 33108
rect 8944 33065 8953 33099
rect 8953 33065 8987 33099
rect 8987 33065 8996 33099
rect 8944 33056 8996 33065
rect 16580 33099 16632 33108
rect 8208 32988 8260 33040
rect 16580 33065 16589 33099
rect 16589 33065 16623 33099
rect 16623 33065 16632 33099
rect 16580 33056 16632 33065
rect 19984 33099 20036 33108
rect 5356 32920 5408 32972
rect 8392 32920 8444 32972
rect 14832 32920 14884 32972
rect 15844 32988 15896 33040
rect 16304 32988 16356 33040
rect 16396 32988 16448 33040
rect 19984 33065 19993 33099
rect 19993 33065 20027 33099
rect 20027 33065 20036 33099
rect 19984 33056 20036 33065
rect 20812 33056 20864 33108
rect 22192 33056 22244 33108
rect 23020 33099 23072 33108
rect 22008 32988 22060 33040
rect 23020 33065 23029 33099
rect 23029 33065 23063 33099
rect 23063 33065 23072 33099
rect 23020 33056 23072 33065
rect 4988 32852 5040 32904
rect 5632 32895 5684 32904
rect 5632 32861 5641 32895
rect 5641 32861 5675 32895
rect 5675 32861 5684 32895
rect 5632 32852 5684 32861
rect 8484 32852 8536 32904
rect 5264 32784 5316 32836
rect 8116 32784 8168 32836
rect 14096 32852 14148 32904
rect 16028 32963 16080 32972
rect 16028 32929 16037 32963
rect 16037 32929 16071 32963
rect 16071 32929 16080 32963
rect 16028 32920 16080 32929
rect 18328 32920 18380 32972
rect 21732 32963 21784 32972
rect 16120 32895 16172 32904
rect 16120 32861 16129 32895
rect 16129 32861 16163 32895
rect 16163 32861 16172 32895
rect 16120 32852 16172 32861
rect 16304 32852 16356 32904
rect 18972 32852 19024 32904
rect 19156 32852 19208 32904
rect 20444 32895 20496 32904
rect 20444 32861 20453 32895
rect 20453 32861 20487 32895
rect 20487 32861 20496 32895
rect 20444 32852 20496 32861
rect 21732 32929 21741 32963
rect 21741 32929 21775 32963
rect 21775 32929 21784 32963
rect 21732 32920 21784 32929
rect 27712 32920 27764 32972
rect 28356 32963 28408 32972
rect 28356 32929 28365 32963
rect 28365 32929 28399 32963
rect 28399 32929 28408 32963
rect 28356 32920 28408 32929
rect 14280 32784 14332 32836
rect 16488 32784 16540 32836
rect 23296 32852 23348 32904
rect 24860 32895 24912 32904
rect 24860 32861 24869 32895
rect 24869 32861 24903 32895
rect 24903 32861 24912 32895
rect 24860 32852 24912 32861
rect 22376 32784 22428 32836
rect 23112 32784 23164 32836
rect 25320 32784 25372 32836
rect 26700 32827 26752 32836
rect 26700 32793 26709 32827
rect 26709 32793 26743 32827
rect 26743 32793 26752 32827
rect 26700 32784 26752 32793
rect 27344 32827 27396 32836
rect 27344 32793 27353 32827
rect 27353 32793 27387 32827
rect 27387 32793 27396 32827
rect 27344 32784 27396 32793
rect 31024 32784 31076 32836
rect 30748 32716 30800 32768
rect 31576 32716 31628 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 5356 32555 5408 32564
rect 5356 32521 5365 32555
rect 5365 32521 5399 32555
rect 5399 32521 5408 32555
rect 5356 32512 5408 32521
rect 7380 32555 7432 32564
rect 7380 32521 7389 32555
rect 7389 32521 7423 32555
rect 7423 32521 7432 32555
rect 7380 32512 7432 32521
rect 9772 32512 9824 32564
rect 16488 32512 16540 32564
rect 18328 32555 18380 32564
rect 18328 32521 18337 32555
rect 18337 32521 18371 32555
rect 18371 32521 18380 32555
rect 18328 32512 18380 32521
rect 20720 32555 20772 32564
rect 20720 32521 20729 32555
rect 20729 32521 20763 32555
rect 20763 32521 20772 32555
rect 20720 32512 20772 32521
rect 22008 32555 22060 32564
rect 22008 32521 22017 32555
rect 22017 32521 22051 32555
rect 22051 32521 22060 32555
rect 22008 32512 22060 32521
rect 25320 32555 25372 32564
rect 7288 32444 7340 32496
rect 8116 32444 8168 32496
rect 14096 32487 14148 32496
rect 14096 32453 14105 32487
rect 14105 32453 14139 32487
rect 14139 32453 14148 32487
rect 14096 32444 14148 32453
rect 14832 32444 14884 32496
rect 21732 32444 21784 32496
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 5172 32419 5224 32428
rect 5172 32385 5181 32419
rect 5181 32385 5215 32419
rect 5215 32385 5224 32419
rect 5172 32376 5224 32385
rect 8484 32419 8536 32428
rect 6276 32308 6328 32360
rect 6184 32240 6236 32292
rect 8484 32385 8493 32419
rect 8493 32385 8527 32419
rect 8527 32385 8536 32419
rect 8484 32376 8536 32385
rect 14280 32419 14332 32428
rect 14280 32385 14289 32419
rect 14289 32385 14323 32419
rect 14323 32385 14332 32419
rect 14280 32376 14332 32385
rect 17776 32376 17828 32428
rect 19156 32419 19208 32428
rect 8392 32351 8444 32360
rect 8392 32317 8401 32351
rect 8401 32317 8435 32351
rect 8435 32317 8444 32351
rect 8392 32308 8444 32317
rect 12716 32351 12768 32360
rect 12716 32317 12725 32351
rect 12725 32317 12759 32351
rect 12759 32317 12768 32351
rect 12716 32308 12768 32317
rect 15292 32351 15344 32360
rect 15292 32317 15301 32351
rect 15301 32317 15335 32351
rect 15335 32317 15344 32351
rect 15292 32308 15344 32317
rect 15752 32308 15804 32360
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 20352 32376 20404 32428
rect 20536 32419 20588 32428
rect 20536 32385 20545 32419
rect 20545 32385 20579 32419
rect 20579 32385 20588 32419
rect 20536 32376 20588 32385
rect 20444 32308 20496 32360
rect 20352 32240 20404 32292
rect 23112 32376 23164 32428
rect 23296 32419 23348 32428
rect 23296 32385 23305 32419
rect 23305 32385 23339 32419
rect 23339 32385 23348 32419
rect 23296 32376 23348 32385
rect 25320 32521 25329 32555
rect 25329 32521 25363 32555
rect 25363 32521 25372 32555
rect 25320 32512 25372 32521
rect 24860 32444 24912 32496
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 29552 32444 29604 32496
rect 32404 32376 32456 32428
rect 32588 32376 32640 32428
rect 33324 32419 33376 32428
rect 33324 32385 33358 32419
rect 33358 32385 33376 32419
rect 33324 32376 33376 32385
rect 28632 32351 28684 32360
rect 22560 32240 22612 32292
rect 28632 32317 28641 32351
rect 28641 32317 28675 32351
rect 28675 32317 28684 32351
rect 28632 32308 28684 32317
rect 29000 32351 29052 32360
rect 29000 32317 29009 32351
rect 29009 32317 29043 32351
rect 29043 32317 29052 32351
rect 29000 32308 29052 32317
rect 32036 32308 32088 32360
rect 25596 32240 25648 32292
rect 1584 32215 1636 32224
rect 1584 32181 1593 32215
rect 1593 32181 1627 32215
rect 1627 32181 1636 32215
rect 1584 32172 1636 32181
rect 7196 32215 7248 32224
rect 7196 32181 7205 32215
rect 7205 32181 7239 32215
rect 7239 32181 7248 32215
rect 8208 32215 8260 32224
rect 7196 32172 7248 32181
rect 8208 32181 8217 32215
rect 8217 32181 8251 32215
rect 8251 32181 8260 32215
rect 8208 32172 8260 32181
rect 18972 32215 19024 32224
rect 18972 32181 18981 32215
rect 18981 32181 19015 32215
rect 19015 32181 19024 32215
rect 18972 32172 19024 32181
rect 19616 32215 19668 32224
rect 19616 32181 19625 32215
rect 19625 32181 19659 32215
rect 19659 32181 19668 32215
rect 19616 32172 19668 32181
rect 22008 32172 22060 32224
rect 23388 32172 23440 32224
rect 23940 32215 23992 32224
rect 23940 32181 23949 32215
rect 23949 32181 23983 32215
rect 23983 32181 23992 32215
rect 23940 32172 23992 32181
rect 33048 32172 33100 32224
rect 34428 32215 34480 32224
rect 34428 32181 34437 32215
rect 34437 32181 34471 32215
rect 34471 32181 34480 32215
rect 34428 32172 34480 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4988 32011 5040 32020
rect 4988 31977 4997 32011
rect 4997 31977 5031 32011
rect 5031 31977 5040 32011
rect 4988 31968 5040 31977
rect 15752 32011 15804 32020
rect 15752 31977 15761 32011
rect 15761 31977 15795 32011
rect 15795 31977 15804 32011
rect 15752 31968 15804 31977
rect 16396 31968 16448 32020
rect 19616 32011 19668 32020
rect 19616 31977 19625 32011
rect 19625 31977 19659 32011
rect 19659 31977 19668 32011
rect 19616 31968 19668 31977
rect 21916 31968 21968 32020
rect 23296 31968 23348 32020
rect 33324 31968 33376 32020
rect 8300 31900 8352 31952
rect 17776 31900 17828 31952
rect 20536 31900 20588 31952
rect 5632 31875 5684 31884
rect 5632 31841 5641 31875
rect 5641 31841 5675 31875
rect 5675 31841 5684 31875
rect 5632 31832 5684 31841
rect 6092 31875 6144 31884
rect 6092 31841 6101 31875
rect 6101 31841 6135 31875
rect 6135 31841 6144 31875
rect 12440 31875 12492 31884
rect 6092 31832 6144 31841
rect 12440 31841 12449 31875
rect 12449 31841 12483 31875
rect 12483 31841 12492 31875
rect 12440 31832 12492 31841
rect 13268 31832 13320 31884
rect 16028 31875 16080 31884
rect 16028 31841 16037 31875
rect 16037 31841 16071 31875
rect 16071 31841 16080 31875
rect 16028 31832 16080 31841
rect 13544 31807 13596 31816
rect 13544 31773 13553 31807
rect 13553 31773 13587 31807
rect 13587 31773 13596 31807
rect 13544 31764 13596 31773
rect 14924 31764 14976 31816
rect 16304 31832 16356 31884
rect 19984 31832 20036 31884
rect 16488 31764 16540 31816
rect 18972 31764 19024 31816
rect 22652 31832 22704 31884
rect 31208 31900 31260 31952
rect 30932 31875 30984 31884
rect 30932 31841 30941 31875
rect 30941 31841 30975 31875
rect 30975 31841 30984 31875
rect 30932 31832 30984 31841
rect 31576 31875 31628 31884
rect 31576 31841 31585 31875
rect 31585 31841 31619 31875
rect 31619 31841 31628 31875
rect 31576 31832 31628 31841
rect 5816 31739 5868 31748
rect 5816 31705 5825 31739
rect 5825 31705 5859 31739
rect 5859 31705 5868 31739
rect 5816 31696 5868 31705
rect 18696 31628 18748 31680
rect 22376 31764 22428 31816
rect 23020 31807 23072 31816
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 33048 31807 33100 31816
rect 33048 31773 33057 31807
rect 33057 31773 33091 31807
rect 33091 31773 33100 31807
rect 33048 31764 33100 31773
rect 22192 31628 22244 31680
rect 23112 31628 23164 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 5540 31467 5592 31476
rect 5540 31433 5549 31467
rect 5549 31433 5583 31467
rect 5583 31433 5592 31467
rect 5540 31424 5592 31433
rect 5816 31424 5868 31476
rect 19984 31424 20036 31476
rect 25504 31424 25556 31476
rect 32404 31424 32456 31476
rect 35348 31424 35400 31476
rect 1584 31356 1636 31408
rect 7288 31399 7340 31408
rect 7288 31365 7297 31399
rect 7297 31365 7331 31399
rect 7331 31365 7340 31399
rect 7288 31356 7340 31365
rect 15292 31356 15344 31408
rect 21732 31356 21784 31408
rect 23296 31356 23348 31408
rect 1400 31331 1452 31340
rect 1400 31297 1409 31331
rect 1409 31297 1443 31331
rect 1443 31297 1452 31331
rect 1400 31288 1452 31297
rect 2504 31220 2556 31272
rect 6368 31288 6420 31340
rect 7472 31331 7524 31340
rect 7472 31297 7481 31331
rect 7481 31297 7515 31331
rect 7515 31297 7524 31331
rect 7472 31288 7524 31297
rect 13544 31288 13596 31340
rect 14924 31331 14976 31340
rect 14924 31297 14933 31331
rect 14933 31297 14967 31331
rect 14967 31297 14976 31331
rect 14924 31288 14976 31297
rect 21456 31288 21508 31340
rect 22560 31331 22612 31340
rect 22560 31297 22569 31331
rect 22569 31297 22603 31331
rect 22603 31297 22612 31331
rect 22560 31288 22612 31297
rect 22836 31331 22888 31340
rect 22836 31297 22845 31331
rect 22845 31297 22879 31331
rect 22879 31297 22888 31331
rect 22836 31288 22888 31297
rect 23112 31288 23164 31340
rect 31024 31356 31076 31408
rect 31484 31356 31536 31408
rect 34428 31356 34480 31408
rect 27344 31288 27396 31340
rect 30932 31288 30984 31340
rect 32128 31331 32180 31340
rect 32128 31297 32137 31331
rect 32137 31297 32171 31331
rect 32171 31297 32180 31331
rect 32128 31288 32180 31297
rect 32404 31331 32456 31340
rect 32404 31297 32413 31331
rect 32413 31297 32447 31331
rect 32447 31297 32456 31331
rect 32404 31288 32456 31297
rect 32496 31331 32548 31340
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 7104 31220 7156 31272
rect 13084 31263 13136 31272
rect 13084 31229 13093 31263
rect 13093 31229 13127 31263
rect 13127 31229 13136 31263
rect 13084 31220 13136 31229
rect 23756 31220 23808 31272
rect 23940 31220 23992 31272
rect 26240 31220 26292 31272
rect 27620 31220 27672 31272
rect 31392 31152 31444 31204
rect 2504 31127 2556 31136
rect 2504 31093 2513 31127
rect 2513 31093 2547 31127
rect 2547 31093 2556 31127
rect 2504 31084 2556 31093
rect 2872 31084 2924 31136
rect 8944 31127 8996 31136
rect 8944 31093 8953 31127
rect 8953 31093 8987 31127
rect 8987 31093 8996 31127
rect 8944 31084 8996 31093
rect 21456 31084 21508 31136
rect 23388 31084 23440 31136
rect 24584 31084 24636 31136
rect 31484 31127 31536 31136
rect 31484 31093 31493 31127
rect 31493 31093 31527 31127
rect 31527 31093 31536 31127
rect 31484 31084 31536 31093
rect 35440 31084 35492 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6368 30923 6420 30932
rect 1400 30855 1452 30864
rect 1400 30821 1409 30855
rect 1409 30821 1443 30855
rect 1443 30821 1452 30855
rect 1400 30812 1452 30821
rect 6368 30889 6377 30923
rect 6377 30889 6411 30923
rect 6411 30889 6420 30923
rect 6368 30880 6420 30889
rect 19984 30880 20036 30932
rect 20812 30880 20864 30932
rect 7012 30812 7064 30864
rect 7196 30812 7248 30864
rect 5540 30744 5592 30796
rect 6276 30744 6328 30796
rect 8944 30787 8996 30796
rect 8944 30753 8953 30787
rect 8953 30753 8987 30787
rect 8987 30753 8996 30787
rect 8944 30744 8996 30753
rect 22008 30880 22060 30932
rect 25504 30880 25556 30932
rect 22100 30855 22152 30864
rect 22100 30821 22109 30855
rect 22109 30821 22143 30855
rect 22143 30821 22152 30855
rect 22100 30812 22152 30821
rect 23940 30812 23992 30864
rect 32128 30880 32180 30932
rect 25412 30744 25464 30796
rect 28632 30744 28684 30796
rect 2780 30719 2832 30728
rect 2780 30685 2789 30719
rect 2789 30685 2823 30719
rect 2823 30685 2832 30719
rect 2780 30676 2832 30685
rect 6184 30719 6236 30728
rect 6184 30685 6193 30719
rect 6193 30685 6227 30719
rect 6227 30685 6236 30719
rect 6184 30676 6236 30685
rect 14464 30676 14516 30728
rect 17592 30676 17644 30728
rect 18696 30719 18748 30728
rect 18696 30685 18705 30719
rect 18705 30685 18739 30719
rect 18739 30685 18748 30719
rect 18696 30676 18748 30685
rect 21916 30719 21968 30728
rect 21916 30685 21925 30719
rect 21925 30685 21959 30719
rect 21959 30685 21968 30719
rect 21916 30676 21968 30685
rect 5080 30608 5132 30660
rect 9128 30651 9180 30660
rect 9128 30617 9137 30651
rect 9137 30617 9171 30651
rect 9171 30617 9180 30651
rect 9128 30608 9180 30617
rect 3240 30540 3292 30592
rect 13084 30608 13136 30660
rect 22192 30676 22244 30728
rect 25780 30676 25832 30728
rect 25596 30651 25648 30660
rect 18512 30583 18564 30592
rect 18512 30549 18521 30583
rect 18521 30549 18555 30583
rect 18555 30549 18564 30583
rect 18512 30540 18564 30549
rect 21456 30540 21508 30592
rect 25596 30617 25605 30651
rect 25605 30617 25639 30651
rect 25639 30617 25648 30651
rect 25596 30608 25648 30617
rect 29368 30608 29420 30660
rect 32404 30744 32456 30796
rect 29644 30608 29696 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5080 30379 5132 30388
rect 5080 30345 5089 30379
rect 5089 30345 5123 30379
rect 5123 30345 5132 30379
rect 5080 30336 5132 30345
rect 18512 30268 18564 30320
rect 22100 30268 22152 30320
rect 25596 30268 25648 30320
rect 31392 30311 31444 30320
rect 31392 30277 31401 30311
rect 31401 30277 31435 30311
rect 31435 30277 31444 30311
rect 31392 30268 31444 30277
rect 2780 30243 2832 30252
rect 2780 30209 2789 30243
rect 2789 30209 2823 30243
rect 2823 30209 2832 30243
rect 2780 30200 2832 30209
rect 5080 30200 5132 30252
rect 7472 30200 7524 30252
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 17592 30243 17644 30252
rect 14464 30200 14516 30209
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 29644 30200 29696 30252
rect 30288 30200 30340 30252
rect 32588 30200 32640 30252
rect 34796 30268 34848 30320
rect 34060 30243 34112 30252
rect 34060 30209 34094 30243
rect 34094 30209 34112 30243
rect 34060 30200 34112 30209
rect 2964 30175 3016 30184
rect 2964 30141 2973 30175
rect 2973 30141 3007 30175
rect 3007 30141 3016 30175
rect 2964 30132 3016 30141
rect 3240 30175 3292 30184
rect 3240 30141 3249 30175
rect 3249 30141 3283 30175
rect 3283 30141 3292 30175
rect 3240 30132 3292 30141
rect 7012 30175 7064 30184
rect 7012 30141 7021 30175
rect 7021 30141 7055 30175
rect 7055 30141 7064 30175
rect 7012 30132 7064 30141
rect 7288 30175 7340 30184
rect 7288 30141 7297 30175
rect 7297 30141 7331 30175
rect 7331 30141 7340 30175
rect 7288 30132 7340 30141
rect 9404 30175 9456 30184
rect 8392 30064 8444 30116
rect 9404 30141 9413 30175
rect 9413 30141 9447 30175
rect 9447 30141 9456 30175
rect 9404 30132 9456 30141
rect 13084 30175 13136 30184
rect 13084 30141 13093 30175
rect 13093 30141 13127 30175
rect 13127 30141 13136 30175
rect 13084 30132 13136 30141
rect 14280 30175 14332 30184
rect 14280 30141 14289 30175
rect 14289 30141 14323 30175
rect 14323 30141 14332 30175
rect 14280 30132 14332 30141
rect 18236 30175 18288 30184
rect 18236 30141 18245 30175
rect 18245 30141 18279 30175
rect 18279 30141 18288 30175
rect 18236 30132 18288 30141
rect 22284 30132 22336 30184
rect 25412 30132 25464 30184
rect 28264 30175 28316 30184
rect 28264 30141 28273 30175
rect 28273 30141 28307 30175
rect 28307 30141 28316 30175
rect 28264 30132 28316 30141
rect 29276 30132 29328 30184
rect 26240 30064 26292 30116
rect 27620 30064 27672 30116
rect 3792 29996 3844 30048
rect 16672 30039 16724 30048
rect 16672 30005 16681 30039
rect 16681 30005 16715 30039
rect 16715 30005 16724 30039
rect 16672 29996 16724 30005
rect 22468 29996 22520 30048
rect 25228 29996 25280 30048
rect 25504 30039 25556 30048
rect 25504 30005 25513 30039
rect 25513 30005 25547 30039
rect 25547 30005 25556 30039
rect 25504 29996 25556 30005
rect 35348 29996 35400 30048
rect 38108 30039 38160 30048
rect 38108 30005 38117 30039
rect 38117 30005 38151 30039
rect 38151 30005 38160 30039
rect 38108 29996 38160 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2504 29792 2556 29844
rect 6184 29792 6236 29844
rect 9128 29835 9180 29844
rect 9128 29801 9137 29835
rect 9137 29801 9171 29835
rect 9171 29801 9180 29835
rect 9128 29792 9180 29801
rect 14188 29792 14240 29844
rect 15108 29792 15160 29844
rect 3792 29699 3844 29708
rect 3792 29665 3801 29699
rect 3801 29665 3835 29699
rect 3835 29665 3844 29699
rect 3792 29656 3844 29665
rect 4620 29699 4672 29708
rect 4620 29665 4629 29699
rect 4629 29665 4663 29699
rect 4663 29665 4672 29699
rect 4620 29656 4672 29665
rect 13268 29699 13320 29708
rect 13268 29665 13277 29699
rect 13277 29665 13311 29699
rect 13311 29665 13320 29699
rect 13268 29656 13320 29665
rect 15016 29656 15068 29708
rect 16672 29699 16724 29708
rect 16672 29665 16681 29699
rect 16681 29665 16715 29699
rect 16715 29665 16724 29699
rect 16672 29656 16724 29665
rect 19340 29656 19392 29708
rect 20720 29699 20772 29708
rect 20720 29665 20729 29699
rect 20729 29665 20763 29699
rect 20763 29665 20772 29699
rect 20720 29656 20772 29665
rect 22284 29699 22336 29708
rect 22284 29665 22293 29699
rect 22293 29665 22327 29699
rect 22327 29665 22336 29699
rect 22284 29656 22336 29665
rect 22468 29699 22520 29708
rect 22468 29665 22477 29699
rect 22477 29665 22511 29699
rect 22511 29665 22520 29699
rect 22468 29656 22520 29665
rect 25228 29699 25280 29708
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 26700 29699 26752 29708
rect 26700 29665 26709 29699
rect 26709 29665 26743 29699
rect 26743 29665 26752 29699
rect 26700 29656 26752 29665
rect 34796 29656 34848 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 3700 29588 3752 29640
rect 6644 29631 6696 29640
rect 6644 29597 6653 29631
rect 6653 29597 6687 29631
rect 6687 29597 6696 29631
rect 6644 29588 6696 29597
rect 8484 29588 8536 29640
rect 12256 29631 12308 29640
rect 8852 29520 8904 29572
rect 12256 29597 12265 29631
rect 12265 29597 12299 29631
rect 12299 29597 12308 29631
rect 12256 29588 12308 29597
rect 13728 29588 13780 29640
rect 14648 29631 14700 29640
rect 14648 29597 14657 29631
rect 14657 29597 14691 29631
rect 14691 29597 14700 29631
rect 14648 29588 14700 29597
rect 20536 29588 20588 29640
rect 22652 29588 22704 29640
rect 24492 29588 24544 29640
rect 14924 29563 14976 29572
rect 14924 29529 14933 29563
rect 14933 29529 14967 29563
rect 14967 29529 14976 29563
rect 14924 29520 14976 29529
rect 16856 29563 16908 29572
rect 16856 29529 16865 29563
rect 16865 29529 16899 29563
rect 16899 29529 16908 29563
rect 16856 29520 16908 29529
rect 4620 29452 4672 29504
rect 9404 29452 9456 29504
rect 12716 29452 12768 29504
rect 22836 29452 22888 29504
rect 36452 29520 36504 29572
rect 35808 29452 35860 29504
rect 37372 29452 37424 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 2964 29248 3016 29300
rect 8392 29291 8444 29300
rect 8392 29257 8401 29291
rect 8401 29257 8435 29291
rect 8435 29257 8444 29291
rect 8392 29248 8444 29257
rect 15384 29291 15436 29300
rect 15384 29257 15393 29291
rect 15393 29257 15427 29291
rect 15427 29257 15436 29291
rect 15384 29248 15436 29257
rect 16856 29291 16908 29300
rect 16856 29257 16865 29291
rect 16865 29257 16899 29291
rect 16899 29257 16908 29291
rect 16856 29248 16908 29257
rect 14924 29223 14976 29232
rect 14924 29189 14933 29223
rect 14933 29189 14967 29223
rect 14967 29189 14976 29223
rect 14924 29180 14976 29189
rect 16580 29180 16632 29232
rect 22836 29180 22888 29232
rect 23020 29248 23072 29300
rect 23664 29248 23716 29300
rect 24308 29248 24360 29300
rect 24492 29291 24544 29300
rect 24492 29257 24501 29291
rect 24501 29257 24535 29291
rect 24535 29257 24544 29291
rect 24492 29248 24544 29257
rect 29276 29291 29328 29300
rect 29276 29257 29285 29291
rect 29285 29257 29319 29291
rect 29319 29257 29328 29291
rect 29276 29248 29328 29257
rect 36452 29291 36504 29300
rect 28264 29180 28316 29232
rect 3240 29112 3292 29164
rect 8392 29112 8444 29164
rect 8852 29155 8904 29164
rect 8852 29121 8861 29155
rect 8861 29121 8895 29155
rect 8895 29121 8904 29155
rect 8852 29112 8904 29121
rect 12256 29155 12308 29164
rect 12256 29121 12265 29155
rect 12265 29121 12299 29155
rect 12299 29121 12308 29155
rect 12256 29112 12308 29121
rect 14648 29112 14700 29164
rect 15200 29155 15252 29164
rect 15200 29121 15209 29155
rect 15209 29121 15243 29155
rect 15243 29121 15252 29155
rect 15200 29112 15252 29121
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 20536 29155 20588 29164
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 22744 29155 22796 29164
rect 3516 29087 3568 29096
rect 3516 29053 3525 29087
rect 3525 29053 3559 29087
rect 3559 29053 3568 29087
rect 3516 29044 3568 29053
rect 3884 29087 3936 29096
rect 3884 29053 3893 29087
rect 3893 29053 3927 29087
rect 3927 29053 3936 29087
rect 9036 29087 9088 29096
rect 3884 29044 3936 29053
rect 9036 29053 9045 29087
rect 9045 29053 9079 29087
rect 9079 29053 9088 29087
rect 9036 29044 9088 29053
rect 12440 29087 12492 29096
rect 12440 29053 12449 29087
rect 12449 29053 12483 29087
rect 12483 29053 12492 29087
rect 12440 29044 12492 29053
rect 12716 29087 12768 29096
rect 12716 29053 12725 29087
rect 12725 29053 12759 29087
rect 12759 29053 12768 29087
rect 12716 29044 12768 29053
rect 15016 29087 15068 29096
rect 15016 29053 15025 29087
rect 15025 29053 15059 29087
rect 15059 29053 15068 29087
rect 15016 29044 15068 29053
rect 19340 29044 19392 29096
rect 20168 29044 20220 29096
rect 18236 28976 18288 29028
rect 19984 28976 20036 29028
rect 20444 28976 20496 29028
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 24308 29155 24360 29164
rect 24308 29121 24317 29155
rect 24317 29121 24351 29155
rect 24351 29121 24360 29155
rect 29092 29155 29144 29164
rect 24308 29112 24360 29121
rect 29092 29121 29101 29155
rect 29101 29121 29135 29155
rect 29135 29121 29144 29155
rect 29092 29112 29144 29121
rect 35348 29180 35400 29232
rect 35808 29155 35860 29164
rect 35808 29121 35817 29155
rect 35817 29121 35851 29155
rect 35851 29121 35860 29155
rect 35808 29112 35860 29121
rect 35992 29155 36044 29164
rect 35992 29121 36001 29155
rect 36001 29121 36035 29155
rect 36035 29121 36044 29155
rect 35992 29112 36044 29121
rect 36452 29257 36461 29291
rect 36461 29257 36495 29291
rect 36495 29257 36504 29291
rect 36452 29248 36504 29257
rect 25596 29044 25648 29096
rect 35900 29044 35952 29096
rect 37372 29112 37424 29164
rect 37004 29044 37056 29096
rect 25412 28976 25464 29028
rect 15108 28908 15160 28960
rect 15476 28908 15528 28960
rect 22100 28908 22152 28960
rect 23756 28908 23808 28960
rect 34704 28908 34756 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3516 28704 3568 28756
rect 3700 28704 3752 28756
rect 4712 28704 4764 28756
rect 7932 28747 7984 28756
rect 7932 28713 7941 28747
rect 7941 28713 7975 28747
rect 7975 28713 7984 28747
rect 7932 28704 7984 28713
rect 8392 28747 8444 28756
rect 8392 28713 8401 28747
rect 8401 28713 8435 28747
rect 8435 28713 8444 28747
rect 8392 28704 8444 28713
rect 9036 28704 9088 28756
rect 15476 28747 15528 28756
rect 15476 28713 15485 28747
rect 15485 28713 15519 28747
rect 15519 28713 15528 28747
rect 15476 28704 15528 28713
rect 29092 28704 29144 28756
rect 35992 28704 36044 28756
rect 15292 28636 15344 28688
rect 4068 28611 4120 28620
rect 4068 28577 4077 28611
rect 4077 28577 4111 28611
rect 4111 28577 4120 28611
rect 4068 28568 4120 28577
rect 5540 28568 5592 28620
rect 8024 28611 8076 28620
rect 8024 28577 8033 28611
rect 8033 28577 8067 28611
rect 8067 28577 8076 28611
rect 8024 28568 8076 28577
rect 12440 28568 12492 28620
rect 14280 28568 14332 28620
rect 14464 28568 14516 28620
rect 18236 28611 18288 28620
rect 18236 28577 18245 28611
rect 18245 28577 18279 28611
rect 18279 28577 18288 28611
rect 18236 28568 18288 28577
rect 20168 28611 20220 28620
rect 20168 28577 20177 28611
rect 20177 28577 20211 28611
rect 20211 28577 20220 28611
rect 20168 28568 20220 28577
rect 34796 28568 34848 28620
rect 37004 28568 37056 28620
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 3700 28500 3752 28552
rect 3884 28500 3936 28552
rect 4160 28500 4212 28552
rect 4988 28500 5040 28552
rect 5264 28500 5316 28552
rect 7840 28500 7892 28552
rect 8208 28543 8260 28552
rect 8208 28509 8217 28543
rect 8217 28509 8251 28543
rect 8251 28509 8260 28543
rect 8208 28500 8260 28509
rect 8944 28543 8996 28552
rect 8944 28509 8953 28543
rect 8953 28509 8987 28543
rect 8987 28509 8996 28543
rect 8944 28500 8996 28509
rect 13544 28543 13596 28552
rect 13544 28509 13553 28543
rect 13553 28509 13587 28543
rect 13587 28509 13596 28543
rect 13544 28500 13596 28509
rect 14096 28543 14148 28552
rect 14096 28509 14105 28543
rect 14105 28509 14139 28543
rect 14139 28509 14148 28543
rect 14096 28500 14148 28509
rect 15108 28500 15160 28552
rect 16856 28543 16908 28552
rect 16856 28509 16865 28543
rect 16865 28509 16899 28543
rect 16899 28509 16908 28543
rect 16856 28500 16908 28509
rect 20076 28500 20128 28552
rect 36452 28500 36504 28552
rect 37372 28543 37424 28552
rect 37372 28509 37381 28543
rect 37381 28509 37415 28543
rect 37415 28509 37424 28543
rect 37372 28500 37424 28509
rect 15384 28475 15436 28484
rect 15384 28441 15393 28475
rect 15393 28441 15427 28475
rect 15427 28441 15436 28475
rect 15384 28432 15436 28441
rect 17040 28475 17092 28484
rect 17040 28441 17049 28475
rect 17049 28441 17083 28475
rect 17083 28441 17092 28475
rect 17040 28432 17092 28441
rect 28080 28475 28132 28484
rect 28080 28441 28089 28475
rect 28089 28441 28123 28475
rect 28123 28441 28132 28475
rect 28080 28432 28132 28441
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 35624 28432 35676 28484
rect 29276 28364 29328 28416
rect 32312 28364 32364 28416
rect 35992 28364 36044 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3700 28203 3752 28212
rect 3700 28169 3709 28203
rect 3709 28169 3743 28203
rect 3743 28169 3752 28203
rect 3700 28160 3752 28169
rect 8484 28160 8536 28212
rect 13728 28203 13780 28212
rect 13728 28169 13737 28203
rect 13737 28169 13771 28203
rect 13771 28169 13780 28203
rect 13728 28160 13780 28169
rect 16672 28160 16724 28212
rect 20812 28160 20864 28212
rect 34060 28203 34112 28212
rect 34060 28169 34069 28203
rect 34069 28169 34103 28203
rect 34103 28169 34112 28203
rect 34060 28160 34112 28169
rect 4160 28135 4212 28144
rect 4160 28101 4169 28135
rect 4169 28101 4203 28135
rect 4203 28101 4212 28135
rect 4160 28092 4212 28101
rect 7840 28092 7892 28144
rect 8300 28092 8352 28144
rect 14372 28092 14424 28144
rect 15384 28092 15436 28144
rect 30288 28135 30340 28144
rect 3700 28024 3752 28076
rect 3884 28067 3936 28076
rect 3884 28033 3893 28067
rect 3893 28033 3927 28067
rect 3927 28033 3936 28067
rect 3884 28024 3936 28033
rect 4068 28024 4120 28076
rect 8208 28067 8260 28076
rect 8208 28033 8217 28067
rect 8217 28033 8251 28067
rect 8251 28033 8260 28067
rect 8208 28024 8260 28033
rect 15108 28067 15160 28076
rect 15108 28033 15117 28067
rect 15117 28033 15151 28067
rect 15151 28033 15160 28067
rect 15108 28024 15160 28033
rect 16856 28024 16908 28076
rect 30288 28101 30297 28135
rect 30297 28101 30331 28135
rect 30331 28101 30340 28135
rect 30288 28092 30340 28101
rect 34704 28092 34756 28144
rect 28172 28024 28224 28076
rect 30472 28067 30524 28076
rect 30472 28033 30481 28067
rect 30481 28033 30515 28067
rect 30515 28033 30524 28067
rect 30472 28024 30524 28033
rect 30932 28024 30984 28076
rect 8024 27999 8076 28008
rect 8024 27965 8033 27999
rect 8033 27965 8067 27999
rect 8067 27965 8076 27999
rect 8024 27956 8076 27965
rect 14464 27956 14516 28008
rect 14556 27956 14608 28008
rect 15016 27956 15068 28008
rect 3792 27888 3844 27940
rect 4804 27888 4856 27940
rect 20260 27888 20312 27940
rect 28632 27888 28684 27940
rect 31392 28067 31444 28076
rect 31392 28033 31401 28067
rect 31401 28033 31435 28067
rect 31435 28033 31444 28067
rect 32128 28067 32180 28076
rect 31392 28024 31444 28033
rect 32128 28033 32137 28067
rect 32137 28033 32171 28067
rect 32171 28033 32180 28067
rect 32128 28024 32180 28033
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 34244 28067 34296 28076
rect 34244 28033 34253 28067
rect 34253 28033 34287 28067
rect 34287 28033 34296 28067
rect 34244 28024 34296 28033
rect 35348 28024 35400 28076
rect 35532 28024 35584 28076
rect 36452 28067 36504 28076
rect 36452 28033 36461 28067
rect 36461 28033 36495 28067
rect 36495 28033 36504 28067
rect 36452 28024 36504 28033
rect 34520 27999 34572 28008
rect 34520 27965 34529 27999
rect 34529 27965 34563 27999
rect 34563 27965 34572 27999
rect 34520 27956 34572 27965
rect 4712 27820 4764 27872
rect 7932 27863 7984 27872
rect 7932 27829 7941 27863
rect 7941 27829 7975 27863
rect 7975 27829 7984 27863
rect 7932 27820 7984 27829
rect 15476 27820 15528 27872
rect 21824 27863 21876 27872
rect 21824 27829 21833 27863
rect 21833 27829 21867 27863
rect 21867 27829 21876 27863
rect 21824 27820 21876 27829
rect 34428 27863 34480 27872
rect 34428 27829 34437 27863
rect 34437 27829 34471 27863
rect 34471 27829 34480 27863
rect 34428 27820 34480 27829
rect 36268 27863 36320 27872
rect 36268 27829 36277 27863
rect 36277 27829 36311 27863
rect 36311 27829 36320 27863
rect 36268 27820 36320 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4712 27616 4764 27668
rect 7932 27659 7984 27668
rect 7932 27625 7941 27659
rect 7941 27625 7975 27659
rect 7975 27625 7984 27659
rect 7932 27616 7984 27625
rect 8944 27616 8996 27668
rect 14096 27659 14148 27668
rect 14096 27625 14105 27659
rect 14105 27625 14139 27659
rect 14139 27625 14148 27659
rect 14096 27616 14148 27625
rect 14188 27616 14240 27668
rect 20076 27659 20128 27668
rect 20076 27625 20085 27659
rect 20085 27625 20119 27659
rect 20119 27625 20128 27659
rect 20076 27616 20128 27625
rect 3240 27548 3292 27600
rect 3976 27548 4028 27600
rect 8024 27523 8076 27532
rect 8024 27489 8033 27523
rect 8033 27489 8067 27523
rect 8067 27489 8076 27523
rect 8024 27480 8076 27489
rect 3700 27412 3752 27464
rect 4160 27412 4212 27464
rect 4620 27412 4672 27464
rect 7104 27412 7156 27464
rect 7840 27412 7892 27464
rect 8208 27455 8260 27464
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 14280 27455 14332 27464
rect 14280 27421 14289 27455
rect 14289 27421 14323 27455
rect 14323 27421 14332 27455
rect 14280 27412 14332 27421
rect 14004 27344 14056 27396
rect 14464 27412 14516 27464
rect 15292 27412 15344 27464
rect 17040 27480 17092 27532
rect 20812 27616 20864 27668
rect 22008 27616 22060 27668
rect 28172 27659 28224 27668
rect 28172 27625 28181 27659
rect 28181 27625 28215 27659
rect 28215 27625 28224 27659
rect 28172 27616 28224 27625
rect 31392 27616 31444 27668
rect 34244 27616 34296 27668
rect 35624 27659 35676 27668
rect 35624 27625 35633 27659
rect 35633 27625 35667 27659
rect 35667 27625 35676 27659
rect 35624 27616 35676 27625
rect 22100 27548 22152 27600
rect 36268 27548 36320 27600
rect 20996 27480 21048 27532
rect 20260 27455 20312 27464
rect 20260 27421 20269 27455
rect 20269 27421 20303 27455
rect 20303 27421 20312 27455
rect 20260 27412 20312 27421
rect 20904 27412 20956 27464
rect 21088 27412 21140 27464
rect 22744 27480 22796 27532
rect 27068 27480 27120 27532
rect 22376 27455 22428 27464
rect 4712 27319 4764 27328
rect 4712 27285 4721 27319
rect 4721 27285 4755 27319
rect 4755 27285 4764 27319
rect 4712 27276 4764 27285
rect 5264 27276 5316 27328
rect 7288 27276 7340 27328
rect 14372 27276 14424 27328
rect 15568 27344 15620 27396
rect 20628 27344 20680 27396
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 22836 27455 22888 27464
rect 22836 27421 22845 27455
rect 22845 27421 22879 27455
rect 22879 27421 22888 27455
rect 22836 27412 22888 27421
rect 26056 27412 26108 27464
rect 27620 27344 27672 27396
rect 28632 27344 28684 27396
rect 32312 27412 32364 27464
rect 35532 27480 35584 27532
rect 34336 27412 34388 27464
rect 32128 27344 32180 27396
rect 35624 27412 35676 27464
rect 35808 27412 35860 27464
rect 22008 27276 22060 27328
rect 26976 27319 27028 27328
rect 26976 27285 26985 27319
rect 26985 27285 27019 27319
rect 27019 27285 27028 27319
rect 26976 27276 27028 27285
rect 27344 27319 27396 27328
rect 27344 27285 27353 27319
rect 27353 27285 27387 27319
rect 27387 27285 27396 27319
rect 27344 27276 27396 27285
rect 28356 27276 28408 27328
rect 29276 27276 29328 27328
rect 33324 27319 33376 27328
rect 33324 27285 33333 27319
rect 33333 27285 33367 27319
rect 33367 27285 33376 27319
rect 36268 27344 36320 27396
rect 33324 27276 33376 27285
rect 34520 27276 34572 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 5540 27072 5592 27124
rect 6644 27072 6696 27124
rect 8208 27072 8260 27124
rect 13544 27072 13596 27124
rect 7288 27004 7340 27056
rect 8300 27004 8352 27056
rect 8760 27004 8812 27056
rect 14372 27004 14424 27056
rect 7656 26936 7708 26988
rect 10048 26979 10100 26988
rect 10048 26945 10057 26979
rect 10057 26945 10091 26979
rect 10091 26945 10100 26979
rect 10048 26936 10100 26945
rect 14004 26911 14056 26920
rect 14004 26877 14013 26911
rect 14013 26877 14047 26911
rect 14047 26877 14056 26911
rect 14004 26868 14056 26877
rect 14740 26936 14792 26988
rect 15108 27072 15160 27124
rect 15476 27115 15528 27124
rect 15476 27081 15485 27115
rect 15485 27081 15519 27115
rect 15519 27081 15528 27115
rect 15476 27072 15528 27081
rect 26056 27115 26108 27124
rect 26056 27081 26065 27115
rect 26065 27081 26099 27115
rect 26099 27081 26108 27115
rect 26056 27072 26108 27081
rect 20628 27004 20680 27056
rect 22008 27047 22060 27056
rect 15660 26979 15712 26988
rect 14280 26868 14332 26920
rect 15016 26868 15068 26920
rect 7840 26800 7892 26852
rect 15108 26800 15160 26852
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 20168 26800 20220 26852
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 22008 27013 22017 27047
rect 22017 27013 22051 27047
rect 22051 27013 22060 27047
rect 22008 27004 22060 27013
rect 33324 27072 33376 27124
rect 34428 27072 34480 27124
rect 26976 27004 27028 27056
rect 30564 27004 30616 27056
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 23388 26936 23440 26988
rect 26332 26936 26384 26988
rect 29276 26936 29328 26988
rect 30288 26936 30340 26988
rect 33600 26936 33652 26988
rect 34336 26936 34388 26988
rect 34704 26979 34756 26988
rect 34704 26945 34713 26979
rect 34713 26945 34747 26979
rect 34747 26945 34756 26979
rect 34704 26936 34756 26945
rect 27160 26911 27212 26920
rect 27160 26877 27169 26911
rect 27169 26877 27203 26911
rect 27203 26877 27212 26911
rect 27160 26868 27212 26877
rect 27344 26868 27396 26920
rect 34428 26868 34480 26920
rect 35900 26936 35952 26988
rect 36268 26868 36320 26920
rect 27620 26800 27672 26852
rect 35532 26800 35584 26852
rect 2780 26732 2832 26784
rect 3700 26732 3752 26784
rect 10600 26732 10652 26784
rect 10784 26732 10836 26784
rect 14188 26775 14240 26784
rect 14188 26741 14197 26775
rect 14197 26741 14231 26775
rect 14231 26741 14240 26775
rect 14188 26732 14240 26741
rect 20812 26775 20864 26784
rect 20812 26741 20821 26775
rect 20821 26741 20855 26775
rect 20855 26741 20864 26775
rect 20812 26732 20864 26741
rect 21732 26732 21784 26784
rect 30380 26732 30432 26784
rect 30932 26732 30984 26784
rect 33600 26775 33652 26784
rect 33600 26741 33609 26775
rect 33609 26741 33643 26775
rect 33643 26741 33652 26775
rect 33600 26732 33652 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 7932 26571 7984 26580
rect 7932 26537 7941 26571
rect 7941 26537 7975 26571
rect 7975 26537 7984 26571
rect 7932 26528 7984 26537
rect 15108 26571 15160 26580
rect 3976 26435 4028 26444
rect 3976 26401 3985 26435
rect 3985 26401 4019 26435
rect 4019 26401 4028 26435
rect 3976 26392 4028 26401
rect 4804 26435 4856 26444
rect 4804 26401 4813 26435
rect 4813 26401 4847 26435
rect 4847 26401 4856 26435
rect 14188 26503 14240 26512
rect 14188 26469 14197 26503
rect 14197 26469 14231 26503
rect 14231 26469 14240 26503
rect 14188 26460 14240 26469
rect 15108 26537 15117 26571
rect 15117 26537 15151 26571
rect 15151 26537 15160 26571
rect 15108 26528 15160 26537
rect 15292 26571 15344 26580
rect 15292 26537 15301 26571
rect 15301 26537 15335 26571
rect 15335 26537 15344 26571
rect 15292 26528 15344 26537
rect 20168 26571 20220 26580
rect 20168 26537 20177 26571
rect 20177 26537 20211 26571
rect 20211 26537 20220 26571
rect 20168 26528 20220 26537
rect 20812 26571 20864 26580
rect 20812 26537 20821 26571
rect 20821 26537 20855 26571
rect 20855 26537 20864 26571
rect 20812 26528 20864 26537
rect 22376 26528 22428 26580
rect 30564 26528 30616 26580
rect 19432 26460 19484 26512
rect 4804 26392 4856 26401
rect 10600 26435 10652 26444
rect 10600 26401 10609 26435
rect 10609 26401 10643 26435
rect 10643 26401 10652 26435
rect 10600 26392 10652 26401
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 14004 26392 14056 26444
rect 14924 26435 14976 26444
rect 14924 26401 14933 26435
rect 14933 26401 14967 26435
rect 14967 26401 14976 26435
rect 14924 26392 14976 26401
rect 5632 26324 5684 26376
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 8024 26367 8076 26376
rect 6920 26324 6972 26333
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 8208 26324 8260 26376
rect 12072 26367 12124 26376
rect 12072 26333 12081 26367
rect 12081 26333 12115 26367
rect 12115 26333 12124 26367
rect 12072 26324 12124 26333
rect 7932 26256 7984 26308
rect 15016 26324 15068 26376
rect 17960 26324 18012 26376
rect 20628 26392 20680 26444
rect 20996 26460 21048 26512
rect 29368 26460 29420 26512
rect 38016 26503 38068 26512
rect 38016 26469 38025 26503
rect 38025 26469 38059 26503
rect 38059 26469 38068 26503
rect 38016 26460 38068 26469
rect 22836 26392 22888 26444
rect 23848 26435 23900 26444
rect 23848 26401 23857 26435
rect 23857 26401 23891 26435
rect 23891 26401 23900 26435
rect 23848 26392 23900 26401
rect 26976 26435 27028 26444
rect 26976 26401 26985 26435
rect 26985 26401 27019 26435
rect 27019 26401 27028 26435
rect 26976 26392 27028 26401
rect 30380 26392 30432 26444
rect 24400 26367 24452 26376
rect 24400 26333 24409 26367
rect 24409 26333 24443 26367
rect 24443 26333 24452 26367
rect 24400 26324 24452 26333
rect 30288 26367 30340 26376
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 37832 26367 37884 26376
rect 37832 26333 37841 26367
rect 37841 26333 37875 26367
rect 37875 26333 37884 26367
rect 37832 26324 37884 26333
rect 14832 26299 14884 26308
rect 3056 26188 3108 26240
rect 3976 26188 4028 26240
rect 8300 26231 8352 26240
rect 8300 26197 8309 26231
rect 8309 26197 8343 26231
rect 8343 26197 8352 26231
rect 8300 26188 8352 26197
rect 14832 26265 14841 26299
rect 14841 26265 14875 26299
rect 14875 26265 14884 26299
rect 14832 26256 14884 26265
rect 15660 26256 15712 26308
rect 19432 26256 19484 26308
rect 20628 26256 20680 26308
rect 22192 26299 22244 26308
rect 22192 26265 22201 26299
rect 22201 26265 22235 26299
rect 22235 26265 22244 26299
rect 22192 26256 22244 26265
rect 26240 26256 26292 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 3056 26027 3108 26036
rect 3056 25993 3065 26027
rect 3065 25993 3099 26027
rect 3099 25993 3108 26027
rect 3056 25984 3108 25993
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 3608 25984 3660 26036
rect 4620 25916 4672 25968
rect 6920 25916 6972 25968
rect 10784 25959 10836 25968
rect 10784 25925 10793 25959
rect 10793 25925 10827 25959
rect 10827 25925 10836 25959
rect 10784 25916 10836 25925
rect 18236 25916 18288 25968
rect 26240 25984 26292 26036
rect 28080 25984 28132 26036
rect 29368 26027 29420 26036
rect 29368 25993 29377 26027
rect 29377 25993 29411 26027
rect 29411 25993 29420 26027
rect 29368 25984 29420 25993
rect 30380 26027 30432 26036
rect 30380 25993 30389 26027
rect 30389 25993 30423 26027
rect 30423 25993 30432 26027
rect 30380 25984 30432 25993
rect 23940 25916 23992 25968
rect 26700 25916 26752 25968
rect 26884 25916 26936 25968
rect 3700 25891 3752 25900
rect 3700 25857 3709 25891
rect 3709 25857 3743 25891
rect 3743 25857 3752 25891
rect 3700 25848 3752 25857
rect 4068 25848 4120 25900
rect 7748 25848 7800 25900
rect 7932 25848 7984 25900
rect 8208 25848 8260 25900
rect 12072 25891 12124 25900
rect 12072 25857 12081 25891
rect 12081 25857 12115 25891
rect 12115 25857 12124 25891
rect 12072 25848 12124 25857
rect 14740 25848 14792 25900
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 24400 25848 24452 25900
rect 4804 25780 4856 25832
rect 8024 25823 8076 25832
rect 8024 25789 8033 25823
rect 8033 25789 8067 25823
rect 8067 25789 8076 25823
rect 8024 25780 8076 25789
rect 9128 25823 9180 25832
rect 9128 25789 9137 25823
rect 9137 25789 9171 25823
rect 9171 25789 9180 25823
rect 9128 25780 9180 25789
rect 13268 25780 13320 25832
rect 13452 25823 13504 25832
rect 13452 25789 13461 25823
rect 13461 25789 13495 25823
rect 13495 25789 13504 25823
rect 13452 25780 13504 25789
rect 9588 25712 9640 25764
rect 15016 25712 15068 25764
rect 15568 25755 15620 25764
rect 15568 25721 15577 25755
rect 15577 25721 15611 25755
rect 15611 25721 15620 25755
rect 15568 25712 15620 25721
rect 17684 25780 17736 25832
rect 19432 25823 19484 25832
rect 19432 25789 19441 25823
rect 19441 25789 19475 25823
rect 19475 25789 19484 25823
rect 19432 25780 19484 25789
rect 22560 25780 22612 25832
rect 24308 25780 24360 25832
rect 27160 25848 27212 25900
rect 30564 25916 30616 25968
rect 31300 25916 31352 25968
rect 29368 25848 29420 25900
rect 34336 25891 34388 25900
rect 34336 25857 34345 25891
rect 34345 25857 34379 25891
rect 34379 25857 34388 25891
rect 34336 25848 34388 25857
rect 34428 25891 34480 25900
rect 34428 25857 34437 25891
rect 34437 25857 34471 25891
rect 34471 25857 34480 25891
rect 34428 25848 34480 25857
rect 25412 25823 25464 25832
rect 25412 25789 25421 25823
rect 25421 25789 25455 25823
rect 25455 25789 25464 25823
rect 25412 25780 25464 25789
rect 27068 25823 27120 25832
rect 27068 25789 27077 25823
rect 27077 25789 27111 25823
rect 27111 25789 27120 25823
rect 27068 25780 27120 25789
rect 34704 25848 34756 25900
rect 35900 25848 35952 25900
rect 23388 25712 23440 25764
rect 29092 25712 29144 25764
rect 33600 25712 33652 25764
rect 34612 25712 34664 25764
rect 2872 25644 2924 25696
rect 4712 25644 4764 25696
rect 7840 25687 7892 25696
rect 7840 25653 7849 25687
rect 7849 25653 7883 25687
rect 7883 25653 7892 25687
rect 7840 25644 7892 25653
rect 10048 25644 10100 25696
rect 30104 25644 30156 25696
rect 34152 25687 34204 25696
rect 34152 25653 34161 25687
rect 34161 25653 34195 25687
rect 34195 25653 34204 25687
rect 34152 25644 34204 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1584 25440 1636 25492
rect 4712 25440 4764 25492
rect 9128 25483 9180 25492
rect 9128 25449 9137 25483
rect 9137 25449 9171 25483
rect 9171 25449 9180 25483
rect 9128 25440 9180 25449
rect 9588 25483 9640 25492
rect 9588 25449 9597 25483
rect 9597 25449 9631 25483
rect 9631 25449 9640 25483
rect 9588 25440 9640 25449
rect 14924 25440 14976 25492
rect 15200 25483 15252 25492
rect 15200 25449 15209 25483
rect 15209 25449 15243 25483
rect 15243 25449 15252 25483
rect 15200 25440 15252 25449
rect 17684 25483 17736 25492
rect 17684 25449 17693 25483
rect 17693 25449 17727 25483
rect 17727 25449 17736 25483
rect 17684 25440 17736 25449
rect 22192 25440 22244 25492
rect 22560 25483 22612 25492
rect 22560 25449 22569 25483
rect 22569 25449 22603 25483
rect 22603 25449 22612 25483
rect 22560 25440 22612 25449
rect 23756 25440 23808 25492
rect 24308 25440 24360 25492
rect 30288 25483 30340 25492
rect 30288 25449 30297 25483
rect 30297 25449 30331 25483
rect 30331 25449 30340 25483
rect 30288 25440 30340 25449
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 4804 25304 4856 25356
rect 15292 25347 15344 25356
rect 15292 25313 15301 25347
rect 15301 25313 15335 25347
rect 15335 25313 15344 25347
rect 15292 25304 15344 25313
rect 24492 25347 24544 25356
rect 24492 25313 24501 25347
rect 24501 25313 24535 25347
rect 24535 25313 24544 25347
rect 24492 25304 24544 25313
rect 1952 25279 2004 25288
rect 1952 25245 1961 25279
rect 1961 25245 1995 25279
rect 1995 25245 2004 25279
rect 1952 25236 2004 25245
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 4068 25279 4120 25288
rect 4068 25245 4077 25279
rect 4077 25245 4111 25279
rect 4111 25245 4120 25279
rect 4068 25236 4120 25245
rect 2412 25211 2464 25220
rect 2412 25177 2421 25211
rect 2421 25177 2455 25211
rect 2455 25177 2464 25211
rect 2412 25168 2464 25177
rect 3884 25168 3936 25220
rect 3056 25143 3108 25152
rect 3056 25109 3065 25143
rect 3065 25109 3099 25143
rect 3099 25109 3108 25143
rect 3056 25100 3108 25109
rect 7656 25236 7708 25288
rect 7932 25279 7984 25288
rect 7932 25245 7941 25279
rect 7941 25245 7975 25279
rect 7975 25245 7984 25279
rect 7932 25236 7984 25245
rect 8300 25236 8352 25288
rect 14648 25236 14700 25288
rect 15016 25236 15068 25288
rect 15384 25279 15436 25288
rect 15384 25245 15393 25279
rect 15393 25245 15427 25279
rect 15427 25245 15436 25279
rect 15384 25236 15436 25245
rect 14832 25168 14884 25220
rect 4344 25100 4396 25152
rect 7748 25143 7800 25152
rect 7748 25109 7757 25143
rect 7757 25109 7791 25143
rect 7791 25109 7800 25143
rect 7748 25100 7800 25109
rect 17500 25279 17552 25288
rect 17500 25245 17509 25279
rect 17509 25245 17543 25279
rect 17543 25245 17552 25279
rect 17500 25236 17552 25245
rect 18144 25279 18196 25288
rect 18144 25245 18153 25279
rect 18153 25245 18187 25279
rect 18187 25245 18196 25279
rect 18144 25236 18196 25245
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 22100 25236 22152 25288
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 24032 25236 24084 25288
rect 29920 25279 29972 25288
rect 29920 25245 29929 25279
rect 29929 25245 29963 25279
rect 29963 25245 29972 25279
rect 29920 25236 29972 25245
rect 30104 25279 30156 25288
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 23480 25168 23532 25220
rect 17868 25100 17920 25152
rect 25596 25100 25648 25152
rect 26884 25143 26936 25152
rect 26884 25109 26893 25143
rect 26893 25109 26927 25143
rect 26927 25109 26936 25143
rect 26884 25100 26936 25109
rect 27068 25100 27120 25152
rect 27804 25100 27856 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 8024 24939 8076 24948
rect 8024 24905 8033 24939
rect 8033 24905 8067 24939
rect 8067 24905 8076 24939
rect 8024 24896 8076 24905
rect 29092 24939 29144 24948
rect 29092 24905 29101 24939
rect 29101 24905 29135 24939
rect 29135 24905 29144 24939
rect 29092 24896 29144 24905
rect 14832 24828 14884 24880
rect 17868 24871 17920 24880
rect 17868 24837 17877 24871
rect 17877 24837 17911 24871
rect 17911 24837 17920 24871
rect 17868 24828 17920 24837
rect 23664 24828 23716 24880
rect 24492 24828 24544 24880
rect 1952 24760 2004 24812
rect 4068 24760 4120 24812
rect 4344 24692 4396 24744
rect 5816 24760 5868 24812
rect 7840 24803 7892 24812
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 23020 24760 23072 24812
rect 23480 24760 23532 24812
rect 24032 24803 24084 24812
rect 24032 24769 24041 24803
rect 24041 24769 24075 24803
rect 24075 24769 24084 24803
rect 24032 24760 24084 24769
rect 10784 24692 10836 24744
rect 13912 24692 13964 24744
rect 15292 24735 15344 24744
rect 15292 24701 15301 24735
rect 15301 24701 15335 24735
rect 15335 24701 15344 24735
rect 15292 24692 15344 24701
rect 18236 24735 18288 24744
rect 4804 24624 4856 24676
rect 7840 24624 7892 24676
rect 15384 24624 15436 24676
rect 17500 24624 17552 24676
rect 18236 24701 18245 24735
rect 18245 24701 18279 24735
rect 18279 24701 18288 24735
rect 18236 24692 18288 24701
rect 18144 24624 18196 24676
rect 23480 24624 23532 24676
rect 25412 24624 25464 24676
rect 5816 24599 5868 24608
rect 5816 24565 5825 24599
rect 5825 24565 5859 24599
rect 5859 24565 5868 24599
rect 5816 24556 5868 24565
rect 6276 24556 6328 24608
rect 6920 24556 6972 24608
rect 15200 24599 15252 24608
rect 15200 24565 15209 24599
rect 15209 24565 15243 24599
rect 15243 24565 15252 24599
rect 15200 24556 15252 24565
rect 23756 24599 23808 24608
rect 23756 24565 23765 24599
rect 23765 24565 23799 24599
rect 23799 24565 23808 24599
rect 23756 24556 23808 24565
rect 27804 24556 27856 24608
rect 30196 24760 30248 24812
rect 36084 24760 36136 24812
rect 36268 24803 36320 24812
rect 36268 24769 36277 24803
rect 36277 24769 36311 24803
rect 36311 24769 36320 24803
rect 36268 24760 36320 24769
rect 35900 24624 35952 24676
rect 30932 24556 30984 24608
rect 34796 24599 34848 24608
rect 34796 24565 34805 24599
rect 34805 24565 34839 24599
rect 34839 24565 34848 24599
rect 34796 24556 34848 24565
rect 35716 24599 35768 24608
rect 35716 24565 35725 24599
rect 35725 24565 35759 24599
rect 35759 24565 35768 24599
rect 35716 24556 35768 24565
rect 37372 24556 37424 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2412 24352 2464 24404
rect 15292 24352 15344 24404
rect 15384 24352 15436 24404
rect 22100 24352 22152 24404
rect 30196 24395 30248 24404
rect 30196 24361 30205 24395
rect 30205 24361 30239 24395
rect 30239 24361 30248 24395
rect 30196 24352 30248 24361
rect 14832 24284 14884 24336
rect 30472 24284 30524 24336
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 7196 24148 7248 24200
rect 14096 24148 14148 24200
rect 14648 24191 14700 24200
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 15200 24148 15252 24200
rect 15752 24148 15804 24200
rect 20444 24148 20496 24200
rect 29920 24191 29972 24200
rect 29920 24157 29929 24191
rect 29929 24157 29963 24191
rect 29963 24157 29972 24191
rect 29920 24148 29972 24157
rect 30288 24148 30340 24200
rect 30840 24191 30892 24200
rect 30840 24157 30849 24191
rect 30849 24157 30883 24191
rect 30883 24157 30892 24191
rect 30840 24148 30892 24157
rect 30932 24148 30984 24200
rect 28816 24123 28868 24132
rect 28816 24089 28825 24123
rect 28825 24089 28859 24123
rect 28859 24089 28868 24123
rect 28816 24080 28868 24089
rect 11796 24012 11848 24064
rect 22100 24055 22152 24064
rect 22100 24021 22109 24055
rect 22109 24021 22143 24055
rect 22143 24021 22152 24055
rect 22100 24012 22152 24021
rect 29828 24012 29880 24064
rect 36176 24284 36228 24336
rect 34152 24148 34204 24200
rect 34796 24148 34848 24200
rect 35716 24148 35768 24200
rect 34888 24080 34940 24132
rect 32496 24012 32548 24064
rect 35532 24012 35584 24064
rect 36268 24148 36320 24200
rect 36820 24191 36872 24200
rect 36820 24157 36829 24191
rect 36829 24157 36863 24191
rect 36863 24157 36872 24191
rect 36820 24148 36872 24157
rect 36084 24080 36136 24132
rect 37004 24080 37056 24132
rect 37280 24055 37332 24064
rect 37280 24021 37289 24055
rect 37289 24021 37323 24055
rect 37323 24021 37332 24055
rect 37280 24012 37332 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 13912 23851 13964 23860
rect 13912 23817 13921 23851
rect 13921 23817 13955 23851
rect 13955 23817 13964 23851
rect 13912 23808 13964 23817
rect 29000 23851 29052 23860
rect 29000 23817 29009 23851
rect 29009 23817 29043 23851
rect 29043 23817 29052 23851
rect 29000 23808 29052 23817
rect 30288 23851 30340 23860
rect 30288 23817 30297 23851
rect 30297 23817 30331 23851
rect 30331 23817 30340 23851
rect 30288 23808 30340 23817
rect 37372 23851 37424 23860
rect 37372 23817 37381 23851
rect 37381 23817 37415 23851
rect 37415 23817 37424 23851
rect 37372 23808 37424 23817
rect 7104 23740 7156 23792
rect 11796 23783 11848 23792
rect 11796 23749 11805 23783
rect 11805 23749 11839 23783
rect 11839 23749 11848 23783
rect 11796 23740 11848 23749
rect 13176 23740 13228 23792
rect 14832 23783 14884 23792
rect 14832 23749 14841 23783
rect 14841 23749 14875 23783
rect 14875 23749 14884 23783
rect 14832 23740 14884 23749
rect 18236 23740 18288 23792
rect 26424 23740 26476 23792
rect 29828 23783 29880 23792
rect 29828 23749 29837 23783
rect 29837 23749 29871 23783
rect 29871 23749 29880 23783
rect 29828 23740 29880 23749
rect 30840 23740 30892 23792
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 14188 23672 14240 23724
rect 20444 23715 20496 23724
rect 20444 23681 20453 23715
rect 20453 23681 20487 23715
rect 20487 23681 20496 23715
rect 20444 23672 20496 23681
rect 22100 23672 22152 23724
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 34520 23740 34572 23792
rect 32496 23715 32548 23724
rect 32496 23681 32530 23715
rect 32530 23681 32548 23715
rect 32496 23672 32548 23681
rect 34888 23715 34940 23724
rect 7380 23647 7432 23656
rect 7380 23613 7389 23647
rect 7389 23613 7423 23647
rect 7423 23613 7432 23647
rect 7380 23604 7432 23613
rect 11612 23647 11664 23656
rect 3424 23536 3476 23588
rect 11612 23613 11621 23647
rect 11621 23613 11655 23647
rect 11655 23613 11664 23647
rect 11612 23604 11664 23613
rect 13544 23604 13596 23656
rect 14464 23604 14516 23656
rect 15292 23604 15344 23656
rect 19432 23604 19484 23656
rect 29092 23604 29144 23656
rect 29736 23604 29788 23656
rect 34888 23681 34897 23715
rect 34897 23681 34931 23715
rect 34931 23681 34940 23715
rect 34888 23672 34940 23681
rect 35532 23740 35584 23792
rect 34796 23604 34848 23656
rect 23480 23536 23532 23588
rect 36728 23579 36780 23588
rect 36728 23545 36737 23579
rect 36737 23545 36771 23579
rect 36771 23545 36780 23579
rect 36728 23536 36780 23545
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 13820 23468 13872 23520
rect 16028 23468 16080 23520
rect 16856 23468 16908 23520
rect 22928 23511 22980 23520
rect 22928 23477 22937 23511
rect 22937 23477 22971 23511
rect 22971 23477 22980 23511
rect 22928 23468 22980 23477
rect 26792 23468 26844 23520
rect 33876 23468 33928 23520
rect 35624 23468 35676 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6552 23307 6604 23316
rect 6552 23273 6561 23307
rect 6561 23273 6595 23307
rect 6595 23273 6604 23307
rect 6552 23264 6604 23273
rect 7380 23264 7432 23316
rect 11612 23264 11664 23316
rect 13820 23264 13872 23316
rect 14096 23307 14148 23316
rect 14096 23273 14105 23307
rect 14105 23273 14139 23307
rect 14139 23273 14148 23307
rect 14096 23264 14148 23273
rect 6644 23196 6696 23248
rect 6736 23196 6788 23248
rect 7840 23196 7892 23248
rect 27160 23264 27212 23316
rect 36820 23264 36872 23316
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2780 23060 2832 23112
rect 5356 23060 5408 23112
rect 7748 23128 7800 23180
rect 14464 23171 14516 23180
rect 14464 23137 14473 23171
rect 14473 23137 14507 23171
rect 14507 23137 14516 23171
rect 14464 23128 14516 23137
rect 16856 23171 16908 23180
rect 16856 23137 16865 23171
rect 16865 23137 16899 23171
rect 16899 23137 16908 23171
rect 16856 23128 16908 23137
rect 22928 23128 22980 23180
rect 23940 23128 23992 23180
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 2964 22924 3016 22976
rect 5632 22924 5684 22976
rect 6368 22992 6420 23044
rect 6460 22992 6512 23044
rect 6736 23060 6788 23112
rect 6828 23060 6880 23112
rect 12900 23103 12952 23112
rect 7656 22992 7708 23044
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 12900 23060 12952 23069
rect 12992 23103 13044 23112
rect 12992 23069 13001 23103
rect 13001 23069 13035 23103
rect 13035 23069 13044 23103
rect 13176 23103 13228 23112
rect 12992 23060 13044 23069
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 14188 23060 14240 23112
rect 14832 23060 14884 23112
rect 15660 23060 15712 23112
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 26792 23103 26844 23112
rect 26792 23069 26810 23103
rect 26810 23069 26844 23103
rect 27068 23103 27120 23112
rect 26792 23060 26844 23069
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 27528 23060 27580 23112
rect 27896 23103 27948 23112
rect 27896 23069 27905 23103
rect 27905 23069 27939 23103
rect 27939 23069 27948 23103
rect 27896 23060 27948 23069
rect 34520 23060 34572 23112
rect 35624 23060 35676 23112
rect 7840 22924 7892 22976
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 19340 22992 19392 23044
rect 22744 22992 22796 23044
rect 25688 22967 25740 22976
rect 25688 22933 25697 22967
rect 25697 22933 25731 22967
rect 25731 22933 25740 22967
rect 25688 22924 25740 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 5356 22763 5408 22772
rect 5356 22729 5365 22763
rect 5365 22729 5399 22763
rect 5399 22729 5408 22763
rect 5356 22720 5408 22729
rect 6828 22763 6880 22772
rect 2964 22695 3016 22704
rect 2964 22661 2973 22695
rect 2973 22661 3007 22695
rect 3007 22661 3016 22695
rect 2964 22652 3016 22661
rect 3608 22652 3660 22704
rect 6368 22695 6420 22704
rect 6368 22661 6377 22695
rect 6377 22661 6411 22695
rect 6411 22661 6420 22695
rect 6368 22652 6420 22661
rect 6828 22729 6837 22763
rect 6837 22729 6871 22763
rect 6871 22729 6880 22763
rect 6828 22720 6880 22729
rect 7840 22695 7892 22704
rect 7840 22661 7849 22695
rect 7849 22661 7883 22695
rect 7883 22661 7892 22695
rect 7840 22652 7892 22661
rect 12900 22720 12952 22772
rect 14188 22720 14240 22772
rect 27528 22763 27580 22772
rect 27528 22729 27537 22763
rect 27537 22729 27571 22763
rect 27571 22729 27580 22763
rect 27528 22720 27580 22729
rect 27896 22720 27948 22772
rect 32036 22720 32088 22772
rect 35900 22720 35952 22772
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 6460 22584 6512 22636
rect 7656 22627 7708 22636
rect 7656 22593 7665 22627
rect 7665 22593 7699 22627
rect 7699 22593 7708 22627
rect 7656 22584 7708 22593
rect 23848 22652 23900 22704
rect 25688 22652 25740 22704
rect 34704 22652 34756 22704
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 6736 22516 6788 22568
rect 11704 22559 11756 22568
rect 11704 22525 11713 22559
rect 11713 22525 11747 22559
rect 11747 22525 11756 22559
rect 11704 22516 11756 22525
rect 13268 22559 13320 22568
rect 13268 22525 13277 22559
rect 13277 22525 13311 22559
rect 13311 22525 13320 22559
rect 13268 22516 13320 22525
rect 18144 22559 18196 22568
rect 18144 22525 18153 22559
rect 18153 22525 18187 22559
rect 18187 22525 18196 22559
rect 18144 22516 18196 22525
rect 18328 22559 18380 22568
rect 18328 22525 18337 22559
rect 18337 22525 18371 22559
rect 18371 22525 18380 22559
rect 18328 22516 18380 22525
rect 24492 22559 24544 22568
rect 19340 22448 19392 22500
rect 24492 22525 24501 22559
rect 24501 22525 24535 22559
rect 24535 22525 24544 22559
rect 24492 22516 24544 22525
rect 26884 22584 26936 22636
rect 29460 22584 29512 22636
rect 30012 22584 30064 22636
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 37188 22584 37240 22636
rect 28172 22516 28224 22568
rect 26332 22491 26384 22500
rect 26332 22457 26341 22491
rect 26341 22457 26375 22491
rect 26375 22457 26384 22491
rect 26332 22448 26384 22457
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 6552 22380 6604 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6552 22176 6604 22228
rect 13820 22176 13872 22228
rect 18144 22176 18196 22228
rect 36176 22108 36228 22160
rect 6644 22040 6696 22092
rect 12992 22083 13044 22092
rect 12992 22049 13001 22083
rect 13001 22049 13035 22083
rect 13035 22049 13044 22083
rect 12992 22040 13044 22049
rect 20996 22040 21048 22092
rect 22744 22083 22796 22092
rect 22744 22049 22753 22083
rect 22753 22049 22787 22083
rect 22787 22049 22796 22083
rect 22744 22040 22796 22049
rect 25688 22083 25740 22092
rect 25688 22049 25697 22083
rect 25697 22049 25731 22083
rect 25731 22049 25740 22083
rect 25688 22040 25740 22049
rect 26424 22083 26476 22092
rect 26424 22049 26433 22083
rect 26433 22049 26467 22083
rect 26467 22049 26476 22083
rect 26424 22040 26476 22049
rect 29460 22040 29512 22092
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 7288 22015 7340 22024
rect 6460 21972 6512 21981
rect 6920 21904 6972 21956
rect 7012 21836 7064 21888
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 10324 21972 10376 22024
rect 12900 22015 12952 22024
rect 10508 21836 10560 21888
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 13176 22015 13228 22024
rect 13176 21981 13185 22015
rect 13185 21981 13219 22015
rect 13219 21981 13228 22015
rect 13176 21972 13228 21981
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 22468 22015 22520 22024
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22468 21972 22520 21981
rect 27712 22015 27764 22024
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 30380 21972 30432 22024
rect 36360 21972 36412 22024
rect 36820 21972 36872 22024
rect 19984 21904 20036 21956
rect 26240 21947 26292 21956
rect 26240 21913 26249 21947
rect 26249 21913 26283 21947
rect 26283 21913 26292 21947
rect 26240 21904 26292 21913
rect 19432 21879 19484 21888
rect 19432 21845 19441 21879
rect 19441 21845 19475 21879
rect 19475 21845 19484 21879
rect 19432 21836 19484 21845
rect 25688 21836 25740 21888
rect 29000 21904 29052 21956
rect 30104 21947 30156 21956
rect 30104 21913 30113 21947
rect 30113 21913 30147 21947
rect 30147 21913 30156 21947
rect 30104 21904 30156 21913
rect 36268 21904 36320 21956
rect 36728 21904 36780 21956
rect 27528 21879 27580 21888
rect 27528 21845 27537 21879
rect 27537 21845 27571 21879
rect 27571 21845 27580 21879
rect 27528 21836 27580 21845
rect 32036 21879 32088 21888
rect 32036 21845 32045 21879
rect 32045 21845 32079 21879
rect 32079 21845 32088 21879
rect 32036 21836 32088 21845
rect 35716 21879 35768 21888
rect 35716 21845 35725 21879
rect 35725 21845 35759 21879
rect 35759 21845 35768 21879
rect 35716 21836 35768 21845
rect 37372 21879 37424 21888
rect 37372 21845 37381 21879
rect 37381 21845 37415 21879
rect 37415 21845 37424 21879
rect 37372 21836 37424 21845
rect 38016 21879 38068 21888
rect 38016 21845 38025 21879
rect 38025 21845 38059 21879
rect 38059 21845 38068 21879
rect 38016 21836 38068 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11704 21632 11756 21684
rect 13176 21632 13228 21684
rect 13360 21632 13412 21684
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 27712 21632 27764 21684
rect 36360 21632 36412 21684
rect 6920 21564 6972 21616
rect 7380 21564 7432 21616
rect 27528 21564 27580 21616
rect 36176 21564 36228 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 6460 21496 6512 21548
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 7012 21496 7064 21548
rect 12716 21496 12768 21548
rect 14004 21496 14056 21548
rect 15200 21496 15252 21548
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 14188 21428 14240 21480
rect 21548 21496 21600 21548
rect 24492 21496 24544 21548
rect 27068 21496 27120 21548
rect 28540 21496 28592 21548
rect 29920 21496 29972 21548
rect 33876 21496 33928 21548
rect 36268 21496 36320 21548
rect 21364 21428 21416 21480
rect 30012 21471 30064 21480
rect 30012 21437 30021 21471
rect 30021 21437 30055 21471
rect 30055 21437 30064 21471
rect 30012 21428 30064 21437
rect 30288 21471 30340 21480
rect 30288 21437 30297 21471
rect 30297 21437 30331 21471
rect 30331 21437 30340 21471
rect 30288 21428 30340 21437
rect 5172 21360 5224 21412
rect 5448 21360 5500 21412
rect 20996 21403 21048 21412
rect 20996 21369 21005 21403
rect 21005 21369 21039 21403
rect 21039 21369 21048 21403
rect 20996 21360 21048 21369
rect 2780 21292 2832 21344
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 6368 21335 6420 21344
rect 6368 21301 6377 21335
rect 6377 21301 6411 21335
rect 6411 21301 6420 21335
rect 6368 21292 6420 21301
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 6736 21292 6788 21344
rect 28264 21292 28316 21344
rect 32588 21335 32640 21344
rect 32588 21301 32597 21335
rect 32597 21301 32631 21335
rect 32631 21301 32640 21335
rect 32588 21292 32640 21301
rect 35624 21292 35676 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1584 21088 1636 21140
rect 2504 21131 2556 21140
rect 2504 21097 2513 21131
rect 2513 21097 2547 21131
rect 2547 21097 2556 21131
rect 2504 21088 2556 21097
rect 14188 21131 14240 21140
rect 14188 21097 14197 21131
rect 14197 21097 14231 21131
rect 14231 21097 14240 21131
rect 14188 21088 14240 21097
rect 21364 21131 21416 21140
rect 3424 21020 3476 21072
rect 2780 20952 2832 21004
rect 5816 20952 5868 21004
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 2596 20927 2648 20936
rect 2596 20893 2605 20927
rect 2605 20893 2639 20927
rect 2639 20893 2648 20927
rect 2596 20884 2648 20893
rect 6368 20884 6420 20936
rect 20904 21020 20956 21072
rect 21364 21097 21373 21131
rect 21373 21097 21407 21131
rect 21407 21097 21416 21131
rect 21364 21088 21416 21097
rect 28540 21131 28592 21140
rect 28540 21097 28549 21131
rect 28549 21097 28583 21131
rect 28583 21097 28592 21131
rect 28540 21088 28592 21097
rect 31484 21088 31536 21140
rect 25504 21020 25556 21072
rect 32128 21088 32180 21140
rect 32312 21020 32364 21072
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 10508 20995 10560 21004
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 14648 20952 14700 21004
rect 15200 20952 15252 21004
rect 16580 20995 16632 21004
rect 16580 20961 16589 20995
rect 16589 20961 16623 20995
rect 16623 20961 16632 20995
rect 16580 20952 16632 20961
rect 18328 20952 18380 21004
rect 14556 20884 14608 20936
rect 16488 20884 16540 20936
rect 18420 20927 18472 20936
rect 18420 20893 18429 20927
rect 18429 20893 18463 20927
rect 18463 20893 18472 20927
rect 18420 20884 18472 20893
rect 19432 20884 19484 20936
rect 19984 20952 20036 21004
rect 26240 20952 26292 21004
rect 27068 20952 27120 21004
rect 20076 20884 20128 20936
rect 20720 20884 20772 20936
rect 21824 20927 21876 20936
rect 12164 20859 12216 20868
rect 12164 20825 12173 20859
rect 12173 20825 12207 20859
rect 12207 20825 12216 20859
rect 12164 20816 12216 20825
rect 20444 20816 20496 20868
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 24400 20927 24452 20936
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 25780 20816 25832 20868
rect 28172 20859 28224 20868
rect 28172 20825 28181 20859
rect 28181 20825 28215 20859
rect 28215 20825 28224 20859
rect 28172 20816 28224 20825
rect 28264 20859 28316 20868
rect 28264 20825 28273 20859
rect 28273 20825 28307 20859
rect 28307 20825 28316 20859
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 32036 20884 32088 20936
rect 34520 20884 34572 20936
rect 28264 20816 28316 20825
rect 30104 20816 30156 20868
rect 31024 20816 31076 20868
rect 1400 20791 1452 20800
rect 1400 20757 1409 20791
rect 1409 20757 1443 20791
rect 1443 20757 1452 20791
rect 1400 20748 1452 20757
rect 2872 20791 2924 20800
rect 2872 20757 2881 20791
rect 2881 20757 2915 20791
rect 2915 20757 2924 20791
rect 2872 20748 2924 20757
rect 4896 20748 4948 20800
rect 23296 20748 23348 20800
rect 27436 20791 27488 20800
rect 27436 20757 27445 20791
rect 27445 20757 27479 20791
rect 27479 20757 27488 20791
rect 27436 20748 27488 20757
rect 29368 20748 29420 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2504 20544 2556 20596
rect 17224 20544 17276 20596
rect 19432 20587 19484 20596
rect 19432 20553 19441 20587
rect 19441 20553 19475 20587
rect 19475 20553 19484 20587
rect 19432 20544 19484 20553
rect 21824 20544 21876 20596
rect 31024 20587 31076 20596
rect 31024 20553 31033 20587
rect 31033 20553 31067 20587
rect 31067 20553 31076 20587
rect 31024 20544 31076 20553
rect 16580 20476 16632 20528
rect 23296 20476 23348 20528
rect 30104 20476 30156 20528
rect 36084 20476 36136 20528
rect 1400 20451 1452 20460
rect 1400 20417 1409 20451
rect 1409 20417 1443 20451
rect 1443 20417 1452 20451
rect 1400 20408 1452 20417
rect 1584 20408 1636 20460
rect 2596 20408 2648 20460
rect 2780 20451 2832 20460
rect 2780 20417 2789 20451
rect 2789 20417 2823 20451
rect 2823 20417 2832 20451
rect 2780 20408 2832 20417
rect 1860 20272 1912 20324
rect 7932 20408 7984 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 18696 20408 18748 20460
rect 20444 20408 20496 20460
rect 20720 20408 20772 20460
rect 28264 20408 28316 20460
rect 30380 20451 30432 20460
rect 30380 20417 30389 20451
rect 30389 20417 30423 20451
rect 30423 20417 30432 20451
rect 30380 20408 30432 20417
rect 12992 20340 13044 20392
rect 15844 20383 15896 20392
rect 15844 20349 15853 20383
rect 15853 20349 15887 20383
rect 15887 20349 15896 20383
rect 15844 20340 15896 20349
rect 16488 20340 16540 20392
rect 19432 20340 19484 20392
rect 20076 20340 20128 20392
rect 27436 20340 27488 20392
rect 30288 20340 30340 20392
rect 34704 20451 34756 20460
rect 34704 20417 34713 20451
rect 34713 20417 34747 20451
rect 34747 20417 34756 20451
rect 34704 20408 34756 20417
rect 35440 20451 35492 20460
rect 35440 20417 35449 20451
rect 35449 20417 35483 20451
rect 35483 20417 35492 20451
rect 35440 20408 35492 20417
rect 35716 20340 35768 20392
rect 36360 20340 36412 20392
rect 18512 20272 18564 20324
rect 21916 20315 21968 20324
rect 21916 20281 21925 20315
rect 21925 20281 21959 20315
rect 21959 20281 21968 20315
rect 21916 20272 21968 20281
rect 2504 20247 2556 20256
rect 2504 20213 2513 20247
rect 2513 20213 2547 20247
rect 2547 20213 2556 20247
rect 2504 20204 2556 20213
rect 3240 20204 3292 20256
rect 3792 20204 3844 20256
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 7380 20204 7432 20256
rect 12072 20204 12124 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 18788 20204 18840 20213
rect 20904 20204 20956 20256
rect 35900 20204 35952 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2964 20000 3016 20052
rect 13820 20000 13872 20052
rect 3056 19932 3108 19984
rect 10324 19932 10376 19984
rect 12440 19932 12492 19984
rect 14740 19932 14792 19984
rect 16672 20000 16724 20052
rect 18420 20000 18472 20052
rect 20904 20043 20956 20052
rect 20904 20009 20913 20043
rect 20913 20009 20947 20043
rect 20947 20009 20956 20043
rect 20904 20000 20956 20009
rect 37648 20043 37700 20052
rect 4712 19907 4764 19916
rect 4712 19873 4721 19907
rect 4721 19873 4755 19907
rect 4755 19873 4764 19907
rect 4712 19864 4764 19873
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 4988 19864 5040 19916
rect 11888 19864 11940 19916
rect 12072 19907 12124 19916
rect 12072 19873 12081 19907
rect 12081 19873 12115 19907
rect 12115 19873 12124 19907
rect 12072 19864 12124 19873
rect 12992 19864 13044 19916
rect 15844 19864 15896 19916
rect 18696 19932 18748 19984
rect 16120 19864 16172 19916
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 3240 19839 3292 19848
rect 3240 19805 3249 19839
rect 3249 19805 3283 19839
rect 3283 19805 3292 19839
rect 3792 19839 3844 19848
rect 3240 19796 3292 19805
rect 3792 19805 3801 19839
rect 3801 19805 3835 19839
rect 3835 19805 3844 19839
rect 3792 19796 3844 19805
rect 2596 19728 2648 19780
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13820 19796 13872 19848
rect 3976 19728 4028 19780
rect 10968 19728 11020 19780
rect 11796 19728 11848 19780
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 4068 19660 4120 19712
rect 4620 19660 4672 19712
rect 11612 19660 11664 19712
rect 16948 19796 17000 19848
rect 18788 19796 18840 19848
rect 20720 19932 20772 19984
rect 20168 19864 20220 19916
rect 32588 19932 32640 19984
rect 25228 19864 25280 19916
rect 28816 19864 28868 19916
rect 30288 19907 30340 19916
rect 30288 19873 30297 19907
rect 30297 19873 30331 19907
rect 30331 19873 30340 19907
rect 30288 19864 30340 19873
rect 20536 19796 20588 19848
rect 21916 19796 21968 19848
rect 35624 19932 35676 19984
rect 16580 19728 16632 19780
rect 18420 19728 18472 19780
rect 18512 19660 18564 19712
rect 25412 19728 25464 19780
rect 26332 19728 26384 19780
rect 27252 19771 27304 19780
rect 27252 19737 27261 19771
rect 27261 19737 27295 19771
rect 27295 19737 27304 19771
rect 27252 19728 27304 19737
rect 22100 19660 22152 19712
rect 29736 19728 29788 19780
rect 35716 19796 35768 19848
rect 36084 19796 36136 19848
rect 36360 19839 36412 19848
rect 36360 19805 36369 19839
rect 36369 19805 36403 19839
rect 36403 19805 36412 19839
rect 36360 19796 36412 19805
rect 37648 20009 37657 20043
rect 37657 20009 37691 20043
rect 37691 20009 37700 20043
rect 37648 20000 37700 20009
rect 37648 19796 37700 19848
rect 32036 19728 32088 19780
rect 35348 19728 35400 19780
rect 30564 19660 30616 19712
rect 31300 19703 31352 19712
rect 31300 19669 31309 19703
rect 31309 19669 31343 19703
rect 31343 19669 31352 19703
rect 31300 19660 31352 19669
rect 34704 19660 34756 19712
rect 35716 19660 35768 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4988 19456 5040 19508
rect 11796 19499 11848 19508
rect 11796 19465 11805 19499
rect 11805 19465 11839 19499
rect 11839 19465 11848 19499
rect 11796 19456 11848 19465
rect 11888 19456 11940 19508
rect 2872 19388 2924 19440
rect 3608 19388 3660 19440
rect 3976 19388 4028 19440
rect 4068 19388 4120 19440
rect 6736 19388 6788 19440
rect 7932 19388 7984 19440
rect 10324 19431 10376 19440
rect 10324 19397 10333 19431
rect 10333 19397 10367 19431
rect 10367 19397 10376 19431
rect 10324 19388 10376 19397
rect 12992 19388 13044 19440
rect 13360 19431 13412 19440
rect 1952 19320 2004 19372
rect 4160 19320 4212 19372
rect 11612 19363 11664 19372
rect 11612 19329 11621 19363
rect 11621 19329 11655 19363
rect 11655 19329 11664 19363
rect 11612 19320 11664 19329
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 13360 19397 13369 19431
rect 13369 19397 13403 19431
rect 13403 19397 13412 19431
rect 13360 19388 13412 19397
rect 14004 19431 14056 19440
rect 14004 19397 14013 19431
rect 14013 19397 14047 19431
rect 14047 19397 14056 19431
rect 14004 19388 14056 19397
rect 14648 19388 14700 19440
rect 13912 19320 13964 19372
rect 16580 19388 16632 19440
rect 18696 19456 18748 19508
rect 18972 19456 19024 19508
rect 24400 19456 24452 19508
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 16488 19320 16540 19372
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 20260 19388 20312 19440
rect 22928 19388 22980 19440
rect 27252 19456 27304 19508
rect 29736 19499 29788 19508
rect 29736 19465 29745 19499
rect 29745 19465 29779 19499
rect 29779 19465 29788 19499
rect 29736 19456 29788 19465
rect 30380 19499 30432 19508
rect 30380 19465 30389 19499
rect 30389 19465 30423 19499
rect 30423 19465 30432 19499
rect 30380 19456 30432 19465
rect 26976 19388 27028 19440
rect 29092 19388 29144 19440
rect 30104 19388 30156 19440
rect 32128 19456 32180 19508
rect 35348 19499 35400 19508
rect 35348 19465 35357 19499
rect 35357 19465 35391 19499
rect 35391 19465 35400 19499
rect 35348 19456 35400 19465
rect 35532 19456 35584 19508
rect 36084 19456 36136 19508
rect 36452 19388 36504 19440
rect 16948 19320 17000 19329
rect 20076 19320 20128 19372
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 22284 19320 22336 19372
rect 3056 19252 3108 19304
rect 14372 19252 14424 19304
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 23020 19295 23072 19304
rect 23020 19261 23029 19295
rect 23029 19261 23063 19295
rect 23063 19261 23072 19295
rect 23020 19252 23072 19261
rect 23296 19320 23348 19372
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 24400 19320 24452 19372
rect 29368 19363 29420 19372
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 30012 19320 30064 19372
rect 31300 19320 31352 19372
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 29828 19252 29880 19304
rect 30196 19252 30248 19304
rect 30012 19184 30064 19236
rect 34704 19363 34756 19372
rect 34704 19329 34713 19363
rect 34713 19329 34747 19363
rect 34747 19329 34756 19363
rect 34704 19320 34756 19329
rect 35716 19320 35768 19372
rect 35440 19252 35492 19304
rect 2964 19116 3016 19168
rect 4712 19116 4764 19168
rect 4896 19116 4948 19168
rect 6460 19159 6512 19168
rect 6460 19125 6469 19159
rect 6469 19125 6503 19159
rect 6503 19125 6512 19159
rect 6460 19116 6512 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 13820 19116 13872 19168
rect 14004 19116 14056 19168
rect 14832 19116 14884 19168
rect 16580 19116 16632 19168
rect 17132 19159 17184 19168
rect 17132 19125 17141 19159
rect 17141 19125 17175 19159
rect 17175 19125 17184 19159
rect 17132 19116 17184 19125
rect 18144 19116 18196 19168
rect 22376 19159 22428 19168
rect 22376 19125 22385 19159
rect 22385 19125 22419 19159
rect 22419 19125 22428 19159
rect 22376 19116 22428 19125
rect 22836 19159 22888 19168
rect 22836 19125 22845 19159
rect 22845 19125 22879 19159
rect 22879 19125 22888 19159
rect 22836 19116 22888 19125
rect 28632 19116 28684 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 4160 18819 4212 18828
rect 4160 18785 4169 18819
rect 4169 18785 4203 18819
rect 4203 18785 4212 18819
rect 4160 18776 4212 18785
rect 4712 18776 4764 18828
rect 5632 18844 5684 18896
rect 9036 18912 9088 18964
rect 21916 18912 21968 18964
rect 22100 18955 22152 18964
rect 22100 18921 22109 18955
rect 22109 18921 22143 18955
rect 22143 18921 22152 18955
rect 22100 18912 22152 18921
rect 22836 18912 22888 18964
rect 24308 18912 24360 18964
rect 32128 18912 32180 18964
rect 35440 18955 35492 18964
rect 35440 18921 35449 18955
rect 35449 18921 35483 18955
rect 35483 18921 35492 18955
rect 35440 18912 35492 18921
rect 37648 18912 37700 18964
rect 14648 18776 14700 18828
rect 26332 18844 26384 18896
rect 22100 18776 22152 18828
rect 23020 18819 23072 18828
rect 23020 18785 23029 18819
rect 23029 18785 23063 18819
rect 23063 18785 23072 18819
rect 23020 18776 23072 18785
rect 26976 18819 27028 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 4620 18708 4672 18760
rect 5172 18708 5224 18760
rect 7104 18708 7156 18760
rect 15200 18708 15252 18760
rect 15844 18708 15896 18760
rect 20168 18708 20220 18760
rect 21916 18708 21968 18760
rect 6460 18640 6512 18692
rect 9772 18640 9824 18692
rect 11980 18640 12032 18692
rect 12256 18640 12308 18692
rect 16580 18683 16632 18692
rect 16580 18649 16589 18683
rect 16589 18649 16623 18683
rect 16623 18649 16632 18683
rect 16580 18640 16632 18649
rect 22376 18708 22428 18760
rect 23112 18708 23164 18760
rect 7472 18615 7524 18624
rect 7472 18581 7481 18615
rect 7481 18581 7515 18615
rect 7515 18581 7524 18615
rect 7472 18572 7524 18581
rect 14372 18572 14424 18624
rect 20076 18615 20128 18624
rect 20076 18581 20085 18615
rect 20085 18581 20119 18615
rect 20119 18581 20128 18615
rect 20076 18572 20128 18581
rect 22836 18640 22888 18692
rect 23296 18640 23348 18692
rect 26976 18785 26985 18819
rect 26985 18785 27019 18819
rect 27019 18785 27028 18819
rect 26976 18776 27028 18785
rect 30564 18776 30616 18828
rect 28908 18708 28960 18760
rect 31576 18708 31628 18760
rect 32036 18751 32088 18760
rect 32036 18717 32045 18751
rect 32045 18717 32079 18751
rect 32079 18717 32088 18751
rect 32036 18708 32088 18717
rect 35624 18708 35676 18760
rect 36452 18708 36504 18760
rect 31300 18640 31352 18692
rect 31668 18640 31720 18692
rect 22284 18572 22336 18624
rect 24768 18572 24820 18624
rect 30012 18572 30064 18624
rect 32312 18572 32364 18624
rect 33600 18572 33652 18624
rect 35808 18572 35860 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 5632 18368 5684 18420
rect 7288 18368 7340 18420
rect 11980 18411 12032 18420
rect 11980 18377 11989 18411
rect 11989 18377 12023 18411
rect 12023 18377 12032 18411
rect 11980 18368 12032 18377
rect 6828 18232 6880 18284
rect 9772 18300 9824 18352
rect 18788 18368 18840 18420
rect 22100 18411 22152 18420
rect 22100 18377 22109 18411
rect 22109 18377 22143 18411
rect 22143 18377 22152 18411
rect 22100 18368 22152 18377
rect 24400 18368 24452 18420
rect 26332 18411 26384 18420
rect 26332 18377 26341 18411
rect 26341 18377 26375 18411
rect 26375 18377 26384 18411
rect 26332 18368 26384 18377
rect 27436 18411 27488 18420
rect 27436 18377 27445 18411
rect 27445 18377 27479 18411
rect 27479 18377 27488 18411
rect 27436 18368 27488 18377
rect 27712 18368 27764 18420
rect 29092 18368 29144 18420
rect 33600 18411 33652 18420
rect 33600 18377 33609 18411
rect 33609 18377 33643 18411
rect 33643 18377 33652 18411
rect 33600 18368 33652 18377
rect 35900 18368 35952 18420
rect 37832 18368 37884 18420
rect 8392 18275 8444 18284
rect 8392 18241 8401 18275
rect 8401 18241 8435 18275
rect 8435 18241 8444 18275
rect 8392 18232 8444 18241
rect 12900 18232 12952 18284
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 18512 18300 18564 18352
rect 19156 18300 19208 18352
rect 19984 18300 20036 18352
rect 22836 18343 22888 18352
rect 14832 18232 14884 18284
rect 15016 18232 15068 18284
rect 22008 18232 22060 18284
rect 3516 18164 3568 18216
rect 9680 18164 9732 18216
rect 11888 18164 11940 18216
rect 12256 18164 12308 18216
rect 13912 18207 13964 18216
rect 13912 18173 13921 18207
rect 13921 18173 13955 18207
rect 13955 18173 13964 18207
rect 13912 18164 13964 18173
rect 15200 18164 15252 18216
rect 9128 18096 9180 18148
rect 22836 18309 22845 18343
rect 22845 18309 22879 18343
rect 22879 18309 22888 18343
rect 22836 18300 22888 18309
rect 23020 18275 23072 18284
rect 23020 18241 23029 18275
rect 23029 18241 23063 18275
rect 23063 18241 23072 18275
rect 23020 18232 23072 18241
rect 23112 18275 23164 18284
rect 23112 18241 23121 18275
rect 23121 18241 23155 18275
rect 23155 18241 23164 18275
rect 24768 18275 24820 18284
rect 23112 18232 23164 18241
rect 24768 18241 24777 18275
rect 24777 18241 24811 18275
rect 24811 18241 24820 18275
rect 24768 18232 24820 18241
rect 26516 18164 26568 18216
rect 27804 18232 27856 18284
rect 34520 18300 34572 18352
rect 35624 18300 35676 18352
rect 32312 18232 32364 18284
rect 34704 18232 34756 18284
rect 35348 18232 35400 18284
rect 35716 18232 35768 18284
rect 36544 18275 36596 18284
rect 36544 18241 36553 18275
rect 36553 18241 36587 18275
rect 36587 18241 36596 18275
rect 36544 18232 36596 18241
rect 37280 18232 37332 18284
rect 27528 18164 27580 18216
rect 35808 18164 35860 18216
rect 29368 18096 29420 18148
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 5356 18028 5408 18080
rect 6552 18071 6604 18080
rect 6552 18037 6561 18071
rect 6561 18037 6595 18071
rect 6595 18037 6604 18071
rect 6552 18028 6604 18037
rect 7932 18071 7984 18080
rect 7932 18037 7941 18071
rect 7941 18037 7975 18071
rect 7975 18037 7984 18071
rect 7932 18028 7984 18037
rect 8944 18028 8996 18080
rect 13360 18028 13412 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 14648 18071 14700 18080
rect 14648 18037 14657 18071
rect 14657 18037 14691 18071
rect 14691 18037 14700 18071
rect 22928 18071 22980 18080
rect 14648 18028 14700 18037
rect 22928 18037 22937 18071
rect 22937 18037 22971 18071
rect 22971 18037 22980 18071
rect 22928 18028 22980 18037
rect 27804 18071 27856 18080
rect 27804 18037 27813 18071
rect 27813 18037 27847 18071
rect 27847 18037 27856 18071
rect 27804 18028 27856 18037
rect 35348 18071 35400 18080
rect 35348 18037 35357 18071
rect 35357 18037 35391 18071
rect 35391 18037 35400 18071
rect 35348 18028 35400 18037
rect 37280 18071 37332 18080
rect 37280 18037 37289 18071
rect 37289 18037 37323 18071
rect 37323 18037 37332 18071
rect 37280 18028 37332 18037
rect 38016 18071 38068 18080
rect 38016 18037 38025 18071
rect 38025 18037 38059 18071
rect 38059 18037 38068 18071
rect 38016 18028 38068 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 8392 17824 8444 17876
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 22008 17824 22060 17876
rect 22928 17867 22980 17876
rect 22928 17833 22937 17867
rect 22937 17833 22971 17867
rect 22971 17833 22980 17867
rect 22928 17824 22980 17833
rect 29276 17824 29328 17876
rect 2596 17756 2648 17808
rect 18420 17756 18472 17808
rect 18788 17756 18840 17808
rect 6552 17688 6604 17740
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 9680 17731 9732 17740
rect 9680 17697 9689 17731
rect 9689 17697 9723 17731
rect 9723 17697 9732 17731
rect 9680 17688 9732 17697
rect 15200 17688 15252 17740
rect 23020 17756 23072 17808
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 30104 17731 30156 17740
rect 30104 17697 30113 17731
rect 30113 17697 30147 17731
rect 30147 17697 30156 17731
rect 30104 17688 30156 17697
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 7932 17620 7984 17672
rect 12348 17663 12400 17672
rect 12348 17629 12357 17663
rect 12357 17629 12391 17663
rect 12391 17629 12400 17663
rect 12348 17620 12400 17629
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 14832 17620 14884 17672
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 7380 17552 7432 17604
rect 14004 17552 14056 17604
rect 15016 17552 15068 17604
rect 22836 17620 22888 17672
rect 23112 17620 23164 17672
rect 6828 17484 6880 17536
rect 10140 17484 10192 17536
rect 12532 17484 12584 17536
rect 15568 17484 15620 17536
rect 20168 17552 20220 17604
rect 27804 17620 27856 17672
rect 28816 17663 28868 17672
rect 28816 17629 28825 17663
rect 28825 17629 28859 17663
rect 28859 17629 28868 17663
rect 28816 17620 28868 17629
rect 29276 17620 29328 17672
rect 27528 17552 27580 17604
rect 30288 17595 30340 17604
rect 30288 17561 30297 17595
rect 30297 17561 30331 17595
rect 30331 17561 30340 17595
rect 30288 17552 30340 17561
rect 31668 17552 31720 17604
rect 34520 17552 34572 17604
rect 20720 17484 20772 17536
rect 23756 17484 23808 17536
rect 27620 17484 27672 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 6644 17280 6696 17332
rect 4896 17212 4948 17264
rect 7380 17280 7432 17332
rect 7748 17280 7800 17332
rect 9036 17280 9088 17332
rect 10140 17280 10192 17332
rect 17592 17280 17644 17332
rect 22836 17280 22888 17332
rect 36544 17280 36596 17332
rect 12532 17255 12584 17264
rect 12532 17221 12541 17255
rect 12541 17221 12575 17255
rect 12575 17221 12584 17255
rect 12532 17212 12584 17221
rect 7564 17144 7616 17196
rect 7748 17187 7800 17196
rect 7748 17153 7757 17187
rect 7757 17153 7791 17187
rect 7791 17153 7800 17187
rect 7748 17144 7800 17153
rect 7932 17144 7984 17196
rect 12348 17187 12400 17196
rect 12348 17153 12357 17187
rect 12357 17153 12391 17187
rect 12391 17153 12400 17187
rect 12348 17144 12400 17153
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 29000 17212 29052 17264
rect 27252 17187 27304 17196
rect 27252 17153 27286 17187
rect 27286 17153 27304 17187
rect 27252 17144 27304 17153
rect 27528 17144 27580 17196
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 2964 17119 3016 17128
rect 2964 17085 2973 17119
rect 2973 17085 3007 17119
rect 3007 17085 3016 17119
rect 2964 17076 3016 17085
rect 6552 17076 6604 17128
rect 14004 17119 14056 17128
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 17960 17119 18012 17128
rect 17960 17085 17969 17119
rect 17969 17085 18003 17119
rect 18003 17085 18012 17119
rect 17960 17076 18012 17085
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 26148 17076 26200 17128
rect 7472 17008 7524 17060
rect 34704 17144 34756 17196
rect 29368 17076 29420 17128
rect 34796 17076 34848 17128
rect 35532 17076 35584 17128
rect 7656 16940 7708 16992
rect 35348 17008 35400 17060
rect 8576 16940 8628 16992
rect 19340 16940 19392 16992
rect 20168 16940 20220 16992
rect 35900 16940 35952 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2780 16736 2832 16788
rect 7472 16736 7524 16788
rect 9036 16779 9088 16788
rect 9036 16745 9045 16779
rect 9045 16745 9079 16779
rect 9079 16745 9088 16779
rect 9036 16736 9088 16745
rect 17776 16736 17828 16788
rect 27252 16736 27304 16788
rect 3424 16668 3476 16720
rect 8300 16668 8352 16720
rect 6552 16600 6604 16652
rect 13912 16600 13964 16652
rect 23756 16600 23808 16652
rect 30288 16600 30340 16652
rect 35624 16643 35676 16652
rect 35624 16609 35633 16643
rect 35633 16609 35667 16643
rect 35667 16609 35676 16643
rect 35624 16600 35676 16609
rect 3792 16575 3844 16584
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 6644 16575 6696 16584
rect 6644 16541 6653 16575
rect 6653 16541 6687 16575
rect 6687 16541 6696 16575
rect 6644 16532 6696 16541
rect 7564 16575 7616 16584
rect 7564 16541 7573 16575
rect 7573 16541 7607 16575
rect 7607 16541 7616 16575
rect 7564 16532 7616 16541
rect 7932 16532 7984 16584
rect 14464 16532 14516 16584
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 27620 16532 27672 16584
rect 35900 16575 35952 16584
rect 35900 16541 35934 16575
rect 35934 16541 35952 16575
rect 35900 16532 35952 16541
rect 7104 16439 7156 16448
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 14096 16396 14148 16448
rect 15660 16396 15712 16448
rect 20168 16439 20220 16448
rect 20168 16405 20177 16439
rect 20177 16405 20211 16439
rect 20211 16405 20220 16439
rect 20168 16396 20220 16405
rect 35808 16396 35860 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2964 16192 3016 16244
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 17960 16192 18012 16244
rect 19248 16192 19300 16244
rect 23572 16192 23624 16244
rect 23756 16235 23808 16244
rect 23756 16201 23765 16235
rect 23765 16201 23799 16235
rect 23799 16201 23808 16235
rect 23756 16192 23808 16201
rect 31208 16192 31260 16244
rect 31576 16192 31628 16244
rect 3884 16124 3936 16176
rect 14096 16167 14148 16176
rect 14096 16133 14105 16167
rect 14105 16133 14139 16167
rect 14139 16133 14148 16167
rect 14096 16124 14148 16133
rect 18604 16124 18656 16176
rect 23296 16167 23348 16176
rect 3608 16056 3660 16108
rect 4620 16056 4672 16108
rect 13912 16099 13964 16108
rect 4804 15988 4856 16040
rect 7196 15988 7248 16040
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 18236 16056 18288 16108
rect 19064 16056 19116 16108
rect 23296 16133 23305 16167
rect 23305 16133 23339 16167
rect 23339 16133 23348 16167
rect 23296 16124 23348 16133
rect 26148 16167 26200 16176
rect 26148 16133 26157 16167
rect 26157 16133 26191 16167
rect 26191 16133 26200 16167
rect 26148 16124 26200 16133
rect 20996 16056 21048 16108
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 32864 16099 32916 16108
rect 2872 15920 2924 15972
rect 3424 15920 3476 15972
rect 13820 15988 13872 16040
rect 15936 15988 15988 16040
rect 18512 15988 18564 16040
rect 22560 15988 22612 16040
rect 32864 16065 32873 16099
rect 32873 16065 32907 16099
rect 32907 16065 32916 16099
rect 32864 16056 32916 16065
rect 35808 16124 35860 16176
rect 24676 16031 24728 16040
rect 24676 15997 24685 16031
rect 24685 15997 24719 16031
rect 24719 15997 24728 16031
rect 24676 15988 24728 15997
rect 29368 15988 29420 16040
rect 34520 16031 34572 16040
rect 21272 15920 21324 15972
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 4068 15852 4120 15904
rect 4712 15852 4764 15904
rect 4896 15895 4948 15904
rect 4896 15861 4905 15895
rect 4905 15861 4939 15895
rect 4939 15861 4948 15895
rect 4896 15852 4948 15861
rect 11704 15852 11756 15904
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 18696 15895 18748 15904
rect 18696 15861 18705 15895
rect 18705 15861 18739 15895
rect 18739 15861 18748 15895
rect 18696 15852 18748 15861
rect 18880 15852 18932 15904
rect 21732 15852 21784 15904
rect 23296 15895 23348 15904
rect 23296 15861 23305 15895
rect 23305 15861 23339 15895
rect 23339 15861 23348 15895
rect 23296 15852 23348 15861
rect 30012 15852 30064 15904
rect 31116 15852 31168 15904
rect 32128 15895 32180 15904
rect 32128 15861 32137 15895
rect 32137 15861 32171 15895
rect 32171 15861 32180 15895
rect 32128 15852 32180 15861
rect 34520 15997 34529 16031
rect 34529 15997 34563 16031
rect 34563 15997 34572 16031
rect 34520 15988 34572 15997
rect 34612 15852 34664 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 7840 15691 7892 15700
rect 7840 15657 7849 15691
rect 7849 15657 7883 15691
rect 7883 15657 7892 15691
rect 7840 15648 7892 15657
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 18696 15691 18748 15700
rect 18696 15657 18705 15691
rect 18705 15657 18739 15691
rect 18739 15657 18748 15691
rect 18696 15648 18748 15657
rect 29000 15691 29052 15700
rect 3792 15555 3844 15564
rect 3792 15521 3801 15555
rect 3801 15521 3835 15555
rect 3835 15521 3844 15555
rect 3792 15512 3844 15521
rect 3976 15512 4028 15564
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 12900 15512 12952 15564
rect 13544 15555 13596 15564
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 15660 15555 15712 15564
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 16672 15512 16724 15521
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 8576 15444 8628 15496
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 19064 15512 19116 15564
rect 19156 15512 19208 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 21364 15512 21416 15564
rect 29000 15657 29009 15691
rect 29009 15657 29043 15691
rect 29043 15657 29052 15691
rect 29000 15648 29052 15657
rect 32128 15648 32180 15700
rect 23572 15555 23624 15564
rect 23572 15521 23581 15555
rect 23581 15521 23615 15555
rect 23615 15521 23624 15555
rect 23572 15512 23624 15521
rect 18512 15487 18564 15496
rect 18512 15453 18521 15487
rect 18521 15453 18555 15487
rect 18555 15453 18564 15487
rect 18512 15444 18564 15453
rect 20168 15444 20220 15496
rect 20812 15487 20864 15496
rect 18696 15419 18748 15428
rect 18696 15385 18705 15419
rect 18705 15385 18739 15419
rect 18739 15385 18748 15419
rect 18696 15376 18748 15385
rect 18880 15376 18932 15428
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 22376 15487 22428 15496
rect 22376 15453 22385 15487
rect 22385 15453 22419 15487
rect 22419 15453 22428 15487
rect 22376 15444 22428 15453
rect 23296 15444 23348 15496
rect 23664 15487 23716 15496
rect 23664 15453 23673 15487
rect 23673 15453 23707 15487
rect 23707 15453 23716 15487
rect 23664 15444 23716 15453
rect 23480 15376 23532 15428
rect 34796 15648 34848 15700
rect 37372 15648 37424 15700
rect 24676 15555 24728 15564
rect 24676 15521 24685 15555
rect 24685 15521 24719 15555
rect 24719 15521 24728 15555
rect 24676 15512 24728 15521
rect 29092 15512 29144 15564
rect 29368 15512 29420 15564
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 34612 15512 34664 15564
rect 35532 15512 35584 15564
rect 28908 15444 28960 15496
rect 31116 15487 31168 15496
rect 31116 15453 31125 15487
rect 31125 15453 31159 15487
rect 31159 15453 31168 15487
rect 31116 15444 31168 15453
rect 31208 15487 31260 15496
rect 31208 15453 31217 15487
rect 31217 15453 31251 15487
rect 31251 15453 31260 15487
rect 31208 15444 31260 15453
rect 34060 15444 34112 15496
rect 34704 15487 34756 15496
rect 34704 15453 34713 15487
rect 34713 15453 34747 15487
rect 34747 15453 34756 15487
rect 34704 15444 34756 15453
rect 8668 15308 8720 15360
rect 17132 15308 17184 15360
rect 25504 15376 25556 15428
rect 30288 15376 30340 15428
rect 36452 15376 36504 15428
rect 23848 15351 23900 15360
rect 23848 15317 23857 15351
rect 23857 15317 23891 15351
rect 23891 15317 23900 15351
rect 23848 15308 23900 15317
rect 29644 15351 29696 15360
rect 29644 15317 29653 15351
rect 29653 15317 29687 15351
rect 29687 15317 29696 15351
rect 29644 15308 29696 15317
rect 30012 15351 30064 15360
rect 30012 15317 30021 15351
rect 30021 15317 30055 15351
rect 30055 15317 30064 15351
rect 30012 15308 30064 15317
rect 32220 15308 32272 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 18972 15104 19024 15156
rect 20812 15104 20864 15156
rect 32864 15104 32916 15156
rect 34612 15147 34664 15156
rect 34612 15113 34621 15147
rect 34621 15113 34655 15147
rect 34655 15113 34664 15147
rect 34612 15104 34664 15113
rect 36452 15104 36504 15156
rect 4712 15079 4764 15088
rect 4712 15045 4721 15079
rect 4721 15045 4755 15079
rect 4755 15045 4764 15079
rect 4712 15036 4764 15045
rect 8668 15079 8720 15088
rect 8668 15045 8677 15079
rect 8677 15045 8711 15079
rect 8711 15045 8720 15079
rect 8668 15036 8720 15045
rect 13268 15036 13320 15088
rect 21640 15036 21692 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 4896 15011 4948 15020
rect 4896 14977 4905 15011
rect 4905 14977 4939 15011
rect 4939 14977 4948 15011
rect 4896 14968 4948 14977
rect 7104 14968 7156 15020
rect 11244 14968 11296 15020
rect 13452 14968 13504 15020
rect 14188 14968 14240 15020
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 17684 14968 17736 15020
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 8944 14900 8996 14952
rect 11704 14943 11756 14952
rect 3424 14832 3476 14884
rect 10232 14832 10284 14884
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 14096 14943 14148 14952
rect 14096 14909 14105 14943
rect 14105 14909 14139 14943
rect 14139 14909 14148 14943
rect 14096 14900 14148 14909
rect 18512 14900 18564 14952
rect 18788 14943 18840 14952
rect 18788 14909 18797 14943
rect 18797 14909 18831 14943
rect 18831 14909 18840 14943
rect 18788 14900 18840 14909
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 16672 14832 16724 14884
rect 19524 14832 19576 14884
rect 21364 14968 21416 15020
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 23572 15036 23624 15088
rect 29000 15036 29052 15088
rect 29736 15036 29788 15088
rect 30288 15036 30340 15088
rect 28816 14968 28868 15020
rect 30472 15011 30524 15020
rect 30472 14977 30490 15011
rect 30490 14977 30524 15011
rect 30472 14968 30524 14977
rect 21180 14900 21232 14952
rect 22008 14900 22060 14952
rect 21640 14832 21692 14884
rect 28632 14832 28684 14884
rect 28908 14832 28960 14884
rect 29368 14875 29420 14884
rect 29368 14841 29377 14875
rect 29377 14841 29411 14875
rect 29411 14841 29420 14875
rect 29368 14832 29420 14841
rect 2780 14764 2832 14816
rect 7748 14764 7800 14816
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 14280 14807 14332 14816
rect 14280 14773 14289 14807
rect 14289 14773 14323 14807
rect 14323 14773 14332 14807
rect 14280 14764 14332 14773
rect 17960 14807 18012 14816
rect 17960 14773 17969 14807
rect 17969 14773 18003 14807
rect 18003 14773 18012 14807
rect 17960 14764 18012 14773
rect 21916 14764 21968 14816
rect 22376 14807 22428 14816
rect 22376 14773 22385 14807
rect 22385 14773 22419 14807
rect 22419 14773 22428 14807
rect 22376 14764 22428 14773
rect 23388 14807 23440 14816
rect 23388 14773 23397 14807
rect 23397 14773 23431 14807
rect 23431 14773 23440 14807
rect 23388 14764 23440 14773
rect 30104 14764 30156 14816
rect 32220 14968 32272 15020
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2504 14603 2556 14612
rect 2504 14569 2513 14603
rect 2513 14569 2547 14603
rect 2547 14569 2556 14603
rect 2504 14560 2556 14569
rect 3056 14560 3108 14612
rect 4068 14560 4120 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 12348 14560 12400 14612
rect 12440 14560 12492 14612
rect 21916 14603 21968 14612
rect 21916 14569 21925 14603
rect 21925 14569 21959 14603
rect 21959 14569 21968 14603
rect 21916 14560 21968 14569
rect 22468 14560 22520 14612
rect 22560 14560 22612 14612
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 4160 14424 4212 14476
rect 4804 14424 4856 14476
rect 11704 14424 11756 14476
rect 14280 14424 14332 14476
rect 16764 14492 16816 14544
rect 19156 14492 19208 14544
rect 19064 14424 19116 14476
rect 1584 14356 1636 14408
rect 2780 14399 2832 14408
rect 2780 14365 2789 14399
rect 2789 14365 2823 14399
rect 2823 14365 2832 14399
rect 2780 14356 2832 14365
rect 3608 14356 3660 14408
rect 4712 14356 4764 14408
rect 8024 14399 8076 14408
rect 8024 14365 8033 14399
rect 8033 14365 8067 14399
rect 8067 14365 8076 14399
rect 8024 14356 8076 14365
rect 13268 14356 13320 14408
rect 17960 14356 18012 14408
rect 18880 14356 18932 14408
rect 18972 14356 19024 14408
rect 19524 14399 19576 14408
rect 19524 14365 19533 14399
rect 19533 14365 19567 14399
rect 19567 14365 19576 14399
rect 19524 14356 19576 14365
rect 21364 14424 21416 14476
rect 21732 14399 21784 14408
rect 3884 14288 3936 14340
rect 2964 14263 3016 14272
rect 2964 14229 2973 14263
rect 2973 14229 3007 14263
rect 3007 14229 3016 14263
rect 2964 14220 3016 14229
rect 3424 14220 3476 14272
rect 9588 14288 9640 14340
rect 14188 14288 14240 14340
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 17684 14220 17736 14272
rect 18696 14288 18748 14340
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 22100 14424 22152 14476
rect 23388 14424 23440 14476
rect 25504 14424 25556 14476
rect 25596 14424 25648 14476
rect 23664 14356 23716 14408
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 27528 14356 27580 14408
rect 28816 14560 28868 14612
rect 30472 14560 30524 14612
rect 34704 14560 34756 14612
rect 29368 14356 29420 14408
rect 29644 14356 29696 14408
rect 34520 14356 34572 14408
rect 35532 14356 35584 14408
rect 38016 14331 38068 14340
rect 38016 14297 38025 14331
rect 38025 14297 38059 14331
rect 38059 14297 38068 14331
rect 38016 14288 38068 14297
rect 21364 14220 21416 14272
rect 28080 14263 28132 14272
rect 28080 14229 28089 14263
rect 28089 14229 28123 14263
rect 28123 14229 28132 14263
rect 28080 14220 28132 14229
rect 37924 14263 37976 14272
rect 37924 14229 37933 14263
rect 37933 14229 37967 14263
rect 37967 14229 37976 14263
rect 37924 14220 37976 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4620 14016 4672 14068
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 13268 14059 13320 14068
rect 13268 14025 13277 14059
rect 13277 14025 13311 14059
rect 13311 14025 13320 14059
rect 13268 14016 13320 14025
rect 3884 13991 3936 14000
rect 3884 13957 3893 13991
rect 3893 13957 3927 13991
rect 3927 13957 3936 13991
rect 3884 13948 3936 13957
rect 7932 13991 7984 14000
rect 7932 13957 7941 13991
rect 7941 13957 7975 13991
rect 7975 13957 7984 13991
rect 7932 13948 7984 13957
rect 14188 13948 14240 14000
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 4160 13812 4212 13864
rect 4620 13880 4672 13932
rect 7748 13923 7800 13932
rect 7748 13889 7757 13923
rect 7757 13889 7791 13923
rect 7791 13889 7800 13923
rect 7748 13880 7800 13889
rect 12348 13923 12400 13932
rect 12348 13889 12357 13923
rect 12357 13889 12391 13923
rect 12391 13889 12400 13923
rect 12348 13880 12400 13889
rect 13452 13923 13504 13932
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 22008 14016 22060 14068
rect 32588 14059 32640 14068
rect 32588 14025 32597 14059
rect 32597 14025 32631 14059
rect 32631 14025 32640 14059
rect 32588 14016 32640 14025
rect 34796 14016 34848 14068
rect 15200 13948 15252 14000
rect 13452 13880 13504 13889
rect 18788 13880 18840 13932
rect 4804 13812 4856 13864
rect 5080 13812 5132 13864
rect 8300 13855 8352 13864
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 14096 13812 14148 13864
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 21364 13948 21416 14000
rect 34060 13991 34112 14000
rect 34060 13957 34069 13991
rect 34069 13957 34103 13991
rect 34103 13957 34112 13991
rect 34060 13948 34112 13957
rect 20720 13880 20772 13932
rect 23848 13880 23900 13932
rect 29920 13880 29972 13932
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 25964 13812 26016 13864
rect 29368 13812 29420 13864
rect 30104 13812 30156 13864
rect 35440 13812 35492 13864
rect 35532 13855 35584 13864
rect 35532 13821 35541 13855
rect 35541 13821 35575 13855
rect 35575 13821 35584 13855
rect 35532 13812 35584 13821
rect 4068 13676 4120 13728
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 13820 13676 13872 13728
rect 14280 13676 14332 13728
rect 20352 13719 20404 13728
rect 20352 13685 20361 13719
rect 20361 13685 20395 13719
rect 20395 13685 20404 13719
rect 20352 13676 20404 13685
rect 20812 13719 20864 13728
rect 20812 13685 20821 13719
rect 20821 13685 20855 13719
rect 20855 13685 20864 13719
rect 20812 13676 20864 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2504 13472 2556 13524
rect 4712 13472 4764 13524
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 20812 13472 20864 13524
rect 21916 13515 21968 13524
rect 21916 13481 21925 13515
rect 21925 13481 21959 13515
rect 21959 13481 21968 13515
rect 21916 13472 21968 13481
rect 4068 13404 4120 13456
rect 24400 13472 24452 13524
rect 29920 13472 29972 13524
rect 30104 13515 30156 13524
rect 30104 13481 30113 13515
rect 30113 13481 30147 13515
rect 30147 13481 30156 13515
rect 30104 13472 30156 13481
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 5540 13336 5592 13388
rect 17408 13336 17460 13388
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 19432 13336 19484 13388
rect 20352 13336 20404 13388
rect 20628 13336 20680 13388
rect 26884 13379 26936 13388
rect 26884 13345 26893 13379
rect 26893 13345 26927 13379
rect 26927 13345 26936 13379
rect 26884 13336 26936 13345
rect 27528 13336 27580 13388
rect 1400 13268 1452 13277
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 6552 13268 6604 13320
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 17224 13268 17276 13320
rect 19984 13268 20036 13320
rect 20720 13268 20772 13320
rect 21732 13311 21784 13320
rect 17500 13200 17552 13252
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 33416 13268 33468 13320
rect 34704 13268 34756 13320
rect 21364 13200 21416 13252
rect 28080 13200 28132 13252
rect 34428 13200 34480 13252
rect 22192 13132 22244 13184
rect 35256 13132 35308 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7840 12928 7892 12980
rect 9588 12903 9640 12912
rect 9588 12869 9597 12903
rect 9597 12869 9631 12903
rect 9631 12869 9640 12903
rect 9588 12860 9640 12869
rect 13176 12860 13228 12912
rect 21732 12928 21784 12980
rect 19064 12860 19116 12912
rect 19984 12860 20036 12912
rect 22008 12860 22060 12912
rect 29092 12928 29144 12980
rect 29736 12971 29788 12980
rect 29736 12937 29745 12971
rect 29745 12937 29779 12971
rect 29779 12937 29788 12971
rect 29736 12928 29788 12937
rect 34796 12928 34848 12980
rect 27712 12860 27764 12912
rect 28816 12860 28868 12912
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 12440 12792 12492 12844
rect 13452 12792 13504 12844
rect 22560 12792 22612 12844
rect 25872 12792 25924 12844
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 9680 12656 9732 12708
rect 11704 12588 11756 12640
rect 11796 12588 11848 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 13084 12631 13136 12640
rect 13084 12597 13093 12631
rect 13093 12597 13127 12631
rect 13127 12597 13136 12631
rect 13084 12588 13136 12597
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 35256 12835 35308 12844
rect 35256 12801 35265 12835
rect 35265 12801 35299 12835
rect 35299 12801 35308 12835
rect 35256 12792 35308 12801
rect 29276 12767 29328 12776
rect 29276 12733 29285 12767
rect 29285 12733 29319 12767
rect 29319 12733 29328 12767
rect 29276 12724 29328 12733
rect 33508 12724 33560 12776
rect 34428 12724 34480 12776
rect 35440 12835 35492 12844
rect 35440 12801 35449 12835
rect 35449 12801 35483 12835
rect 35483 12801 35492 12835
rect 35440 12792 35492 12801
rect 13820 12588 13872 12640
rect 21916 12631 21968 12640
rect 21916 12597 21925 12631
rect 21925 12597 21959 12631
rect 21959 12597 21968 12631
rect 21916 12588 21968 12597
rect 22284 12588 22336 12640
rect 22468 12588 22520 12640
rect 23756 12588 23808 12640
rect 24308 12631 24360 12640
rect 24308 12597 24317 12631
rect 24317 12597 24351 12631
rect 24351 12597 24360 12631
rect 24308 12588 24360 12597
rect 26884 12588 26936 12640
rect 30472 12588 30524 12640
rect 36084 12588 36136 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3608 12384 3660 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 6460 12384 6512 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 17408 12384 17460 12436
rect 17500 12384 17552 12436
rect 9680 12316 9732 12368
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 4712 12248 4764 12300
rect 12164 12316 12216 12368
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 1400 12180 1452 12189
rect 2596 12044 2648 12096
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 4620 12180 4672 12232
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 9128 12180 9180 12232
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17592 12248 17644 12300
rect 20444 12384 20496 12436
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 22468 12427 22520 12436
rect 22468 12393 22477 12427
rect 22477 12393 22511 12427
rect 22511 12393 22520 12427
rect 22468 12384 22520 12393
rect 32588 12427 32640 12436
rect 32588 12393 32597 12427
rect 32597 12393 32631 12427
rect 32631 12393 32640 12427
rect 32588 12384 32640 12393
rect 35440 12384 35492 12436
rect 35808 12384 35860 12436
rect 22100 12248 22152 12300
rect 25964 12291 26016 12300
rect 25964 12257 25973 12291
rect 25973 12257 26007 12291
rect 26007 12257 26016 12291
rect 25964 12248 26016 12257
rect 27252 12291 27304 12300
rect 27252 12257 27261 12291
rect 27261 12257 27295 12291
rect 27295 12257 27304 12291
rect 27252 12248 27304 12257
rect 29736 12248 29788 12300
rect 12440 12180 12492 12189
rect 11520 12155 11572 12164
rect 11520 12121 11529 12155
rect 11529 12121 11563 12155
rect 11563 12121 11572 12155
rect 11520 12112 11572 12121
rect 17224 12223 17276 12232
rect 4160 12044 4212 12096
rect 8208 12044 8260 12096
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 21640 12180 21692 12232
rect 22560 12180 22612 12232
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 12256 12087 12308 12096
rect 12256 12053 12265 12087
rect 12265 12053 12299 12087
rect 12299 12053 12308 12087
rect 12256 12044 12308 12053
rect 18880 12112 18932 12164
rect 25044 12155 25096 12164
rect 25044 12121 25053 12155
rect 25053 12121 25087 12155
rect 25087 12121 25096 12155
rect 25044 12112 25096 12121
rect 32588 12180 32640 12232
rect 33140 12180 33192 12232
rect 27436 12112 27488 12164
rect 29920 12112 29972 12164
rect 33416 12223 33468 12232
rect 33416 12189 33425 12223
rect 33425 12189 33459 12223
rect 33459 12189 33468 12223
rect 33416 12180 33468 12189
rect 33508 12112 33560 12164
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 18512 12044 18564 12096
rect 23112 12044 23164 12096
rect 32404 12044 32456 12096
rect 33692 12087 33744 12096
rect 33692 12053 33701 12087
rect 33701 12053 33735 12087
rect 33735 12053 33744 12087
rect 33692 12044 33744 12053
rect 35348 12044 35400 12096
rect 36084 12180 36136 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 7656 11840 7708 11892
rect 17868 11840 17920 11892
rect 28908 11840 28960 11892
rect 29736 11840 29788 11892
rect 4160 11815 4212 11824
rect 4160 11781 4169 11815
rect 4169 11781 4203 11815
rect 4203 11781 4212 11815
rect 4160 11772 4212 11781
rect 10968 11815 11020 11824
rect 6460 11704 6512 11756
rect 4620 11636 4672 11688
rect 10968 11781 10977 11815
rect 10977 11781 11011 11815
rect 11011 11781 11020 11815
rect 10968 11772 11020 11781
rect 13176 11815 13228 11824
rect 13176 11781 13185 11815
rect 13185 11781 13219 11815
rect 13219 11781 13228 11815
rect 13176 11772 13228 11781
rect 13544 11772 13596 11824
rect 7380 11704 7432 11756
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 11520 11704 11572 11756
rect 13084 11704 13136 11756
rect 17224 11772 17276 11824
rect 17500 11772 17552 11824
rect 10600 11636 10652 11688
rect 12532 11636 12584 11688
rect 13360 11636 13412 11688
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 23756 11704 23808 11756
rect 29920 11815 29972 11824
rect 29920 11781 29929 11815
rect 29929 11781 29963 11815
rect 29963 11781 29972 11815
rect 29920 11772 29972 11781
rect 30472 11772 30524 11824
rect 33140 11772 33192 11824
rect 29184 11704 29236 11756
rect 29552 11704 29604 11756
rect 27344 11636 27396 11688
rect 28816 11636 28868 11688
rect 13268 11500 13320 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 14096 11500 14148 11552
rect 16212 11500 16264 11552
rect 29644 11568 29696 11620
rect 30288 11704 30340 11756
rect 30104 11636 30156 11688
rect 33416 11840 33468 11892
rect 34428 11840 34480 11892
rect 33692 11772 33744 11824
rect 33508 11636 33560 11688
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 20168 11500 20220 11552
rect 20812 11500 20864 11552
rect 28356 11500 28408 11552
rect 28816 11543 28868 11552
rect 28816 11509 28825 11543
rect 28825 11509 28859 11543
rect 28859 11509 28868 11543
rect 28816 11500 28868 11509
rect 32680 11543 32732 11552
rect 32680 11509 32689 11543
rect 32689 11509 32723 11543
rect 32723 11509 32732 11543
rect 32680 11500 32732 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3976 11339 4028 11348
rect 3976 11305 3985 11339
rect 3985 11305 4019 11339
rect 4019 11305 4028 11339
rect 3976 11296 4028 11305
rect 4896 11296 4948 11348
rect 5540 11296 5592 11348
rect 5724 11296 5776 11348
rect 8208 11296 8260 11348
rect 10600 11339 10652 11348
rect 10600 11305 10609 11339
rect 10609 11305 10643 11339
rect 10643 11305 10652 11339
rect 10600 11296 10652 11305
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 19340 11339 19392 11348
rect 19340 11305 19349 11339
rect 19349 11305 19383 11339
rect 19383 11305 19392 11339
rect 19340 11296 19392 11305
rect 20628 11339 20680 11348
rect 20628 11305 20637 11339
rect 20637 11305 20671 11339
rect 20671 11305 20680 11339
rect 20628 11296 20680 11305
rect 21456 11296 21508 11348
rect 29552 11339 29604 11348
rect 29552 11305 29561 11339
rect 29561 11305 29595 11339
rect 29595 11305 29604 11339
rect 29552 11296 29604 11305
rect 30472 11339 30524 11348
rect 30472 11305 30481 11339
rect 30481 11305 30515 11339
rect 30515 11305 30524 11339
rect 30472 11296 30524 11305
rect 34428 11296 34480 11348
rect 3424 11228 3476 11280
rect 8760 11228 8812 11280
rect 9772 11228 9824 11280
rect 19984 11228 20036 11280
rect 27436 11228 27488 11280
rect 4160 11160 4212 11212
rect 12256 11203 12308 11212
rect 12256 11169 12265 11203
rect 12265 11169 12299 11203
rect 12299 11169 12308 11203
rect 12256 11160 12308 11169
rect 13360 11203 13412 11212
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 16672 11203 16724 11212
rect 16672 11169 16681 11203
rect 16681 11169 16715 11203
rect 16715 11169 16724 11203
rect 16672 11160 16724 11169
rect 18880 11160 18932 11212
rect 20536 11160 20588 11212
rect 22192 11203 22244 11212
rect 22192 11169 22201 11203
rect 22201 11169 22235 11203
rect 22235 11169 22244 11203
rect 22192 11160 22244 11169
rect 29276 11160 29328 11212
rect 32404 11160 32456 11212
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4712 11092 4764 11144
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5448 11092 5500 11144
rect 5908 11092 5960 11144
rect 6828 11092 6880 11144
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 8208 11092 8260 11144
rect 11796 11092 11848 11144
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 24676 11092 24728 11144
rect 25320 11092 25372 11144
rect 30288 11092 30340 11144
rect 34888 11135 34940 11144
rect 34888 11101 34897 11135
rect 34897 11101 34931 11135
rect 34931 11101 34940 11135
rect 34888 11092 34940 11101
rect 5172 11024 5224 11076
rect 26976 11024 27028 11076
rect 29276 11024 29328 11076
rect 34152 11024 34204 11076
rect 35900 11135 35952 11144
rect 35900 11101 35910 11135
rect 35910 11101 35944 11135
rect 35944 11101 35952 11135
rect 35900 11092 35952 11101
rect 35808 11024 35860 11076
rect 8208 10999 8260 11008
rect 8208 10965 8217 10999
rect 8217 10965 8251 10999
rect 8251 10965 8260 10999
rect 8208 10956 8260 10965
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 13084 10956 13136 10965
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 18328 10999 18380 11008
rect 18328 10965 18337 10999
rect 18337 10965 18371 10999
rect 18371 10965 18380 10999
rect 18328 10956 18380 10965
rect 20812 10956 20864 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4160 10752 4212 10804
rect 6460 10752 6512 10804
rect 6828 10752 6880 10804
rect 8116 10752 8168 10804
rect 3240 10684 3292 10736
rect 22100 10752 22152 10804
rect 24584 10752 24636 10804
rect 26976 10795 27028 10804
rect 26976 10761 26985 10795
rect 26985 10761 27019 10795
rect 27019 10761 27028 10795
rect 26976 10752 27028 10761
rect 27436 10752 27488 10804
rect 29736 10752 29788 10804
rect 30288 10752 30340 10804
rect 33232 10752 33284 10804
rect 18328 10684 18380 10736
rect 19064 10727 19116 10736
rect 19064 10693 19073 10727
rect 19073 10693 19107 10727
rect 19107 10693 19116 10727
rect 19064 10684 19116 10693
rect 20260 10684 20312 10736
rect 24676 10727 24728 10736
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3332 10616 3384 10668
rect 4620 10616 4672 10668
rect 5080 10616 5132 10668
rect 6736 10616 6788 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 19340 10616 19392 10668
rect 19984 10616 20036 10668
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 3056 10548 3108 10600
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 20628 10548 20680 10600
rect 20996 10616 21048 10668
rect 24676 10693 24685 10727
rect 24685 10693 24719 10727
rect 24719 10693 24728 10727
rect 24676 10684 24728 10693
rect 25044 10684 25096 10736
rect 29092 10684 29144 10736
rect 29644 10727 29696 10736
rect 29644 10693 29653 10727
rect 29653 10693 29687 10727
rect 29687 10693 29696 10727
rect 29644 10684 29696 10693
rect 34888 10752 34940 10804
rect 27160 10659 27212 10668
rect 6276 10480 6328 10532
rect 21916 10548 21968 10600
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 29368 10616 29420 10668
rect 35900 10684 35952 10736
rect 35808 10616 35860 10668
rect 24584 10548 24636 10600
rect 30196 10548 30248 10600
rect 34796 10548 34848 10600
rect 35716 10548 35768 10600
rect 26424 10480 26476 10532
rect 2412 10412 2464 10464
rect 2964 10412 3016 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 12440 10412 12492 10464
rect 14096 10412 14148 10464
rect 20720 10412 20772 10464
rect 27988 10412 28040 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 5264 10208 5316 10260
rect 6828 10208 6880 10260
rect 17224 10208 17276 10260
rect 20536 10208 20588 10260
rect 27436 10208 27488 10260
rect 29460 10208 29512 10260
rect 29736 10208 29788 10260
rect 4804 10140 4856 10192
rect 6736 10140 6788 10192
rect 14372 10140 14424 10192
rect 18604 10140 18656 10192
rect 5632 10072 5684 10124
rect 5908 10072 5960 10124
rect 14096 10115 14148 10124
rect 2228 10004 2280 10056
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 5172 10004 5224 10056
rect 5540 10004 5592 10056
rect 6276 10004 6328 10056
rect 7472 10004 7524 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 11888 10004 11940 10056
rect 3148 9936 3200 9988
rect 4252 9936 4304 9988
rect 8852 9936 8904 9988
rect 11980 9936 12032 9988
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 14096 10072 14148 10081
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 19340 10004 19392 10056
rect 20720 10140 20772 10192
rect 21548 10140 21600 10192
rect 21916 10140 21968 10192
rect 29644 10140 29696 10192
rect 20628 10072 20680 10124
rect 27344 10115 27396 10124
rect 27344 10081 27353 10115
rect 27353 10081 27387 10115
rect 27387 10081 27396 10115
rect 27344 10072 27396 10081
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23112 10004 23164 10013
rect 27528 10047 27580 10056
rect 27528 10013 27537 10047
rect 27537 10013 27571 10047
rect 27571 10013 27580 10047
rect 27528 10004 27580 10013
rect 29460 10004 29512 10056
rect 29644 10047 29696 10056
rect 29644 10013 29653 10047
rect 29653 10013 29687 10047
rect 29687 10013 29696 10047
rect 29644 10004 29696 10013
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 30288 10072 30340 10124
rect 38108 10047 38160 10056
rect 25688 9979 25740 9988
rect 16580 9868 16632 9920
rect 18512 9868 18564 9920
rect 25688 9945 25697 9979
rect 25697 9945 25731 9979
rect 25731 9945 25740 9979
rect 25688 9936 25740 9945
rect 27988 9936 28040 9988
rect 29276 9936 29328 9988
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 30748 9936 30800 9988
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 22836 9868 22888 9920
rect 22928 9911 22980 9920
rect 22928 9877 22937 9911
rect 22937 9877 22971 9911
rect 22971 9877 22980 9911
rect 22928 9868 22980 9877
rect 30656 9868 30708 9920
rect 32128 9911 32180 9920
rect 32128 9877 32137 9911
rect 32137 9877 32171 9911
rect 32171 9877 32180 9911
rect 32128 9868 32180 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3424 9664 3476 9716
rect 10784 9664 10836 9716
rect 16580 9664 16632 9716
rect 2964 9596 3016 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3240 9528 3292 9580
rect 4252 9596 4304 9648
rect 4896 9596 4948 9648
rect 5632 9596 5684 9648
rect 7288 9596 7340 9648
rect 7472 9639 7524 9648
rect 7472 9605 7481 9639
rect 7481 9605 7515 9639
rect 7515 9605 7524 9639
rect 7472 9596 7524 9605
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 14004 9596 14056 9648
rect 17684 9664 17736 9716
rect 20260 9664 20312 9716
rect 20628 9664 20680 9716
rect 27160 9664 27212 9716
rect 29828 9664 29880 9716
rect 3056 9460 3108 9512
rect 5816 9528 5868 9580
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 18604 9639 18656 9648
rect 18604 9605 18613 9639
rect 18613 9605 18647 9639
rect 18647 9605 18656 9639
rect 18604 9596 18656 9605
rect 25044 9596 25096 9648
rect 25412 9596 25464 9648
rect 15660 9528 15712 9537
rect 4160 9460 4212 9512
rect 4988 9460 5040 9512
rect 12716 9460 12768 9512
rect 15752 9503 15804 9512
rect 15108 9392 15160 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 8852 9324 8904 9376
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 16948 9571 17000 9580
rect 16580 9460 16632 9512
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 20076 9528 20128 9580
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 18144 9460 18196 9512
rect 19064 9460 19116 9512
rect 20812 9460 20864 9512
rect 22836 9503 22888 9512
rect 19340 9392 19392 9444
rect 20720 9392 20772 9444
rect 22836 9469 22845 9503
rect 22845 9469 22879 9503
rect 22879 9469 22888 9503
rect 22836 9460 22888 9469
rect 23664 9503 23716 9512
rect 23664 9469 23673 9503
rect 23673 9469 23707 9503
rect 23707 9469 23716 9503
rect 23664 9460 23716 9469
rect 26424 9571 26476 9580
rect 26424 9537 26433 9571
rect 26433 9537 26467 9571
rect 26467 9537 26476 9571
rect 26424 9528 26476 9537
rect 27344 9571 27396 9580
rect 26976 9460 27028 9512
rect 27344 9537 27353 9571
rect 27353 9537 27387 9571
rect 27387 9537 27396 9571
rect 27344 9528 27396 9537
rect 29368 9596 29420 9648
rect 30196 9596 30248 9648
rect 32128 9639 32180 9648
rect 32128 9605 32137 9639
rect 32137 9605 32171 9639
rect 32171 9605 32180 9639
rect 32128 9596 32180 9605
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 29552 9528 29604 9580
rect 35440 9528 35492 9580
rect 33232 9460 33284 9512
rect 35348 9503 35400 9512
rect 23388 9392 23440 9444
rect 27344 9392 27396 9444
rect 32404 9435 32456 9444
rect 32404 9401 32413 9435
rect 32413 9401 32447 9435
rect 32447 9401 32456 9435
rect 32404 9392 32456 9401
rect 16580 9324 16632 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 17132 9367 17184 9376
rect 16672 9324 16724 9333
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 25320 9324 25372 9376
rect 26148 9324 26200 9376
rect 30288 9324 30340 9376
rect 32588 9367 32640 9376
rect 32588 9333 32597 9367
rect 32597 9333 32631 9367
rect 32631 9333 32640 9367
rect 32588 9324 32640 9333
rect 34612 9324 34664 9376
rect 35348 9469 35357 9503
rect 35357 9469 35391 9503
rect 35391 9469 35400 9503
rect 35348 9460 35400 9469
rect 35992 9324 36044 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 3056 9120 3108 9172
rect 5356 9120 5408 9172
rect 8208 9163 8260 9172
rect 1400 9095 1452 9104
rect 1400 9061 1409 9095
rect 1409 9061 1443 9095
rect 1443 9061 1452 9095
rect 1400 9052 1452 9061
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 1584 8916 1636 8968
rect 5264 8984 5316 9036
rect 5540 8984 5592 9036
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 15752 9120 15804 9172
rect 16856 9120 16908 9172
rect 20536 9163 20588 9172
rect 20536 9129 20545 9163
rect 20545 9129 20579 9163
rect 20579 9129 20588 9163
rect 20536 9120 20588 9129
rect 26976 9163 27028 9172
rect 26976 9129 26985 9163
rect 26985 9129 27019 9163
rect 27019 9129 27028 9163
rect 26976 9120 27028 9129
rect 29000 9163 29052 9172
rect 29000 9129 29009 9163
rect 29009 9129 29043 9163
rect 29043 9129 29052 9163
rect 29000 9120 29052 9129
rect 29460 9120 29512 9172
rect 35440 9120 35492 9172
rect 15108 9052 15160 9104
rect 19432 9052 19484 9104
rect 18512 8984 18564 9036
rect 32680 8984 32732 9036
rect 5080 8916 5132 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 2412 8848 2464 8900
rect 5632 8848 5684 8900
rect 7288 8848 7340 8900
rect 8208 8916 8260 8968
rect 26148 8959 26200 8968
rect 26148 8925 26157 8959
rect 26157 8925 26191 8959
rect 26191 8925 26200 8959
rect 26148 8916 26200 8925
rect 27436 8916 27488 8968
rect 29092 8916 29144 8968
rect 34612 8916 34664 8968
rect 35348 8984 35400 9036
rect 34888 8959 34940 8968
rect 34888 8925 34897 8959
rect 34897 8925 34931 8959
rect 34931 8925 34940 8959
rect 34888 8916 34940 8925
rect 30472 8848 30524 8900
rect 30656 8848 30708 8900
rect 34428 8848 34480 8900
rect 35900 8916 35952 8968
rect 25964 8823 26016 8832
rect 25964 8789 25973 8823
rect 25973 8789 26007 8823
rect 26007 8789 26016 8823
rect 25964 8780 26016 8789
rect 26332 8823 26384 8832
rect 26332 8789 26341 8823
rect 26341 8789 26375 8823
rect 26375 8789 26384 8823
rect 26332 8780 26384 8789
rect 29000 8780 29052 8832
rect 35532 8780 35584 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 8852 8619 8904 8628
rect 8852 8585 8861 8619
rect 8861 8585 8895 8619
rect 8895 8585 8904 8619
rect 8852 8576 8904 8585
rect 3424 8508 3476 8560
rect 15660 8576 15712 8628
rect 29092 8619 29144 8628
rect 29092 8585 29101 8619
rect 29101 8585 29135 8619
rect 29135 8585 29144 8619
rect 29092 8576 29144 8585
rect 30012 8576 30064 8628
rect 30472 8576 30524 8628
rect 30748 8619 30800 8628
rect 30748 8585 30757 8619
rect 30757 8585 30791 8619
rect 30791 8585 30800 8619
rect 30748 8576 30800 8585
rect 34888 8576 34940 8628
rect 5724 8440 5776 8492
rect 5816 8440 5868 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 11980 8508 12032 8560
rect 22928 8508 22980 8560
rect 24492 8508 24544 8560
rect 29000 8508 29052 8560
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 24308 8440 24360 8492
rect 29644 8440 29696 8492
rect 30104 8483 30156 8492
rect 30104 8449 30113 8483
rect 30113 8449 30147 8483
rect 30147 8449 30156 8483
rect 30104 8440 30156 8449
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 32588 8508 32640 8560
rect 8024 8372 8076 8424
rect 8852 8372 8904 8424
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 27528 8372 27580 8424
rect 11060 8304 11112 8356
rect 23388 8304 23440 8356
rect 26332 8304 26384 8356
rect 30012 8304 30064 8356
rect 35900 8440 35952 8492
rect 33692 8372 33744 8424
rect 34428 8415 34480 8424
rect 34428 8381 34437 8415
rect 34437 8381 34471 8415
rect 34471 8381 34480 8415
rect 34428 8372 34480 8381
rect 34336 8304 34388 8356
rect 37832 8304 37884 8356
rect 3700 8279 3752 8288
rect 3700 8245 3709 8279
rect 3709 8245 3743 8279
rect 3743 8245 3752 8279
rect 3700 8236 3752 8245
rect 7840 8279 7892 8288
rect 7840 8245 7849 8279
rect 7849 8245 7883 8279
rect 7883 8245 7892 8279
rect 7840 8236 7892 8245
rect 9220 8236 9272 8288
rect 17592 8236 17644 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2504 8032 2556 8084
rect 5724 8032 5776 8084
rect 6644 8075 6696 8084
rect 6644 8041 6653 8075
rect 6653 8041 6687 8075
rect 6687 8041 6696 8075
rect 6644 8032 6696 8041
rect 7840 8032 7892 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 26332 8032 26384 8084
rect 3700 7896 3752 7948
rect 8300 7964 8352 8016
rect 14004 7964 14056 8016
rect 8024 7939 8076 7948
rect 8024 7905 8033 7939
rect 8033 7905 8067 7939
rect 8067 7905 8076 7939
rect 8024 7896 8076 7905
rect 8852 7896 8904 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 24860 7939 24912 7948
rect 24860 7905 24869 7939
rect 24869 7905 24903 7939
rect 24903 7905 24912 7939
rect 25320 7939 25372 7948
rect 24860 7896 24912 7905
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 6644 7828 6696 7880
rect 7380 7828 7432 7880
rect 7748 7828 7800 7880
rect 8208 7871 8260 7880
rect 3608 7760 3660 7812
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 9680 7828 9732 7880
rect 14004 7828 14056 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 20720 7871 20772 7880
rect 20720 7837 20729 7871
rect 20729 7837 20763 7871
rect 20763 7837 20772 7871
rect 20720 7828 20772 7837
rect 22100 7828 22152 7880
rect 25964 7828 26016 7880
rect 30012 7760 30064 7812
rect 8208 7692 8260 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 10600 7692 10652 7744
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 16764 7692 16816 7701
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3608 7531 3660 7540
rect 3608 7497 3617 7531
rect 3617 7497 3651 7531
rect 3651 7497 3660 7531
rect 3608 7488 3660 7497
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 7748 7463 7800 7472
rect 7748 7429 7757 7463
rect 7757 7429 7791 7463
rect 7791 7429 7800 7463
rect 7748 7420 7800 7429
rect 8392 7420 8444 7472
rect 14004 7463 14056 7472
rect 14004 7429 14013 7463
rect 14013 7429 14047 7463
rect 14047 7429 14056 7463
rect 14004 7420 14056 7429
rect 17592 7463 17644 7472
rect 17592 7429 17601 7463
rect 17601 7429 17635 7463
rect 17635 7429 17644 7463
rect 17592 7420 17644 7429
rect 18880 7420 18932 7472
rect 26884 7420 26936 7472
rect 27528 7420 27580 7472
rect 30104 7420 30156 7472
rect 30472 7420 30524 7472
rect 5724 7352 5776 7404
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 8208 7352 8260 7404
rect 4712 7284 4764 7336
rect 5356 7284 5408 7336
rect 7656 7284 7708 7336
rect 3424 7216 3476 7268
rect 13820 7284 13872 7336
rect 14372 7284 14424 7336
rect 17960 7284 18012 7336
rect 30748 7395 30800 7404
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 18144 7216 18196 7268
rect 23388 7327 23440 7336
rect 23388 7293 23397 7327
rect 23397 7293 23431 7327
rect 23431 7293 23440 7327
rect 27252 7327 27304 7336
rect 23388 7284 23440 7293
rect 27252 7293 27261 7327
rect 27261 7293 27295 7327
rect 27295 7293 27304 7327
rect 27252 7284 27304 7293
rect 30104 7284 30156 7336
rect 30748 7361 30757 7395
rect 30757 7361 30791 7395
rect 30791 7361 30800 7395
rect 30748 7352 30800 7361
rect 30932 7395 30984 7404
rect 30932 7361 30941 7395
rect 30941 7361 30975 7395
rect 30975 7361 30984 7395
rect 30932 7352 30984 7361
rect 31208 7352 31260 7404
rect 34060 7352 34112 7404
rect 34336 7395 34388 7404
rect 34336 7361 34345 7395
rect 34345 7361 34379 7395
rect 34379 7361 34388 7395
rect 34336 7352 34388 7361
rect 32680 7284 32732 7336
rect 37924 7216 37976 7268
rect 4620 7148 4672 7200
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 8668 7148 8720 7200
rect 19432 7148 19484 7200
rect 23112 7148 23164 7200
rect 27252 7148 27304 7200
rect 30932 7148 30984 7200
rect 33048 7148 33100 7200
rect 34520 7148 34572 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4712 6987 4764 6996
rect 4712 6953 4721 6987
rect 4721 6953 4755 6987
rect 4755 6953 4764 6987
rect 4712 6944 4764 6953
rect 4804 6944 4856 6996
rect 5356 6944 5408 6996
rect 7840 6987 7892 6996
rect 7840 6953 7849 6987
rect 7849 6953 7883 6987
rect 7883 6953 7892 6987
rect 7840 6944 7892 6953
rect 30748 6944 30800 6996
rect 34336 6944 34388 6996
rect 34520 6876 34572 6928
rect 35164 6876 35216 6928
rect 4068 6808 4120 6860
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 13820 6808 13872 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4528 6740 4580 6792
rect 8208 6740 8260 6792
rect 8668 6740 8720 6792
rect 12900 6740 12952 6792
rect 15108 6808 15160 6860
rect 16764 6851 16816 6860
rect 16764 6817 16773 6851
rect 16773 6817 16807 6851
rect 16807 6817 16816 6851
rect 16764 6808 16816 6817
rect 19432 6851 19484 6860
rect 4620 6672 4672 6724
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 5172 6672 5224 6681
rect 7748 6715 7800 6724
rect 7748 6681 7757 6715
rect 7757 6681 7791 6715
rect 7791 6681 7800 6715
rect 7748 6672 7800 6681
rect 13268 6672 13320 6724
rect 15936 6740 15988 6792
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 14372 6715 14424 6724
rect 14372 6681 14381 6715
rect 14381 6681 14415 6715
rect 14415 6681 14424 6715
rect 14372 6672 14424 6681
rect 14740 6604 14792 6656
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 16764 6672 16816 6724
rect 19432 6817 19441 6851
rect 19441 6817 19475 6851
rect 19475 6817 19484 6851
rect 19432 6808 19484 6817
rect 20720 6851 20772 6860
rect 20720 6817 20729 6851
rect 20729 6817 20763 6851
rect 20763 6817 20772 6851
rect 20720 6808 20772 6817
rect 23388 6808 23440 6860
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 22100 6740 22152 6792
rect 23940 6740 23992 6792
rect 20168 6672 20220 6724
rect 23572 6672 23624 6724
rect 30472 6808 30524 6860
rect 34060 6808 34112 6860
rect 30380 6783 30432 6792
rect 30380 6749 30389 6783
rect 30389 6749 30423 6783
rect 30423 6749 30432 6783
rect 30380 6740 30432 6749
rect 33048 6740 33100 6792
rect 34152 6783 34204 6792
rect 33876 6715 33928 6724
rect 33876 6681 33885 6715
rect 33885 6681 33919 6715
rect 33919 6681 33928 6715
rect 33876 6672 33928 6681
rect 34152 6749 34161 6783
rect 34161 6749 34195 6783
rect 34195 6749 34204 6783
rect 34152 6740 34204 6749
rect 34612 6808 34664 6860
rect 35808 6851 35860 6860
rect 35808 6817 35817 6851
rect 35817 6817 35851 6851
rect 35851 6817 35860 6851
rect 35808 6808 35860 6817
rect 17040 6604 17092 6656
rect 18512 6604 18564 6656
rect 23204 6604 23256 6656
rect 23480 6604 23532 6656
rect 34060 6647 34112 6656
rect 34060 6613 34069 6647
rect 34069 6613 34103 6647
rect 34103 6613 34112 6647
rect 34060 6604 34112 6613
rect 34704 6647 34756 6656
rect 34704 6613 34713 6647
rect 34713 6613 34747 6647
rect 34747 6613 34756 6647
rect 34704 6604 34756 6613
rect 34888 6672 34940 6724
rect 35164 6783 35216 6792
rect 35164 6749 35173 6783
rect 35173 6749 35207 6783
rect 35207 6749 35216 6783
rect 35164 6740 35216 6749
rect 35348 6783 35400 6792
rect 35348 6749 35357 6783
rect 35357 6749 35391 6783
rect 35391 6749 35400 6783
rect 35348 6740 35400 6749
rect 37740 6647 37792 6656
rect 37740 6613 37749 6647
rect 37749 6613 37783 6647
rect 37783 6613 37792 6647
rect 37740 6604 37792 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 14280 6400 14332 6452
rect 16396 6400 16448 6452
rect 18512 6400 18564 6452
rect 20904 6400 20956 6452
rect 22284 6400 22336 6452
rect 23940 6443 23992 6452
rect 23940 6409 23949 6443
rect 23949 6409 23983 6443
rect 23983 6409 23992 6443
rect 23940 6400 23992 6409
rect 34888 6400 34940 6452
rect 7748 6332 7800 6384
rect 14096 6332 14148 6384
rect 20168 6332 20220 6384
rect 23204 6332 23256 6384
rect 27344 6332 27396 6384
rect 28080 6332 28132 6384
rect 34704 6332 34756 6384
rect 4528 6264 4580 6316
rect 4712 6264 4764 6316
rect 8208 6264 8260 6316
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 19064 6307 19116 6316
rect 19064 6273 19073 6307
rect 19073 6273 19107 6307
rect 19107 6273 19116 6307
rect 19064 6264 19116 6273
rect 33140 6307 33192 6316
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 4896 6196 4948 6248
rect 7840 6196 7892 6248
rect 4804 6128 4856 6180
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 10324 6060 10376 6112
rect 14372 6128 14424 6180
rect 14004 6060 14056 6112
rect 23388 6196 23440 6248
rect 33140 6273 33149 6307
rect 33149 6273 33183 6307
rect 33183 6273 33192 6307
rect 33140 6264 33192 6273
rect 34152 6264 34204 6316
rect 35808 6264 35860 6316
rect 37832 6307 37884 6316
rect 37832 6273 37841 6307
rect 37841 6273 37875 6307
rect 37875 6273 37884 6307
rect 37832 6264 37884 6273
rect 33048 6196 33100 6248
rect 33876 6196 33928 6248
rect 33968 6239 34020 6248
rect 33968 6205 33977 6239
rect 33977 6205 34011 6239
rect 34011 6205 34020 6239
rect 33968 6196 34020 6205
rect 15108 6128 15160 6180
rect 25688 6128 25740 6180
rect 25780 6128 25832 6180
rect 33692 6171 33744 6180
rect 33692 6137 33701 6171
rect 33701 6137 33735 6171
rect 33735 6137 33744 6171
rect 33692 6128 33744 6137
rect 16212 6060 16264 6112
rect 19156 6103 19208 6112
rect 19156 6069 19165 6103
rect 19165 6069 19199 6103
rect 19199 6069 19208 6103
rect 19156 6060 19208 6069
rect 23204 6060 23256 6112
rect 33876 6103 33928 6112
rect 33876 6069 33885 6103
rect 33885 6069 33919 6103
rect 33919 6069 33928 6103
rect 33876 6060 33928 6069
rect 34060 6060 34112 6112
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2688 5899 2740 5908
rect 2688 5865 2697 5899
rect 2697 5865 2731 5899
rect 2731 5865 2740 5899
rect 2688 5856 2740 5865
rect 2872 5856 2924 5908
rect 4804 5899 4856 5908
rect 4804 5865 4813 5899
rect 4813 5865 4847 5899
rect 4847 5865 4856 5899
rect 4804 5856 4856 5865
rect 14004 5856 14056 5908
rect 15936 5856 15988 5908
rect 16856 5856 16908 5908
rect 21180 5856 21232 5908
rect 3424 5788 3476 5840
rect 16396 5788 16448 5840
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 11980 5720 12032 5772
rect 13084 5763 13136 5772
rect 13084 5729 13093 5763
rect 13093 5729 13127 5763
rect 13127 5729 13136 5763
rect 13084 5720 13136 5729
rect 13360 5720 13412 5772
rect 16212 5720 16264 5772
rect 29736 5788 29788 5840
rect 30380 5788 30432 5840
rect 32864 5856 32916 5908
rect 34612 5856 34664 5908
rect 33140 5831 33192 5840
rect 33140 5797 33149 5831
rect 33149 5797 33183 5831
rect 33183 5797 33192 5831
rect 33140 5788 33192 5797
rect 3792 5652 3844 5704
rect 4620 5652 4672 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 8300 5652 8352 5704
rect 15936 5695 15988 5704
rect 4160 5584 4212 5636
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16396 5652 16448 5704
rect 16948 5695 17000 5704
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 19432 5652 19484 5704
rect 22560 5720 22612 5772
rect 22744 5720 22796 5772
rect 23112 5763 23164 5772
rect 23112 5729 23121 5763
rect 23121 5729 23155 5763
rect 23155 5729 23164 5763
rect 23112 5720 23164 5729
rect 33876 5720 33928 5772
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 20904 5652 20956 5704
rect 23204 5695 23256 5704
rect 23204 5661 23213 5695
rect 23213 5661 23247 5695
rect 23247 5661 23256 5695
rect 23204 5652 23256 5661
rect 10600 5584 10652 5636
rect 10784 5627 10836 5636
rect 10784 5593 10793 5627
rect 10793 5593 10827 5627
rect 10827 5593 10836 5627
rect 10784 5584 10836 5593
rect 12900 5584 12952 5636
rect 4620 5516 4672 5568
rect 13084 5516 13136 5568
rect 13636 5516 13688 5568
rect 15936 5516 15988 5568
rect 17040 5584 17092 5636
rect 19064 5584 19116 5636
rect 23296 5584 23348 5636
rect 16764 5516 16816 5568
rect 17408 5516 17460 5568
rect 19984 5516 20036 5568
rect 20720 5516 20772 5568
rect 23572 5652 23624 5704
rect 30104 5695 30156 5704
rect 30104 5661 30113 5695
rect 30113 5661 30147 5695
rect 30147 5661 30156 5695
rect 30104 5652 30156 5661
rect 33140 5652 33192 5704
rect 33232 5695 33284 5704
rect 33232 5661 33241 5695
rect 33241 5661 33275 5695
rect 33275 5661 33284 5695
rect 33232 5652 33284 5661
rect 37740 5584 37792 5636
rect 25136 5516 25188 5568
rect 32220 5516 32272 5568
rect 33324 5516 33376 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2228 5312 2280 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 16212 5312 16264 5364
rect 16948 5312 17000 5364
rect 17132 5312 17184 5364
rect 17960 5312 18012 5364
rect 4160 5287 4212 5296
rect 4160 5253 4169 5287
rect 4169 5253 4203 5287
rect 4203 5253 4212 5287
rect 4160 5244 4212 5253
rect 10324 5287 10376 5296
rect 10324 5253 10333 5287
rect 10333 5253 10367 5287
rect 10367 5253 10376 5287
rect 10324 5244 10376 5253
rect 3976 5176 4028 5228
rect 5172 5176 5224 5228
rect 12348 5244 12400 5296
rect 17040 5287 17092 5296
rect 17040 5253 17049 5287
rect 17049 5253 17083 5287
rect 17083 5253 17092 5287
rect 17040 5244 17092 5253
rect 19156 5244 19208 5296
rect 20812 5287 20864 5296
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 8760 5108 8812 5160
rect 10508 5151 10560 5160
rect 2872 4972 2924 5024
rect 4804 5040 4856 5092
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 13268 5219 13320 5228
rect 10508 5108 10560 5117
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13636 5219 13688 5228
rect 13360 5176 13412 5185
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 14188 5219 14240 5228
rect 13636 5176 13688 5185
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17132 5176 17184 5228
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 18144 5176 18196 5228
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 16212 5108 16264 5160
rect 17040 5108 17092 5160
rect 19432 5108 19484 5160
rect 19984 5176 20036 5228
rect 20536 5219 20588 5228
rect 20536 5185 20545 5219
rect 20545 5185 20579 5219
rect 20579 5185 20588 5219
rect 20536 5176 20588 5185
rect 20812 5253 20821 5287
rect 20821 5253 20855 5287
rect 20855 5253 20864 5287
rect 20812 5244 20864 5253
rect 20260 5108 20312 5160
rect 22284 5312 22336 5364
rect 23112 5312 23164 5364
rect 23480 5287 23532 5296
rect 23480 5253 23489 5287
rect 23489 5253 23523 5287
rect 23523 5253 23532 5287
rect 23480 5244 23532 5253
rect 25136 5355 25188 5364
rect 23296 5219 23348 5228
rect 23296 5185 23305 5219
rect 23305 5185 23339 5219
rect 23339 5185 23348 5219
rect 23296 5176 23348 5185
rect 23572 5219 23624 5228
rect 23572 5185 23581 5219
rect 23581 5185 23615 5219
rect 23615 5185 23624 5219
rect 23572 5176 23624 5185
rect 25136 5321 25145 5355
rect 25145 5321 25179 5355
rect 25179 5321 25188 5355
rect 25136 5312 25188 5321
rect 27620 5312 27672 5364
rect 27344 5287 27396 5296
rect 27344 5253 27353 5287
rect 27353 5253 27387 5287
rect 27387 5253 27396 5287
rect 30840 5312 30892 5364
rect 33232 5312 33284 5364
rect 33968 5312 34020 5364
rect 27344 5244 27396 5253
rect 25964 5219 26016 5228
rect 25964 5185 25973 5219
rect 25973 5185 26007 5219
rect 26007 5185 26016 5219
rect 25964 5176 26016 5185
rect 22744 5151 22796 5160
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 4712 4972 4764 5024
rect 5080 4972 5132 5024
rect 9680 4972 9732 5024
rect 26884 5108 26936 5160
rect 27528 5151 27580 5160
rect 27528 5117 27537 5151
rect 27537 5117 27571 5151
rect 27571 5117 27580 5151
rect 27528 5108 27580 5117
rect 30104 5108 30156 5160
rect 30380 5108 30432 5160
rect 31944 5176 31996 5228
rect 33324 5176 33376 5228
rect 34520 5244 34572 5296
rect 34152 5219 34204 5228
rect 34152 5185 34161 5219
rect 34161 5185 34195 5219
rect 34195 5185 34204 5219
rect 34152 5176 34204 5185
rect 33140 5108 33192 5160
rect 13176 4972 13228 5024
rect 15936 4972 15988 5024
rect 19432 5015 19484 5024
rect 19432 4981 19441 5015
rect 19441 4981 19475 5015
rect 19475 4981 19484 5015
rect 19432 4972 19484 4981
rect 21272 4972 21324 5024
rect 24584 4972 24636 5024
rect 33692 5040 33744 5092
rect 28356 4972 28408 5024
rect 28448 4972 28500 5024
rect 29736 4972 29788 5024
rect 33416 5015 33468 5024
rect 33416 4981 33425 5015
rect 33425 4981 33459 5015
rect 33459 4981 33468 5015
rect 33416 4972 33468 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11888 4768 11940 4820
rect 16764 4811 16816 4820
rect 16764 4777 16773 4811
rect 16773 4777 16807 4811
rect 16807 4777 16816 4811
rect 16764 4768 16816 4777
rect 20168 4768 20220 4820
rect 23572 4768 23624 4820
rect 19064 4700 19116 4752
rect 20260 4700 20312 4752
rect 25780 4768 25832 4820
rect 26884 4811 26936 4820
rect 26884 4777 26893 4811
rect 26893 4777 26927 4811
rect 26927 4777 26936 4811
rect 26884 4768 26936 4777
rect 34152 4811 34204 4820
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 9588 4632 9640 4684
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 4620 4564 4672 4616
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 13268 4632 13320 4684
rect 22560 4675 22612 4684
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 10784 4564 10836 4616
rect 12348 4607 12400 4616
rect 11888 4496 11940 4548
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 14004 4564 14056 4616
rect 15108 4564 15160 4616
rect 22560 4641 22569 4675
rect 22569 4641 22603 4675
rect 22603 4641 22612 4675
rect 22560 4632 22612 4641
rect 34152 4777 34161 4811
rect 34161 4777 34195 4811
rect 34195 4777 34204 4811
rect 34152 4768 34204 4777
rect 17040 4564 17092 4616
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 19248 4607 19300 4616
rect 4620 4428 4672 4480
rect 8392 4428 8444 4480
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 15752 4496 15804 4548
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22744 4607 22796 4616
rect 19340 4496 19392 4548
rect 22100 4496 22152 4548
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 27344 4675 27396 4684
rect 27344 4641 27353 4675
rect 27353 4641 27387 4675
rect 27387 4641 27396 4675
rect 27344 4632 27396 4641
rect 27528 4675 27580 4684
rect 27528 4641 27537 4675
rect 27537 4641 27571 4675
rect 27571 4641 27580 4675
rect 27528 4632 27580 4641
rect 27620 4564 27672 4616
rect 34796 4700 34848 4752
rect 28448 4607 28500 4616
rect 28448 4573 28457 4607
rect 28457 4573 28491 4607
rect 28491 4573 28500 4607
rect 28448 4564 28500 4573
rect 29184 4564 29236 4616
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 32220 4607 32272 4616
rect 31944 4496 31996 4548
rect 32220 4573 32229 4607
rect 32229 4573 32263 4607
rect 32263 4573 32272 4607
rect 32220 4564 32272 4573
rect 32864 4564 32916 4616
rect 33416 4564 33468 4616
rect 33324 4496 33376 4548
rect 17040 4428 17092 4480
rect 17224 4471 17276 4480
rect 17224 4437 17233 4471
rect 17233 4437 17267 4471
rect 17267 4437 17276 4471
rect 17224 4428 17276 4437
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 28356 4471 28408 4480
rect 28356 4437 28365 4471
rect 28365 4437 28399 4471
rect 28399 4437 28408 4471
rect 28356 4428 28408 4437
rect 29736 4428 29788 4480
rect 32128 4471 32180 4480
rect 32128 4437 32137 4471
rect 32137 4437 32171 4471
rect 32171 4437 32180 4471
rect 32128 4428 32180 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 8300 4267 8352 4276
rect 8300 4233 8309 4267
rect 8309 4233 8343 4267
rect 8343 4233 8352 4267
rect 8300 4224 8352 4233
rect 15752 4267 15804 4276
rect 15752 4233 15761 4267
rect 15761 4233 15795 4267
rect 15795 4233 15804 4267
rect 15752 4224 15804 4233
rect 17040 4224 17092 4276
rect 2872 4199 2924 4208
rect 2872 4165 2881 4199
rect 2881 4165 2915 4199
rect 2915 4165 2924 4199
rect 2872 4156 2924 4165
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 4896 4088 4948 4140
rect 9404 4131 9456 4140
rect 9404 4097 9422 4131
rect 9422 4097 9456 4131
rect 9404 4088 9456 4097
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 15936 4131 15988 4140
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 9864 4020 9916 4072
rect 10876 4020 10928 4072
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 17224 4156 17276 4208
rect 18052 4224 18104 4276
rect 19340 4267 19392 4276
rect 19340 4233 19349 4267
rect 19349 4233 19383 4267
rect 19383 4233 19392 4267
rect 19340 4224 19392 4233
rect 22284 4224 22336 4276
rect 27620 4267 27672 4276
rect 27620 4233 27629 4267
rect 27629 4233 27663 4267
rect 27663 4233 27672 4267
rect 27620 4224 27672 4233
rect 30840 4267 30892 4276
rect 30840 4233 30849 4267
rect 30849 4233 30883 4267
rect 30883 4233 30892 4267
rect 30840 4224 30892 4233
rect 32864 4224 32916 4276
rect 23664 4156 23716 4208
rect 28356 4156 28408 4208
rect 18972 4088 19024 4140
rect 15108 4020 15160 4072
rect 19248 4088 19300 4140
rect 22100 4131 22152 4140
rect 22100 4097 22134 4131
rect 22134 4097 22152 4131
rect 24400 4131 24452 4140
rect 2596 3884 2648 3936
rect 8944 3884 8996 3936
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 12440 3884 12492 3936
rect 19432 4020 19484 4072
rect 17960 3884 18012 3936
rect 22100 4088 22152 4097
rect 24400 4097 24409 4131
rect 24409 4097 24443 4131
rect 24443 4097 24452 4131
rect 24400 4088 24452 4097
rect 29736 4131 29788 4140
rect 29736 4097 29770 4131
rect 29770 4097 29788 4131
rect 29736 4088 29788 4097
rect 24860 4020 24912 4072
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 24676 3884 24728 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 3424 3680 3476 3732
rect 4988 3612 5040 3664
rect 2596 3587 2648 3596
rect 2596 3553 2605 3587
rect 2605 3553 2639 3587
rect 2639 3553 2648 3587
rect 2596 3544 2648 3553
rect 4712 3544 4764 3596
rect 1584 3476 1636 3528
rect 8392 3476 8444 3528
rect 4712 3451 4764 3460
rect 4712 3417 4721 3451
rect 4721 3417 4755 3451
rect 4755 3417 4764 3451
rect 4712 3408 4764 3417
rect 10508 3612 10560 3664
rect 10876 3655 10928 3664
rect 10876 3621 10885 3655
rect 10885 3621 10919 3655
rect 10919 3621 10928 3655
rect 10876 3612 10928 3621
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 11612 3680 11664 3732
rect 14004 3680 14056 3732
rect 17960 3680 18012 3732
rect 13360 3612 13412 3664
rect 24860 3680 24912 3732
rect 25964 3723 26016 3732
rect 25964 3689 25973 3723
rect 25973 3689 26007 3723
rect 26007 3689 26016 3723
rect 25964 3680 26016 3689
rect 29460 3680 29512 3732
rect 31944 3680 31996 3732
rect 12440 3519 12492 3528
rect 12440 3485 12474 3519
rect 12474 3485 12492 3519
rect 12440 3476 12492 3485
rect 24676 3476 24728 3528
rect 32864 3476 32916 3528
rect 20536 3408 20588 3460
rect 32128 3408 32180 3460
rect 10232 3340 10284 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5172 3136 5224 3188
rect 9404 3136 9456 3188
rect 11612 3136 11664 3188
rect 24860 3136 24912 3188
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 10140 3000 10192 3052
rect 1400 2839 1452 2848
rect 1400 2805 1409 2839
rect 1409 2805 1443 2839
rect 1443 2805 1452 2839
rect 1400 2796 1452 2805
rect 1860 2796 1912 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 2872 2592 2924 2644
rect 5264 2524 5316 2576
rect 2780 2388 2832 2440
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 37740 2388 37792 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 3330 39672 3386 39681
rect 3330 39607 3386 39616
rect 3238 38992 3294 39001
rect 3238 38927 3294 38936
rect 3252 37398 3280 38927
rect 3240 37392 3292 37398
rect 3240 37334 3292 37340
rect 2320 36712 2372 36718
rect 2320 36654 2372 36660
rect 2872 36712 2924 36718
rect 2872 36654 2924 36660
rect 2332 36378 2360 36654
rect 2320 36372 2372 36378
rect 2320 36314 2372 36320
rect 2780 36168 2832 36174
rect 2780 36110 2832 36116
rect 2792 35834 2820 36110
rect 2780 35828 2832 35834
rect 2780 35770 2832 35776
rect 2884 35154 2912 36654
rect 3344 35894 3372 39607
rect 9692 39222 9904 39250
rect 3422 38312 3478 38321
rect 3422 38247 3478 38256
rect 3436 37466 3464 38247
rect 4066 37632 4122 37641
rect 4066 37567 4122 37576
rect 3424 37460 3476 37466
rect 3424 37402 3476 37408
rect 4080 37346 4108 37567
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4080 37318 4200 37346
rect 3974 36952 4030 36961
rect 3974 36887 4030 36896
rect 3988 36310 4016 36887
rect 4172 36718 4200 37318
rect 4160 36712 4212 36718
rect 4160 36654 4212 36660
rect 4712 36712 4764 36718
rect 4712 36654 4764 36660
rect 4620 36576 4672 36582
rect 4620 36518 4672 36524
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 3976 36304 4028 36310
rect 3976 36246 4028 36252
rect 4066 36272 4122 36281
rect 4066 36207 4068 36216
rect 4120 36207 4122 36216
rect 4068 36178 4120 36184
rect 3344 35866 3648 35894
rect 2964 35624 3016 35630
rect 2964 35566 3016 35572
rect 3148 35624 3200 35630
rect 3148 35566 3200 35572
rect 3422 35592 3478 35601
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 2976 34610 3004 35566
rect 3160 34921 3188 35566
rect 3422 35527 3478 35536
rect 3146 34912 3202 34921
rect 3146 34847 3202 34856
rect 3436 34678 3464 35527
rect 3424 34672 3476 34678
rect 3424 34614 3476 34620
rect 2964 34604 3016 34610
rect 2964 34546 3016 34552
rect 2870 34232 2926 34241
rect 2870 34167 2926 34176
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 2412 33992 2464 33998
rect 2412 33934 2464 33940
rect 1412 33590 1440 33934
rect 1400 33584 1452 33590
rect 1398 33552 1400 33561
rect 1452 33552 1454 33561
rect 2424 33522 2452 33934
rect 2504 33856 2556 33862
rect 2504 33798 2556 33804
rect 2596 33856 2648 33862
rect 2596 33798 2648 33804
rect 1398 33487 1454 33496
rect 2412 33516 2464 33522
rect 2412 33458 2464 33464
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1412 32201 1440 32370
rect 1584 32224 1636 32230
rect 1398 32192 1454 32201
rect 1584 32166 1636 32172
rect 1398 32127 1454 32136
rect 1596 31414 1624 32166
rect 1584 31408 1636 31414
rect 1584 31350 1636 31356
rect 1400 31340 1452 31346
rect 1400 31282 1452 31288
rect 1412 30870 1440 31282
rect 2516 31278 2544 33798
rect 2608 33590 2636 33798
rect 2596 33584 2648 33590
rect 2596 33526 2648 33532
rect 2884 33454 2912 34167
rect 2872 33448 2924 33454
rect 2872 33390 2924 33396
rect 3238 31512 3294 31521
rect 3238 31447 3294 31456
rect 2504 31272 2556 31278
rect 2504 31214 2556 31220
rect 2504 31136 2556 31142
rect 2504 31078 2556 31084
rect 2872 31136 2924 31142
rect 2872 31078 2924 31084
rect 1400 30864 1452 30870
rect 1398 30832 1400 30841
rect 1452 30832 1454 30841
rect 1398 30767 1454 30776
rect 2516 29850 2544 31078
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2792 30258 2820 30670
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 2504 29844 2556 29850
rect 2504 29786 2556 29792
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29481 1440 29582
rect 1398 29472 1454 29481
rect 1398 29407 1454 29416
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1412 28121 1440 28494
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1398 28112 1454 28121
rect 1398 28047 1454 28056
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1412 26761 1440 26930
rect 1398 26752 1454 26761
rect 1398 26687 1454 26696
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 25401 1440 25842
rect 1596 25498 1624 28358
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 1584 25492 1636 25498
rect 1584 25434 1636 25440
rect 1398 25392 1454 25401
rect 2792 25362 2820 26726
rect 2884 26234 2912 31078
rect 3252 30598 3280 31447
rect 3240 30592 3292 30598
rect 3240 30534 3292 30540
rect 3252 30190 3280 30534
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 3240 30184 3292 30190
rect 3240 30126 3292 30132
rect 2976 29306 3004 30126
rect 2964 29300 3016 29306
rect 2964 29242 3016 29248
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3252 27606 3280 29106
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3528 28762 3556 29038
rect 3516 28756 3568 28762
rect 3516 28698 3568 28704
rect 3240 27600 3292 27606
rect 3240 27542 3292 27548
rect 3056 26240 3108 26246
rect 2884 26206 3004 26234
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 1398 25327 1454 25336
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2884 25294 2912 25638
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 2872 25288 2924 25294
rect 2872 25230 2924 25236
rect 1964 24818 1992 25230
rect 2412 25220 2464 25226
rect 2412 25162 2464 25168
rect 1952 24812 2004 24818
rect 1952 24754 2004 24760
rect 2424 24410 2452 25162
rect 2412 24404 2464 24410
rect 2412 24346 2464 24352
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 24041 1440 24142
rect 1398 24032 1454 24041
rect 1398 23967 1454 23976
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 2780 23112 2832 23118
rect 2976 23066 3004 26206
rect 3056 26182 3108 26188
rect 3068 26042 3096 26182
rect 3620 26042 3648 35866
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4632 35154 4660 36518
rect 4724 35766 4752 36654
rect 8944 36576 8996 36582
rect 8944 36518 8996 36524
rect 5540 36304 5592 36310
rect 5540 36246 5592 36252
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 5000 35834 5028 36042
rect 5552 36038 5580 36246
rect 6920 36236 6972 36242
rect 6920 36178 6972 36184
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 4988 35828 5040 35834
rect 4988 35770 5040 35776
rect 4712 35760 4764 35766
rect 4712 35702 4764 35708
rect 5172 35692 5224 35698
rect 5172 35634 5224 35640
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 3976 35080 4028 35086
rect 3976 35022 4028 35028
rect 3988 34746 4016 35022
rect 4620 35012 4672 35018
rect 4620 34954 4672 34960
rect 3976 34740 4028 34746
rect 3976 34682 4028 34688
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 3976 33992 4028 33998
rect 3976 33934 4028 33940
rect 3988 33658 4016 33934
rect 3976 33652 4028 33658
rect 3976 33594 4028 33600
rect 4080 33114 4108 34478
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4632 34134 4660 34954
rect 4896 34604 4948 34610
rect 4896 34546 4948 34552
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 4724 34202 4752 34342
rect 4712 34196 4764 34202
rect 4712 34138 4764 34144
rect 4620 34128 4672 34134
rect 4620 34070 4672 34076
rect 4908 33998 4936 34546
rect 4988 34536 5040 34542
rect 4988 34478 5040 34484
rect 5000 34066 5028 34478
rect 5184 34202 5212 35634
rect 5552 35154 5580 35974
rect 6932 35222 6960 36178
rect 7288 35624 7340 35630
rect 7288 35566 7340 35572
rect 7564 35624 7616 35630
rect 7564 35566 7616 35572
rect 7300 35290 7328 35566
rect 7288 35284 7340 35290
rect 7288 35226 7340 35232
rect 6920 35216 6972 35222
rect 6920 35158 6972 35164
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 7576 34746 7604 35566
rect 8956 35154 8984 36518
rect 9588 36100 9640 36106
rect 9588 36042 9640 36048
rect 8944 35148 8996 35154
rect 8944 35090 8996 35096
rect 8576 35012 8628 35018
rect 8576 34954 8628 34960
rect 8588 34746 8616 34954
rect 7564 34740 7616 34746
rect 7564 34682 7616 34688
rect 8576 34740 8628 34746
rect 8576 34682 8628 34688
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 7380 34604 7432 34610
rect 7380 34546 7432 34552
rect 8392 34604 8444 34610
rect 8392 34546 8444 34552
rect 5736 34406 5764 34546
rect 5540 34400 5592 34406
rect 5540 34342 5592 34348
rect 5724 34400 5776 34406
rect 5724 34342 5776 34348
rect 5552 34202 5580 34342
rect 5172 34196 5224 34202
rect 5172 34138 5224 34144
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 4988 34060 5040 34066
rect 4988 34002 5040 34008
rect 4620 33992 4672 33998
rect 4620 33934 4672 33940
rect 4896 33992 4948 33998
rect 4948 33940 5028 33946
rect 4896 33934 5028 33940
rect 4632 33454 4660 33934
rect 4908 33918 5028 33934
rect 5000 33522 5028 33918
rect 4988 33516 5040 33522
rect 4988 33458 5040 33464
rect 5264 33516 5316 33522
rect 5264 33458 5316 33464
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 5000 32910 5028 33458
rect 4988 32904 5040 32910
rect 4618 32872 4674 32881
rect 4988 32846 5040 32852
rect 4618 32807 4674 32816
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 3882 30152 3938 30161
rect 3882 30087 3938 30096
rect 3792 30048 3844 30054
rect 3792 29990 3844 29996
rect 3804 29714 3832 29990
rect 3792 29708 3844 29714
rect 3792 29650 3844 29656
rect 3700 29640 3752 29646
rect 3700 29582 3752 29588
rect 3712 28762 3740 29582
rect 3896 29102 3924 30087
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4632 29714 4660 32807
rect 5000 32026 5028 32846
rect 5276 32842 5304 33458
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5368 32978 5396 33390
rect 5552 33318 5580 34138
rect 5736 33862 5764 34342
rect 5724 33856 5776 33862
rect 5724 33798 5776 33804
rect 5736 33658 5764 33798
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 6092 33380 6144 33386
rect 6092 33322 6144 33328
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5552 33114 5580 33254
rect 5540 33108 5592 33114
rect 5540 33050 5592 33056
rect 5356 32972 5408 32978
rect 5356 32914 5408 32920
rect 5264 32836 5316 32842
rect 5264 32778 5316 32784
rect 5172 32428 5224 32434
rect 5172 32370 5224 32376
rect 4988 32020 5040 32026
rect 4988 31962 5040 31968
rect 5080 30660 5132 30666
rect 5080 30602 5132 30608
rect 5092 30410 5120 30602
rect 5000 30394 5120 30410
rect 5000 30388 5132 30394
rect 5000 30382 5080 30388
rect 4620 29708 4672 29714
rect 4620 29650 4672 29656
rect 4632 29510 4660 29650
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 3884 29096 3936 29102
rect 3884 29038 3936 29044
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 3790 28792 3846 28801
rect 3700 28756 3752 28762
rect 4214 28784 4522 28804
rect 3790 28727 3846 28736
rect 4712 28756 4764 28762
rect 3700 28698 3752 28704
rect 3700 28552 3752 28558
rect 3700 28494 3752 28500
rect 3712 28218 3740 28494
rect 3700 28212 3752 28218
rect 3700 28154 3752 28160
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 3712 27470 3740 28018
rect 3804 27946 3832 28727
rect 4712 28698 4764 28704
rect 4068 28620 4120 28626
rect 4068 28562 4120 28568
rect 3884 28552 3936 28558
rect 3884 28494 3936 28500
rect 3896 28082 3924 28494
rect 4080 28098 4108 28562
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 4172 28150 4200 28494
rect 3988 28082 4108 28098
rect 4160 28144 4212 28150
rect 4160 28086 4212 28092
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3988 28076 4120 28082
rect 3988 28070 4068 28076
rect 3792 27940 3844 27946
rect 3792 27882 3844 27888
rect 3988 27606 4016 28070
rect 4068 28018 4120 28024
rect 4172 27962 4200 28086
rect 4080 27934 4200 27962
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 4080 27554 4108 27934
rect 4724 27878 4752 28698
rect 5000 28558 5028 30382
rect 5080 30330 5132 30336
rect 5080 30252 5132 30258
rect 5080 30194 5132 30200
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 4804 27940 4856 27946
rect 4804 27882 4856 27888
rect 4712 27872 4764 27878
rect 4712 27814 4764 27820
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4724 27674 4752 27814
rect 4712 27668 4764 27674
rect 4712 27610 4764 27616
rect 4080 27526 4200 27554
rect 4172 27470 4200 27526
rect 3700 27464 3752 27470
rect 4160 27464 4212 27470
rect 3700 27406 3752 27412
rect 4066 27432 4122 27441
rect 3712 26790 3740 27406
rect 4160 27406 4212 27412
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4066 27367 4122 27376
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3056 26036 3108 26042
rect 3056 25978 3108 25984
rect 3608 26036 3660 26042
rect 3608 25978 3660 25984
rect 3712 25906 3740 26726
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 3988 26246 4016 26386
rect 3976 26240 4028 26246
rect 3976 26182 4028 26188
rect 4080 26058 4108 27367
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 3988 26030 4108 26058
rect 4526 26072 4582 26081
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3884 25220 3936 25226
rect 3884 25162 3936 25168
rect 3056 25152 3108 25158
rect 3056 25094 3108 25100
rect 2780 23054 2832 23060
rect 1412 22681 1440 23054
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1398 22672 1454 22681
rect 1398 22607 1454 22616
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21321 1440 21490
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 1596 21146 1624 22918
rect 2792 22642 2820 23054
rect 2884 23038 3004 23066
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2884 21298 2912 23038
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2976 22710 3004 22918
rect 2964 22704 3016 22710
rect 2964 22646 3016 22652
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1412 20466 1440 20742
rect 2516 20602 2544 21082
rect 2792 21010 2820 21286
rect 2884 21270 3004 21298
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2504 20596 2556 20602
rect 2504 20538 2556 20544
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1412 19961 1440 20402
rect 1398 19952 1454 19961
rect 1398 19887 1454 19896
rect 1596 18970 1624 20402
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 1872 19854 1900 20266
rect 2516 20262 2544 20538
rect 2608 20466 2636 20878
rect 2792 20466 2820 20946
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 2608 19786 2636 20402
rect 2596 19780 2648 19786
rect 2596 19722 2648 19728
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 19378 1992 19654
rect 2884 19446 2912 20742
rect 2976 20058 3004 21270
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 2976 19854 3004 19994
rect 3068 19990 3096 25094
rect 3422 24712 3478 24721
rect 3422 24647 3478 24656
rect 3436 23594 3464 24647
rect 3424 23588 3476 23594
rect 3344 23548 3424 23576
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3056 19984 3108 19990
rect 3056 19926 3108 19932
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 2976 19174 3004 19790
rect 3068 19310 3096 19926
rect 3252 19854 3280 20198
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 18601 1440 18702
rect 1398 18592 1454 18601
rect 1398 18527 1454 18536
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 17241 1440 17614
rect 1398 17232 1454 17241
rect 1398 17167 1454 17176
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15881 1440 16050
rect 1584 15904 1636 15910
rect 1398 15872 1454 15881
rect 1584 15846 1636 15852
rect 1398 15807 1454 15816
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14521 1440 14962
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1596 14414 1624 15846
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 2516 13530 2544 14554
rect 2608 14482 2636 17750
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2792 16794 2820 17070
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2976 16250 3004 17070
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2792 14414 2820 14758
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 13161 1440 13262
rect 1398 13152 1454 13161
rect 1398 13087 1454 13096
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11801 1440 12174
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 1398 11792 1454 11801
rect 1398 11727 1454 11736
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10441 1440 10610
rect 2412 10464 2464 10470
rect 1398 10432 1454 10441
rect 2412 10406 2464 10412
rect 1398 10367 1454 10376
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9586 2268 9998
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 1412 9110 1440 9522
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1400 9104 1452 9110
rect 1398 9072 1400 9081
rect 1452 9072 1454 9081
rect 1398 9007 1454 9016
rect 1596 8974 1624 9318
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7721 1440 7822
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6361 1440 6734
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 5001 1440 5170
rect 1398 4992 1454 5001
rect 1398 4927 1454 4936
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 3641 1440 4082
rect 1398 3632 1454 3641
rect 1398 3567 1454 3576
rect 1596 3534 1624 6598
rect 2240 5370 2268 9522
rect 2424 8906 2452 10406
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2516 8090 2544 9114
rect 2608 9042 2636 12038
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2884 6914 2912 15914
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3068 14618 3096 15438
rect 3344 14958 3372 23548
rect 3424 23530 3476 23536
rect 3606 23352 3662 23361
rect 3606 23287 3662 23296
rect 3620 22710 3648 23287
rect 3608 22704 3660 22710
rect 3608 22646 3660 22652
rect 3422 21992 3478 22001
rect 3422 21927 3478 21936
rect 3436 21078 3464 21927
rect 3424 21072 3476 21078
rect 3424 21014 3476 21020
rect 3620 19446 3648 22646
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 19854 3832 20198
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3608 19440 3660 19446
rect 3608 19382 3660 19388
rect 3514 19272 3570 19281
rect 3514 19207 3570 19216
rect 3528 18222 3556 19207
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3422 17912 3478 17921
rect 3422 17847 3478 17856
rect 3436 16726 3464 17847
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3422 16552 3478 16561
rect 3422 16487 3478 16496
rect 3436 15978 3464 16487
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3422 15192 3478 15201
rect 3422 15127 3478 15136
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3436 14890 3464 15127
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 2976 10470 3004 14214
rect 3436 13841 3464 14214
rect 3422 13832 3478 13841
rect 3422 13767 3478 13776
rect 3238 12472 3294 12481
rect 3238 12407 3294 12416
rect 3252 10742 3280 12407
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3436 11121 3464 11222
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 10266 3004 10406
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2976 9654 3004 10202
rect 3068 10062 3096 10542
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3068 9518 3096 9998
rect 3160 9994 3188 10610
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3344 9602 3372 10610
rect 3422 9752 3478 9761
rect 3422 9687 3424 9696
rect 3476 9687 3478 9696
rect 3424 9658 3476 9664
rect 3252 9586 3372 9602
rect 3240 9580 3372 9586
rect 3292 9574 3372 9580
rect 3240 9522 3292 9528
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 9178 3096 9454
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3436 8401 3464 8502
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3436 7041 3464 7210
rect 3422 7032 3478 7041
rect 3422 6967 3478 6976
rect 3528 6914 3556 18158
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3620 14414 3648 16050
rect 3804 15570 3832 16526
rect 3896 16182 3924 25162
rect 3988 25106 4016 26030
rect 4526 26007 4582 26016
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 4080 25294 4108 25842
rect 4540 25684 4568 26007
rect 4632 25974 4660 27406
rect 4724 27334 4752 27610
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4620 25968 4672 25974
rect 4620 25910 4672 25916
rect 4724 25702 4752 27270
rect 4816 26450 4844 27882
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4712 25696 4764 25702
rect 4540 25656 4660 25684
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4344 25152 4396 25158
rect 3988 25078 4108 25106
rect 4344 25094 4396 25100
rect 4080 24818 4108 25078
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4356 24750 4384 25094
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4632 22642 4660 25656
rect 4712 25638 4764 25644
rect 4724 25498 4752 25638
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 4816 25362 4844 25774
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4816 24682 4844 25298
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 3974 20632 4030 20641
rect 3974 20567 4030 20576
rect 3988 19786 4016 20567
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4632 19802 4660 22578
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4724 19922 4752 20198
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 3976 19780 4028 19786
rect 4632 19774 4752 19802
rect 3976 19722 4028 19728
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4080 19446 4108 19654
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3620 13938 3648 14350
rect 3896 14346 3924 16118
rect 3988 15570 4016 19382
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4172 19258 4200 19314
rect 4080 19230 4200 19258
rect 4080 18850 4108 19230
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4080 18834 4200 18850
rect 4080 18828 4212 18834
rect 4080 18822 4160 18828
rect 4160 18770 4212 18776
rect 4632 18766 4660 19654
rect 4724 19174 4752 19774
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4724 18086 4752 18770
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 4080 14618 4108 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3896 14006 3924 14282
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 4080 13734 4108 14554
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4172 13870 4200 14418
rect 4632 14074 4660 16050
rect 4816 16046 4844 24618
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4908 19922 4936 20742
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 5000 19514 5028 19858
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 17270 4936 19110
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4724 15094 4752 15846
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4816 14482 4844 15982
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4908 15026 4936 15846
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13462 4108 13670
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3620 12442 3648 12718
rect 4080 12442 4108 13398
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4080 12322 4108 12378
rect 3988 12294 4108 12322
rect 3988 11354 4016 12294
rect 4632 12238 4660 13874
rect 4724 13530 4752 14350
rect 5092 14074 5120 30194
rect 5184 21418 5212 32370
rect 5276 28558 5304 32778
rect 5368 32570 5396 32914
rect 5356 32564 5408 32570
rect 5356 32506 5408 32512
rect 5552 31482 5580 33050
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5644 31890 5672 32846
rect 6104 31890 6132 33322
rect 7392 32570 7420 34546
rect 8404 33114 8432 34546
rect 9036 34536 9088 34542
rect 9036 34478 9088 34484
rect 9220 34536 9272 34542
rect 9220 34478 9272 34484
rect 8944 33992 8996 33998
rect 8944 33934 8996 33940
rect 8760 33856 8812 33862
rect 8760 33798 8812 33804
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8208 33040 8260 33046
rect 8208 32982 8260 32988
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 7380 32564 7432 32570
rect 7380 32506 7432 32512
rect 8128 32502 8156 32778
rect 7288 32496 7340 32502
rect 7288 32438 7340 32444
rect 8116 32496 8168 32502
rect 8116 32438 8168 32444
rect 6276 32360 6328 32366
rect 6276 32302 6328 32308
rect 6184 32292 6236 32298
rect 6184 32234 6236 32240
rect 5632 31884 5684 31890
rect 5632 31826 5684 31832
rect 6092 31884 6144 31890
rect 6092 31826 6144 31832
rect 5816 31748 5868 31754
rect 5816 31690 5868 31696
rect 5828 31482 5856 31690
rect 5540 31476 5592 31482
rect 5540 31418 5592 31424
rect 5816 31476 5868 31482
rect 5816 31418 5868 31424
rect 5540 30796 5592 30802
rect 5540 30738 5592 30744
rect 5552 28626 5580 30738
rect 6196 30734 6224 32234
rect 6288 30802 6316 32302
rect 7196 32224 7248 32230
rect 7196 32166 7248 32172
rect 6368 31340 6420 31346
rect 6368 31282 6420 31288
rect 6380 30938 6408 31282
rect 7104 31272 7156 31278
rect 7104 31214 7156 31220
rect 6368 30932 6420 30938
rect 6368 30874 6420 30880
rect 7012 30864 7064 30870
rect 7012 30806 7064 30812
rect 6276 30796 6328 30802
rect 6276 30738 6328 30744
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 6196 29850 6224 30670
rect 7024 30190 7052 30806
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 6184 29844 6236 29850
rect 6184 29786 6236 29792
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5264 28552 5316 28558
rect 5264 28494 5316 28500
rect 5264 27328 5316 27334
rect 5264 27270 5316 27276
rect 5552 27282 5580 28562
rect 5172 21412 5224 21418
rect 5172 21354 5224 21360
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5092 13870 5120 14010
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4724 12306 4752 13466
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3976 11144 4028 11150
rect 4080 11098 4108 12174
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11830 4200 12038
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4028 11092 4108 11098
rect 3976 11086 4108 11092
rect 3988 11070 4108 11086
rect 4080 10146 4108 11070
rect 4172 10810 4200 11154
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4632 10674 4660 11630
rect 4724 11150 4752 12242
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4816 10198 4844 13806
rect 5184 12594 5212 18702
rect 5276 13326 5304 27270
rect 5552 27254 5672 27282
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5368 22778 5396 23054
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5184 12566 5304 12594
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 11354 4936 12174
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5276 11150 5304 12566
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 4804 10192 4856 10198
rect 4080 10118 4200 10146
rect 4804 10134 4856 10140
rect 4172 9518 4200 10118
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4264 9654 4292 9930
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 7954 3740 8230
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3620 7546 3648 7754
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4632 6914 4660 7142
rect 4724 7002 4752 7278
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 2884 6886 3280 6914
rect 3528 6886 3924 6914
rect 3252 6254 3280 6886
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 2700 5914 2728 6190
rect 2884 5914 2912 6190
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3436 5681 3464 5782
rect 3804 5710 3832 6598
rect 3792 5704 3844 5710
rect 3422 5672 3478 5681
rect 3792 5646 3844 5652
rect 3422 5607 3478 5616
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 4146 2728 4558
rect 2884 4214 2912 4966
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 3896 4078 3924 6886
rect 4540 6886 4660 6914
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 5234 4016 6734
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4080 5166 4108 6802
rect 4540 6798 4568 6886
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6322 4568 6734
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4632 5710 4660 6666
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4724 5710 4752 6258
rect 4816 6186 4844 6938
rect 4908 6338 4936 9590
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5000 6866 5028 9454
rect 5092 8974 5120 10610
rect 5184 10062 5212 11018
rect 5276 10266 5304 11086
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4908 6310 5028 6338
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4816 5914 4844 6122
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4172 5302 4200 5578
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4632 4622 4660 5510
rect 4816 5098 4844 5850
rect 4908 5778 4936 6190
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1412 377 1440 2790
rect 1872 2378 1900 2790
rect 2516 2650 2544 3674
rect 2608 3602 2636 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 2650 2912 2994
rect 3436 2961 3464 3674
rect 4632 3482 4660 4422
rect 4724 3602 4752 4966
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4908 4146 4936 4558
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5000 3670 5028 6310
rect 5092 5114 5120 8910
rect 5184 6730 5212 9998
rect 5368 9178 5396 18022
rect 5460 11150 5488 21354
rect 5552 13394 5580 27066
rect 5644 26382 5672 27254
rect 6656 27130 6684 29582
rect 7116 27470 7144 31214
rect 7208 30870 7236 32166
rect 7300 31414 7328 32438
rect 8220 32230 8248 32982
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8404 32366 8432 32914
rect 8484 32904 8536 32910
rect 8484 32846 8536 32852
rect 8496 32434 8524 32846
rect 8484 32428 8536 32434
rect 8484 32370 8536 32376
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 8300 31952 8352 31958
rect 8300 31894 8352 31900
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 7472 31340 7524 31346
rect 7472 31282 7524 31288
rect 7196 30864 7248 30870
rect 7196 30806 7248 30812
rect 7484 30258 7512 31282
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7288 30184 7340 30190
rect 7288 30126 7340 30132
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 5632 26376 5684 26382
rect 5632 26318 5684 26324
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6932 25974 6960 26318
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5828 24614 5856 24754
rect 6932 24614 6960 25910
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5644 18902 5672 22918
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 21010 5856 21286
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5644 18426 5672 18838
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 11354 5580 13330
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5552 9042 5580 9998
rect 5644 9654 5672 10066
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5234 5212 6054
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5092 5086 5212 5114
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4690 5120 4966
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4632 3466 4752 3482
rect 4632 3460 4764 3466
rect 4632 3454 4712 3460
rect 4712 3402 4764 3408
rect 5184 3194 5212 5086
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 3422 2952 3478 2961
rect 3422 2887 3478 2896
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 5276 2582 5304 8978
rect 5644 8906 5672 9590
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5736 8498 5764 11290
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5920 10130 5948 11086
rect 6288 10538 6316 24550
rect 7116 23798 7144 27406
rect 7300 27334 7328 30126
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 7840 28552 7892 28558
rect 7840 28494 7892 28500
rect 7852 28150 7880 28494
rect 7840 28144 7892 28150
rect 7840 28086 7892 28092
rect 7852 27470 7880 28086
rect 7944 27878 7972 28698
rect 8024 28620 8076 28626
rect 8024 28562 8076 28568
rect 8036 28014 8064 28562
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8220 28082 8248 28494
rect 8312 28150 8340 31894
rect 8392 30116 8444 30122
rect 8392 30058 8444 30064
rect 8404 29306 8432 30058
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8404 28762 8432 29106
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 8496 28218 8524 29582
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8300 28144 8352 28150
rect 8300 28086 8352 28092
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7944 27674 7972 27814
rect 7932 27668 7984 27674
rect 7932 27610 7984 27616
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 7104 23792 7156 23798
rect 7104 23734 7156 23740
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6564 23322 6592 23462
rect 6552 23316 6604 23322
rect 6552 23258 6604 23264
rect 6368 23044 6420 23050
rect 6368 22986 6420 22992
rect 6460 23044 6512 23050
rect 6460 22986 6512 22992
rect 6380 22710 6408 22986
rect 6368 22704 6420 22710
rect 6368 22646 6420 22652
rect 6472 22642 6500 22986
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6472 22030 6500 22578
rect 6564 22438 6592 23258
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6736 23248 6788 23254
rect 6736 23190 6788 23196
rect 6656 22522 6684 23190
rect 6748 23118 6776 23190
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6840 22778 6868 23054
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6736 22568 6788 22574
rect 6656 22516 6736 22522
rect 6656 22510 6788 22516
rect 6656 22494 6776 22510
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6564 22234 6592 22374
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 21554 6500 21966
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6564 21350 6592 22170
rect 6656 22098 6684 22494
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6656 21554 6684 22034
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 6932 21622 6960 21898
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 7024 21554 7052 21830
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6380 20942 6408 21286
rect 6748 21010 6776 21286
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18698 6500 19110
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6472 12442 6500 18634
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6564 17746 6592 18022
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6564 17134 6592 17682
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 16658 6592 17070
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6656 16590 6684 17274
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6472 11762 6500 12378
rect 6564 11898 6592 13262
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 10810 6500 11698
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6748 10674 6776 19382
rect 7116 18766 7144 23734
rect 7208 23730 7236 24142
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7300 22030 7328 26998
rect 7656 26988 7708 26994
rect 7656 26930 7708 26936
rect 7668 25294 7696 26930
rect 7852 26858 7880 27406
rect 7840 26852 7892 26858
rect 7840 26794 7892 26800
rect 7944 26586 7972 27610
rect 8036 27538 8064 27950
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7944 26466 7972 26522
rect 7852 26438 7972 26466
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 7760 25158 7788 25842
rect 7852 25702 7880 26438
rect 8036 26382 8064 27474
rect 8220 27470 8248 28018
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8220 27130 8248 27406
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8220 26382 8248 27066
rect 8312 27062 8340 28086
rect 8772 27062 8800 33798
rect 8956 33114 8984 33934
rect 9048 33522 9076 34478
rect 9232 34202 9260 34478
rect 9600 34202 9628 36042
rect 9220 34196 9272 34202
rect 9220 34138 9272 34144
rect 9588 34196 9640 34202
rect 9588 34138 9640 34144
rect 9036 33516 9088 33522
rect 9036 33458 9088 33464
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8944 31136 8996 31142
rect 8944 31078 8996 31084
rect 8956 30802 8984 31078
rect 8944 30796 8996 30802
rect 8944 30738 8996 30744
rect 9128 30660 9180 30666
rect 9128 30602 9180 30608
rect 9140 29850 9168 30602
rect 9404 30184 9456 30190
rect 9404 30126 9456 30132
rect 9128 29844 9180 29850
rect 9128 29786 9180 29792
rect 8852 29572 8904 29578
rect 8852 29514 8904 29520
rect 8864 29170 8892 29514
rect 9416 29510 9444 30126
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 9036 29096 9088 29102
rect 9036 29038 9088 29044
rect 9048 28762 9076 29038
rect 9036 28756 9088 28762
rect 9036 28698 9088 28704
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 8956 27674 8984 28494
rect 8944 27668 8996 27674
rect 8944 27610 8996 27616
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 8760 27056 8812 27062
rect 8760 26998 8812 27004
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 7932 26308 7984 26314
rect 7932 26250 7984 26256
rect 7944 25906 7972 26250
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 8036 25838 8064 26318
rect 8220 25906 8248 26318
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7392 23322 7420 23598
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7760 23186 7788 25094
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7852 24682 7880 24754
rect 7840 24676 7892 24682
rect 7840 24618 7892 24624
rect 7852 23254 7880 24618
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7668 22642 7696 22986
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22710 7880 22918
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7300 18426 7328 21966
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7392 20262 7420 21558
rect 7944 20466 7972 25230
rect 8036 24954 8064 25774
rect 8312 25294 8340 26182
rect 9128 25832 9180 25838
rect 9128 25774 9180 25780
rect 9140 25498 9168 25774
rect 9588 25764 9640 25770
rect 9588 25706 9640 25712
rect 9600 25498 9628 25706
rect 9128 25492 9180 25498
rect 9128 25434 9180 25440
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8024 24948 8076 24954
rect 8024 24890 8076 24896
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6840 17542 6868 18226
rect 7392 17610 7420 20198
rect 7944 19446 7972 20402
rect 9692 20369 9720 39222
rect 9876 39114 9904 39222
rect 9954 39200 10010 40000
rect 29918 39200 29974 40000
rect 9968 39114 9996 39200
rect 9876 39086 9996 39114
rect 23940 37460 23992 37466
rect 23940 37402 23992 37408
rect 13360 37392 13412 37398
rect 13360 37334 13412 37340
rect 12900 36712 12952 36718
rect 12900 36654 12952 36660
rect 12912 36378 12940 36654
rect 12900 36372 12952 36378
rect 12900 36314 12952 36320
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11808 35154 11836 35566
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 13268 35012 13320 35018
rect 13268 34954 13320 34960
rect 13280 34610 13308 34954
rect 13268 34604 13320 34610
rect 13268 34546 13320 34552
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9784 32570 9812 33934
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 12452 31890 12480 33390
rect 12716 32360 12768 32366
rect 12716 32302 12768 32308
rect 12440 31884 12492 31890
rect 12440 31826 12492 31832
rect 12256 29640 12308 29646
rect 12256 29582 12308 29588
rect 12268 29170 12296 29582
rect 12728 29510 12756 32302
rect 13268 31884 13320 31890
rect 13268 31826 13320 31832
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 13096 30666 13124 31214
rect 13084 30660 13136 30666
rect 13084 30602 13136 30608
rect 13096 30190 13124 30602
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13280 29714 13308 31826
rect 13372 31754 13400 37334
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 14372 36848 14424 36854
rect 14372 36790 14424 36796
rect 13820 36712 13872 36718
rect 13820 36654 13872 36660
rect 13636 36168 13688 36174
rect 13636 36110 13688 36116
rect 13648 35698 13676 36110
rect 13832 36106 13860 36654
rect 13820 36100 13872 36106
rect 13820 36042 13872 36048
rect 13636 35692 13688 35698
rect 13636 35634 13688 35640
rect 13452 35624 13504 35630
rect 13452 35566 13504 35572
rect 13464 34610 13492 35566
rect 13544 35488 13596 35494
rect 13544 35430 13596 35436
rect 13556 35154 13584 35430
rect 14384 35154 14412 36790
rect 16776 35698 16804 37266
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 22204 36786 22232 37198
rect 22192 36780 22244 36786
rect 22192 36722 22244 36728
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22100 36644 22152 36650
rect 22100 36586 22152 36592
rect 18696 36576 18748 36582
rect 18696 36518 18748 36524
rect 18708 36242 18736 36518
rect 22112 36242 22140 36586
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 22100 36236 22152 36242
rect 22100 36178 22152 36184
rect 16856 36100 16908 36106
rect 16856 36042 16908 36048
rect 19340 36100 19392 36106
rect 19340 36042 19392 36048
rect 21824 36100 21876 36106
rect 21824 36042 21876 36048
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15488 35154 15516 35430
rect 16868 35154 16896 36042
rect 18420 36032 18472 36038
rect 18420 35974 18472 35980
rect 17132 35624 17184 35630
rect 17132 35566 17184 35572
rect 13544 35148 13596 35154
rect 13544 35090 13596 35096
rect 14372 35148 14424 35154
rect 14372 35090 14424 35096
rect 15476 35148 15528 35154
rect 15476 35090 15528 35096
rect 16856 35148 16908 35154
rect 16856 35090 16908 35096
rect 14188 35080 14240 35086
rect 14188 35022 14240 35028
rect 13452 34604 13504 34610
rect 13452 34546 13504 34552
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 14108 32502 14136 32846
rect 14096 32496 14148 32502
rect 14096 32438 14148 32444
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13372 31726 13492 31754
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12728 29102 12756 29446
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12452 28626 12480 29038
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 10048 26988 10100 26994
rect 10048 26930 10100 26936
rect 10060 25702 10088 26930
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10612 26450 10640 26726
rect 10796 26450 10824 26726
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 10784 25968 10836 25974
rect 10784 25910 10836 25916
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10796 24750 10824 25910
rect 12084 25906 12112 26318
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 13464 25838 13492 31726
rect 13556 31346 13584 31758
rect 13544 31340 13596 31346
rect 13544 31282 13596 31288
rect 14200 29850 14228 35022
rect 15660 35012 15712 35018
rect 15660 34954 15712 34960
rect 15672 34746 15700 34954
rect 15660 34740 15712 34746
rect 15660 34682 15712 34688
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 15384 34604 15436 34610
rect 15384 34546 15436 34552
rect 14280 33992 14332 33998
rect 14280 33934 14332 33940
rect 14292 33522 14320 33934
rect 14280 33516 14332 33522
rect 14280 33458 14332 33464
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 14292 32434 14320 32778
rect 14844 32502 14872 32914
rect 14832 32496 14884 32502
rect 14832 32438 14884 32444
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 14924 31816 14976 31822
rect 14924 31758 14976 31764
rect 14936 31346 14964 31758
rect 14924 31340 14976 31346
rect 14924 31282 14976 31288
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14476 30258 14504 30670
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14280 30184 14332 30190
rect 14280 30126 14332 30132
rect 14188 29844 14240 29850
rect 14188 29786 14240 29792
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13556 27130 13584 28494
rect 13740 28218 13768 29582
rect 14292 28626 14320 30126
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 15016 29708 15068 29714
rect 15016 29650 15068 29656
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14660 29170 14688 29582
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 14936 29238 14964 29514
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 15028 29102 15056 29650
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 14280 28620 14332 28626
rect 14280 28562 14332 28568
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 14108 27674 14136 28494
rect 14372 28144 14424 28150
rect 14372 28086 14424 28092
rect 14096 27668 14148 27674
rect 14096 27610 14148 27616
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 14016 26926 14044 27338
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14016 26450 14044 26862
rect 14200 26790 14228 27610
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14292 26926 14320 27406
rect 14384 27334 14412 28086
rect 14476 28014 14504 28562
rect 15028 28014 15056 29038
rect 15120 28966 15148 29786
rect 15212 29288 15240 34546
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15304 31414 15332 32302
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15396 29306 15424 34546
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15672 34202 15700 34478
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 16396 34196 16448 34202
rect 16396 34138 16448 34144
rect 16028 34060 16080 34066
rect 16028 34002 16080 34008
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 15856 33046 15884 33934
rect 15844 33040 15896 33046
rect 15844 32982 15896 32988
rect 16040 32978 16068 34002
rect 16120 33924 16172 33930
rect 16120 33866 16172 33872
rect 16028 32972 16080 32978
rect 16028 32914 16080 32920
rect 15752 32360 15804 32366
rect 15752 32302 15804 32308
rect 15764 32026 15792 32302
rect 15752 32020 15804 32026
rect 15752 31962 15804 31968
rect 16040 31890 16068 32914
rect 16132 32910 16160 33866
rect 16408 33046 16436 34138
rect 16580 33448 16632 33454
rect 16580 33390 16632 33396
rect 16592 33114 16620 33390
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16304 33040 16356 33046
rect 16304 32982 16356 32988
rect 16396 33040 16448 33046
rect 16396 32982 16448 32988
rect 16316 32910 16344 32982
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16316 31890 16344 32846
rect 16408 32026 16436 32982
rect 16488 32836 16540 32842
rect 16488 32778 16540 32784
rect 16500 32570 16528 32778
rect 16488 32564 16540 32570
rect 16488 32506 16540 32512
rect 16396 32020 16448 32026
rect 16396 31962 16448 31968
rect 16028 31884 16080 31890
rect 16028 31826 16080 31832
rect 16304 31884 16356 31890
rect 16304 31826 16356 31832
rect 16500 31822 16528 32506
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16684 29714 16712 29990
rect 16672 29708 16724 29714
rect 16672 29650 16724 29656
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 16868 29306 16896 29514
rect 15384 29300 15436 29306
rect 15212 29260 15332 29288
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 15108 28960 15160 28966
rect 15108 28902 15160 28908
rect 15212 28778 15240 29106
rect 15120 28750 15240 28778
rect 15120 28558 15148 28750
rect 15304 28694 15332 29260
rect 15384 29242 15436 29248
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15488 28762 15516 28902
rect 15476 28756 15528 28762
rect 15476 28698 15528 28704
rect 15292 28688 15344 28694
rect 15292 28630 15344 28636
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15120 28082 15148 28494
rect 15384 28484 15436 28490
rect 15384 28426 15436 28432
rect 15396 28150 15424 28426
rect 15384 28144 15436 28150
rect 15384 28086 15436 28092
rect 15108 28076 15160 28082
rect 15108 28018 15160 28024
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 14476 27470 14504 27950
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14384 27062 14412 27270
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14200 26518 14228 26726
rect 14188 26512 14240 26518
rect 14188 26454 14240 26460
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 13268 25832 13320 25838
rect 13268 25774 13320 25780
rect 13452 25832 13504 25838
rect 13452 25774 13504 25780
rect 13280 24818 13308 25774
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23798 11836 24006
rect 13924 23866 13952 24686
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 13176 23792 13228 23798
rect 13176 23734 13228 23740
rect 11612 23656 11664 23662
rect 11612 23598 11664 23604
rect 11624 23322 11652 23598
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 13188 23118 13216 23734
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10336 21010 10364 21966
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21010 10548 21830
rect 11716 21690 11744 22510
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 12728 21554 12756 22918
rect 12912 22778 12940 23054
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12912 22030 12940 22714
rect 13004 22098 13032 23054
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 12164 20868 12216 20874
rect 12164 20810 12216 20816
rect 9678 20360 9734 20369
rect 9678 20295 9734 20304
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 10324 19984 10376 19990
rect 10324 19926 10376 19932
rect 10336 19446 10364 19926
rect 12084 19922 12112 20198
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9048 18970 9076 19110
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7484 17882 7512 18566
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 11150 6868 17478
rect 7392 17338 7420 17546
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7484 17066 7512 17818
rect 7944 17678 7972 18022
rect 8404 17882 8432 18226
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8956 17746 8984 18022
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7760 17202 7788 17274
rect 7944 17202 7972 17614
rect 9048 17338 9076 18906
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9784 18358 9812 18634
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9140 17746 9168 18090
rect 9692 17746 9720 18158
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 16794 7512 17002
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7576 16590 7604 17138
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 15026 7144 16390
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 15706 7236 15982
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7668 15502 7696 16934
rect 7944 16590 7972 17138
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15706 7880 15982
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7760 13938 7788 14758
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7760 12850 7788 13262
rect 7852 12986 7880 14214
rect 7944 14006 7972 14758
rect 8036 14414 8064 16390
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8312 13870 8340 16662
rect 8588 15502 8616 16934
rect 9048 16794 9076 17274
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8680 15094 8708 15302
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8956 14618 8984 14894
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11150 7420 11698
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 6840 10810 6868 11086
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6288 10062 6316 10474
rect 6748 10198 6776 10610
rect 6840 10266 6868 10746
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7484 9654 7512 9998
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 8634 5856 9522
rect 7300 8906 7328 9590
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5828 8498 5856 8570
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5736 8090 5764 8434
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 5736 7410 5764 8026
rect 6656 7886 6684 8026
rect 7392 7886 7420 8910
rect 7668 8498 7696 11834
rect 8220 11354 8248 12038
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8220 11150 8248 11290
rect 8208 11144 8260 11150
rect 8128 11092 8208 11098
rect 8128 11086 8260 11092
rect 8128 11070 8248 11086
rect 8128 10810 8156 11070
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8220 9178 8248 10950
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8220 8974 8248 9114
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 7668 7342 7696 8434
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 8090 7880 8230
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7478 7788 7822
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 5368 7002 5396 7278
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 7760 6730 7788 7414
rect 7852 7206 7880 8026
rect 8036 7954 8064 8366
rect 8312 8022 8340 13806
rect 9600 12918 9628 14282
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11762 9168 12174
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8036 7698 8064 7890
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7750 8248 7822
rect 7944 7670 8064 7698
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 7944 7410 7972 7670
rect 8220 7410 8248 7686
rect 8404 7478 8432 7686
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 7002 7880 7142
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7840 6860 7892 6866
rect 7944 6848 7972 7346
rect 7892 6820 7972 6848
rect 7840 6802 7892 6808
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7760 6390 7788 6666
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7852 6254 7880 6802
rect 8220 6798 8248 7346
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6798 8708 7142
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8220 6322 8248 6598
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 4282 8340 5646
rect 8772 5166 8800 11222
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8864 9382 8892 9930
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8864 8634 8892 9318
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8864 8430 8892 8570
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8864 7954 8892 8366
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 8090 9260 8230
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7546 8892 7890
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 5778 9168 6598
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 9600 4690 9628 12854
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9692 12374 9720 12650
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9784 11286 9812 18294
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 17338 10180 17478
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9692 7886 9720 8434
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9692 4622 9720 4966
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8404 3534 8432 4422
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3602 8984 3878
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 9416 3194 9444 4082
rect 9876 4078 9904 4558
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 10152 3058 10180 3878
rect 10244 3398 10272 14826
rect 10980 11830 11008 19722
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11624 19378 11652 19654
rect 11808 19514 11836 19722
rect 11900 19514 11928 19858
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11992 18426 12020 18634
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15570 11744 15846
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 15026 11284 15438
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14482 11744 14894
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11716 12306 11744 12582
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 11532 11762 11560 12106
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10612 11354 10640 11630
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 11808 11150 11836 12582
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 10062 10456 10406
rect 11900 10062 11928 18158
rect 12176 12374 12204 20810
rect 13004 20398 13032 22034
rect 13188 22030 13216 23054
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13188 21690 13216 21966
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12268 18222 12296 18634
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17202 12388 17614
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12452 14618 12480 19926
rect 13004 19922 13032 20334
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13004 19446 13032 19858
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 13096 19378 13124 19790
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18290 12940 19110
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17270 12572 17478
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15570 12940 15846
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 13280 15094 13308 22510
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13372 19854 13400 21626
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 19446 13400 19790
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17678 13400 18022
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13556 15570 13584 23598
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13832 23322 13860 23462
rect 14108 23322 14136 24142
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 13832 22234 13860 23258
rect 14200 23118 14228 23666
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14476 23186 14504 23598
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14200 22778 14228 23054
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13832 19854 13860 19994
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13832 19174 13860 19790
rect 14016 19446 14044 21490
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14200 21146 14228 21422
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14568 20942 14596 27950
rect 15120 27130 15148 28018
rect 15488 27878 15516 28698
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14752 25906 14780 26930
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 14924 26444 14976 26450
rect 14924 26386 14976 26392
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14660 24206 14688 25230
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14660 21010 14688 24142
rect 14752 22642 14780 25842
rect 14844 25226 14872 26250
rect 14936 25498 14964 26386
rect 15028 26382 15056 26862
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15120 26586 15148 26794
rect 15304 26586 15332 27406
rect 15488 27130 15516 27814
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15476 27124 15528 27130
rect 15476 27066 15528 27072
rect 15108 26580 15160 26586
rect 15108 26522 15160 26528
rect 15292 26580 15344 26586
rect 15292 26522 15344 26528
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 15028 25770 15056 26318
rect 15120 26234 15148 26522
rect 15120 26206 15240 26234
rect 15016 25764 15068 25770
rect 15016 25706 15068 25712
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 15028 25294 15056 25706
rect 15212 25498 15240 26206
rect 15580 25770 15608 27338
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15672 26314 15700 26930
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 15568 25764 15620 25770
rect 15568 25706 15620 25712
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14844 24886 14872 25162
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14844 24342 14872 24822
rect 15212 24614 15240 25434
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15304 24750 15332 25298
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15396 24818 15424 25230
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15304 24410 15332 24686
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 15396 24410 15424 24618
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 14832 24336 14884 24342
rect 14832 24278 14884 24284
rect 14844 23798 14872 24278
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 14832 23792 14884 23798
rect 14832 23734 14884 23740
rect 14844 23118 14872 23734
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14660 20466 14688 20946
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14660 19446 14688 20402
rect 14752 19990 14780 22578
rect 15212 21554 15240 24142
rect 15304 23662 15332 24346
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15672 23118 15700 26250
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15764 24206 15792 25842
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 16040 23118 16068 23462
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 15672 22094 15700 23054
rect 15672 22066 15884 22094
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15212 21010 15240 21490
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15856 20398 15884 22066
rect 16592 21010 16620 29174
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16684 28218 16712 29106
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16868 28082 16896 28494
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 17052 27538 17080 28426
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16868 23186 16896 23462
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 17144 21690 17172 35566
rect 18432 35154 18460 35974
rect 19352 35698 19380 36042
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 21836 35834 21864 36042
rect 21824 35828 21876 35834
rect 21824 35770 21876 35776
rect 22112 35766 22140 36178
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 19064 35624 19116 35630
rect 19064 35566 19116 35572
rect 19076 35290 19104 35566
rect 21744 35290 21772 35634
rect 22388 35290 22416 36654
rect 23480 36236 23532 36242
rect 23480 36178 23532 36184
rect 23492 35698 23520 36178
rect 23952 35894 23980 37402
rect 29932 37262 29960 39200
rect 38014 37904 38070 37913
rect 38014 37839 38070 37848
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 38028 37466 38056 37839
rect 38016 37460 38068 37466
rect 38016 37402 38068 37408
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 29184 37120 29236 37126
rect 29184 37062 29236 37068
rect 25412 36576 25464 36582
rect 25412 36518 25464 36524
rect 25424 36242 25452 36518
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 25596 36100 25648 36106
rect 25596 36042 25648 36048
rect 27252 36100 27304 36106
rect 27252 36042 27304 36048
rect 23860 35866 23980 35894
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 19064 35284 19116 35290
rect 19524 35284 19576 35290
rect 19064 35226 19116 35232
rect 19352 35244 19524 35272
rect 18420 35148 18472 35154
rect 18420 35090 18472 35096
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17972 34134 18000 34546
rect 18052 34536 18104 34542
rect 18052 34478 18104 34484
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 17960 34128 18012 34134
rect 17960 34070 18012 34076
rect 18064 33522 18092 34478
rect 19260 34082 19288 34478
rect 19352 34406 19380 35244
rect 19524 35226 19576 35232
rect 21732 35284 21784 35290
rect 21732 35226 21784 35232
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 20812 35216 20864 35222
rect 20812 35158 20864 35164
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34678 20024 35022
rect 20720 35012 20772 35018
rect 20720 34954 20772 34960
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19352 34202 19380 34342
rect 19340 34196 19392 34202
rect 19340 34138 19392 34144
rect 19260 34054 19380 34082
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 18340 32978 18368 33934
rect 18328 32972 18380 32978
rect 18328 32914 18380 32920
rect 18340 32570 18368 32914
rect 18972 32904 19024 32910
rect 18972 32846 19024 32852
rect 19156 32904 19208 32910
rect 19156 32846 19208 32852
rect 18328 32564 18380 32570
rect 18328 32506 18380 32512
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17788 31958 17816 32370
rect 18984 32230 19012 32846
rect 19168 32434 19196 32846
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 18972 32224 19024 32230
rect 18972 32166 19024 32172
rect 17776 31952 17828 31958
rect 17776 31894 17828 31900
rect 17592 30728 17644 30734
rect 17592 30670 17644 30676
rect 17604 30258 17632 30670
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17684 25832 17736 25838
rect 17684 25774 17736 25780
rect 17696 25498 17724 25774
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17512 24682 17540 25230
rect 17500 24676 17552 24682
rect 17500 24618 17552 24624
rect 17788 22094 17816 31894
rect 18984 31822 19012 32166
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18696 31680 18748 31686
rect 18696 31622 18748 31628
rect 18708 30734 18736 31622
rect 18696 30728 18748 30734
rect 18696 30670 18748 30676
rect 18512 30592 18564 30598
rect 18512 30534 18564 30540
rect 18524 30326 18552 30534
rect 18512 30320 18564 30326
rect 18512 30262 18564 30268
rect 18236 30184 18288 30190
rect 18236 30126 18288 30132
rect 18248 29034 18276 30126
rect 19352 29714 19380 34054
rect 19996 33998 20024 34614
rect 20732 34610 20760 34954
rect 20720 34604 20772 34610
rect 20720 34546 20772 34552
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19996 33114 20024 33934
rect 20364 33522 20392 34342
rect 20732 33590 20760 34546
rect 20824 34542 20852 35158
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 20812 34536 20864 34542
rect 20812 34478 20864 34484
rect 20720 33584 20772 33590
rect 20720 33526 20772 33532
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20352 33380 20404 33386
rect 20352 33322 20404 33328
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 20364 32434 20392 33322
rect 20444 32904 20496 32910
rect 20444 32846 20496 32852
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20364 32298 20392 32370
rect 20456 32366 20484 32846
rect 20732 32570 20760 33526
rect 20824 33454 20852 34478
rect 20812 33448 20864 33454
rect 20812 33390 20864 33396
rect 20824 33114 20852 33390
rect 22204 33114 22232 35022
rect 22480 34746 22508 35634
rect 23860 35630 23888 35866
rect 23848 35624 23900 35630
rect 23848 35566 23900 35572
rect 23860 35018 23888 35566
rect 23848 35012 23900 35018
rect 23848 34954 23900 34960
rect 25044 35012 25096 35018
rect 25044 34954 25096 34960
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 23020 34536 23072 34542
rect 23020 34478 23072 34484
rect 22928 33516 22980 33522
rect 22928 33458 22980 33464
rect 22836 33312 22888 33318
rect 22836 33254 22888 33260
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22008 33040 22060 33046
rect 22008 32982 22060 32988
rect 21732 32972 21784 32978
rect 21732 32914 21784 32920
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 21744 32502 21772 32914
rect 22020 32570 22048 32982
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22008 32564 22060 32570
rect 22008 32506 22060 32512
rect 21732 32496 21784 32502
rect 21732 32438 21784 32444
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20444 32360 20496 32366
rect 20444 32302 20496 32308
rect 20352 32292 20404 32298
rect 20352 32234 20404 32240
rect 19616 32224 19668 32230
rect 19616 32166 19668 32172
rect 19628 32026 19656 32166
rect 19616 32020 19668 32026
rect 19616 31962 19668 31968
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19996 31482 20024 31826
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19996 30938 20024 31418
rect 19984 30932 20036 30938
rect 19984 30874 20036 30880
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19352 29102 19380 29650
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 18236 29028 18288 29034
rect 18236 28970 18288 28976
rect 19984 29028 20036 29034
rect 19984 28970 20036 28976
rect 18248 28626 18276 28970
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 26512 19484 26518
rect 19432 26454 19484 26460
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17972 25906 18000 26318
rect 19444 26314 19472 26454
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17880 24886 17908 25094
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 18156 24682 18184 25230
rect 18248 24750 18276 25910
rect 19444 25838 19472 26250
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 18236 24744 18288 24750
rect 18236 24686 18288 24692
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18248 23798 18276 24686
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18156 22234 18184 22510
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 17788 22066 17908 22094
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 20398 16528 20878
rect 16592 20534 16620 20946
rect 17236 20602 17264 21490
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 15856 19922 15884 20334
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18086 13860 19110
rect 13924 18222 13952 19314
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18290 14044 19110
rect 14384 18630 14412 19246
rect 14660 18834 14688 19382
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 14016 17610 14044 18226
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 16114 13952 16594
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13832 15162 13860 15982
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12360 13938 12388 14554
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13280 14074 13308 14350
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13464 13938 13492 14962
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12452 12238 12480 12786
rect 12544 12782 12572 13670
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12544 12306 12572 12718
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12636 12442 12664 12582
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11218 12296 12038
rect 12544 11694 12572 12242
rect 13096 11762 13124 12582
rect 13188 12102 13216 12854
rect 13464 12850 13492 13874
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13832 12646 13860 13670
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11830 13216 12038
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 13280 11150 13308 11494
rect 13372 11218 13400 11630
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11354 13492 11494
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13556 11150 13584 11766
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11992 9994 12020 11086
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10674 13124 10950
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 6866 10640 7686
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5302 10364 6054
rect 10796 5642 10824 9658
rect 12452 9654 12480 10406
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12728 9518 12756 9998
rect 14016 9654 14044 17070
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 16182 14136 16390
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14108 13870 14136 14894
rect 14200 14346 14228 14962
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14292 14482 14320 14758
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14200 14006 14228 14282
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14292 13734 14320 14418
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11150 14136 11494
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10130 14136 10406
rect 14292 10130 14320 10950
rect 14384 10198 14412 18566
rect 14844 18290 14872 19110
rect 15856 18766 15884 19858
rect 16132 19378 16160 19858
rect 16500 19378 16528 20334
rect 16592 19786 16620 20470
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16684 20058 16712 20198
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16592 19446 16620 19722
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16580 19168 16632 19174
rect 16684 19156 16712 19994
rect 16960 19854 16988 20402
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16960 19378 16988 19790
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16632 19128 16712 19156
rect 16580 19110 16632 19116
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14476 16590 14504 18022
rect 14660 17882 14688 18022
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14844 17678 14872 18226
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15028 17610 15056 18226
rect 15212 18222 15240 18702
rect 16592 18698 16620 19110
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15212 17746 15240 18158
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 15212 14006 15240 17682
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 16590 15608 17478
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 15570 15700 16390
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 15026 15516 15438
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 15948 10130 15976 15982
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11218 16252 11494
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16592 10418 16620 18634
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 14890 16712 15506
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 11218 16712 14826
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16776 13326 16804 14486
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16592 10390 16712 10418
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9722 16620 9862
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 7954 11100 8298
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11992 5778 12020 8502
rect 14016 8022 14044 9590
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15120 9110 15148 9386
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15672 8634 15700 9522
rect 16592 9518 16620 9658
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 15764 9178 15792 9454
rect 16684 9382 16712 10390
rect 16960 9586 16988 19314
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 15366 17172 19110
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 17338 17632 17614
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17788 16794 17816 17070
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17696 14278 17724 14962
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17236 13326 17264 13806
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17420 13394 17448 13466
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17052 11558 17080 12378
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11762 17172 12242
rect 17236 12238 17264 13262
rect 17420 12442 17448 13330
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17512 12442 17540 13194
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 11830 17264 12174
rect 17512 11830 17540 12378
rect 17604 12306 17632 13330
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10266 17264 10542
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17696 9722 17724 14214
rect 17880 12238 17908 22066
rect 18340 21010 18368 22510
rect 19352 22506 19380 22986
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18432 20058 18460 20878
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18156 19174 18184 19858
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17972 16250 18000 17070
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14414 18000 14758
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11898 17908 12174
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 18156 9518 18184 19110
rect 18432 17814 18460 19722
rect 18524 19718 18552 20266
rect 18708 19990 18736 20402
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18524 18358 18552 19654
rect 18708 19514 18736 19926
rect 18800 19854 18828 20198
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18800 18426 18828 19790
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18248 15706 18276 16050
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18524 15502 18552 15982
rect 18616 15586 18644 16118
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18708 15706 18736 15846
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18616 15558 18736 15586
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18524 14958 18552 15438
rect 18708 15434 18736 15558
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18708 14346 18736 15370
rect 18800 14958 18828 17750
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 15434 18920 15846
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18800 13938 18828 14894
rect 18892 14414 18920 15370
rect 18984 15162 19012 19450
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19076 15570 19104 16050
rect 19168 15570 19196 18294
rect 19260 16250 19288 21966
rect 19352 17134 19380 22442
rect 19444 21894 19472 23598
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 21962 20024 28970
rect 20180 28626 20208 29038
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 20088 27674 20116 28494
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 20272 27470 20300 27882
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20168 26852 20220 26858
rect 20168 26794 20220 26800
rect 20180 26586 20208 26794
rect 20168 26580 20220 26586
rect 20168 26522 20220 26528
rect 20364 26234 20392 32234
rect 20456 29034 20484 32302
rect 20548 31958 20576 32370
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 21744 31414 21772 32438
rect 22020 32230 22048 32506
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21468 31142 21496 31282
rect 21456 31136 21508 31142
rect 21456 31078 21508 31084
rect 20812 30932 20864 30938
rect 20812 30874 20864 30880
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 20536 29640 20588 29646
rect 20536 29582 20588 29588
rect 20548 29170 20576 29582
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20444 29028 20496 29034
rect 20444 28970 20496 28976
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20640 27062 20668 27338
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 20640 26450 20668 26998
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20628 26308 20680 26314
rect 20732 26296 20760 29650
rect 20824 28218 20852 30874
rect 21468 30598 21496 31078
rect 21928 30734 21956 31962
rect 22020 30938 22048 32166
rect 22388 31822 22416 32778
rect 22560 32292 22612 32298
rect 22560 32234 22612 32240
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 22100 30864 22152 30870
rect 22100 30806 22152 30812
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 21456 30592 21508 30598
rect 21456 30534 21508 30540
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20824 27826 20852 28154
rect 20824 27798 20944 27826
rect 20812 27668 20864 27674
rect 20812 27610 20864 27616
rect 20824 26790 20852 27610
rect 20916 27470 20944 27798
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 21008 26994 21036 27474
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26586 20852 26726
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 21008 26518 21036 26930
rect 20996 26512 21048 26518
rect 20996 26454 21048 26460
rect 21008 26330 21036 26454
rect 20680 26268 20760 26296
rect 20916 26302 21036 26330
rect 20628 26250 20680 26256
rect 20364 26206 20576 26234
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20456 23730 20484 24142
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21010 20024 21898
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19444 20602 19472 20878
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 20088 20398 20116 20878
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20456 20466 20484 20810
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18984 14414 19012 15098
rect 19076 14958 19104 15506
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14482 19104 14894
rect 19168 14550 19196 15506
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18892 12170 18920 14350
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11150 18552 12038
rect 18892 11218 18920 12106
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10742 18368 10950
rect 19076 10742 19104 12854
rect 19352 11354 19380 16934
rect 19444 13394 19472 20334
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 20180 19378 20208 19858
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18358 20024 19246
rect 20088 18630 20116 19314
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19536 14414 19564 14826
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19996 12918 20024 13262
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 19352 10674 19380 11290
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19996 10674 20024 11222
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 16592 7886 16620 9318
rect 16868 9178 16896 9454
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 17144 8498 17172 9318
rect 18524 9042 18552 9862
rect 18616 9654 18644 10134
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 14016 7478 14044 7822
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 6866 13860 7278
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12912 5642 12940 6734
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4146 10364 4422
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10520 3670 10548 5102
rect 10612 4622 10640 5578
rect 10796 4622 10824 5578
rect 13096 5574 13124 5714
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11900 4826 11928 5170
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 11900 4554 11928 4762
rect 12360 4622 12388 5238
rect 13280 5234 13308 6666
rect 14108 6390 14136 7686
rect 14292 6458 14320 7822
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 6730 14412 7278
rect 16776 6866 16804 7686
rect 17604 7478 17632 8230
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18892 7342 18920 7414
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14384 6186 14412 6666
rect 15120 6662 15148 6802
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 14752 6322 14780 6598
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 15120 6186 15148 6598
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5914 14044 6054
rect 15948 5914 15976 6734
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13372 5234 13400 5714
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5234 13676 5510
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 13188 4146 13216 4966
rect 13280 4690 13308 5170
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3670 10916 4014
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 11624 3738 11652 3878
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 11624 3194 11652 3674
rect 12452 3534 12480 3878
rect 13372 3670 13400 5170
rect 14016 4622 14044 5850
rect 15948 5710 15976 5850
rect 16224 5778 16252 6054
rect 16408 5846 16436 6394
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 5234 15976 5510
rect 16224 5370 16252 5714
rect 16408 5710 16436 5782
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16776 5574 16804 6666
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 14200 5137 14228 5170
rect 16224 5166 16252 5306
rect 16212 5160 16264 5166
rect 14186 5128 14242 5137
rect 16212 5102 16264 5108
rect 14186 5063 14242 5072
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14016 3738 14044 4558
rect 15120 4078 15148 4558
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15764 4282 15792 4490
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15948 4146 15976 4966
rect 16776 4826 16804 5510
rect 16868 5234 16896 5850
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 5370 16988 5646
rect 17052 5642 17080 6598
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 17052 5302 17080 5578
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17144 5234 17172 5306
rect 17222 5264 17278 5273
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17132 5228 17184 5234
rect 17222 5199 17224 5208
rect 17132 5170 17184 5176
rect 17276 5199 17278 5208
rect 17224 5170 17276 5176
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17052 4622 17080 5102
rect 17420 4622 17448 5510
rect 17972 5370 18000 7278
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17972 4570 18000 5306
rect 18156 5234 18184 7210
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 6458 18552 6598
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 19076 6322 19104 9454
rect 19352 9450 19380 9998
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 20088 9586 20116 18566
rect 20180 17610 20208 18702
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 16998 20208 17546
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20180 15502 20208 16390
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 11558 20208 15438
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20272 10742 20300 19382
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 13394 20392 13670
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20456 12442 20484 20402
rect 20548 19854 20576 26206
rect 20916 21434 20944 26302
rect 21100 26234 21128 27406
rect 21008 26206 21128 26234
rect 21008 22098 21036 26206
rect 20996 22094 21048 22098
rect 20996 22092 21128 22094
rect 21048 22066 21128 22092
rect 20996 22034 21048 22040
rect 20916 21418 21036 21434
rect 20916 21412 21048 21418
rect 20916 21406 20996 21412
rect 20996 21354 21048 21360
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20466 20760 20878
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20732 19990 20760 20402
rect 20916 20262 20944 21014
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 20058 20944 20198
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 13938 20760 17478
rect 21008 16114 21036 21354
rect 21100 19802 21128 22066
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21376 21146 21404 21422
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21100 19774 21220 19802
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20824 15162 20852 15438
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 21192 14958 21220 19774
rect 21272 15972 21324 15978
rect 21272 15914 21324 15920
rect 21284 15570 21312 15914
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21376 15026 21404 15506
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21376 14278 21404 14418
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 14006 21404 14214
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20640 13394 20668 13806
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20732 13326 20760 13874
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20824 13530 20852 13670
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 21376 13258 21404 13942
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20272 9722 20300 10678
rect 20548 10266 20576 11154
rect 20640 10606 20668 11290
rect 20824 11014 20852 11494
rect 21468 11354 21496 30534
rect 22112 30326 22140 30806
rect 22204 30734 22232 31622
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22100 30320 22152 30326
rect 22100 30262 22152 30268
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22296 29714 22324 30126
rect 22284 29708 22336 29714
rect 22284 29650 22336 29656
rect 22100 28960 22152 28966
rect 22020 28908 22100 28914
rect 22020 28902 22152 28908
rect 22020 28886 22140 28902
rect 21824 27872 21876 27878
rect 21824 27814 21876 27820
rect 21836 26994 21864 27814
rect 22020 27674 22048 28886
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 22100 27600 22152 27606
rect 22388 27554 22416 31758
rect 22572 31346 22600 32234
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22480 29714 22508 29990
rect 22468 29708 22520 29714
rect 22468 29650 22520 29656
rect 22664 29646 22692 31826
rect 22848 31346 22876 33254
rect 22940 31804 22968 33458
rect 23032 33114 23060 34478
rect 23020 33108 23072 33114
rect 23020 33050 23072 33056
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23112 32836 23164 32842
rect 23112 32778 23164 32784
rect 23124 32434 23152 32778
rect 23308 32434 23336 32846
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23020 31816 23072 31822
rect 22940 31776 23020 31804
rect 23020 31758 23072 31764
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22848 29238 22876 29446
rect 23032 29306 23060 31758
rect 23124 31686 23152 32370
rect 23308 32026 23336 32370
rect 23388 32224 23440 32230
rect 23388 32166 23440 32172
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 23124 31346 23152 31622
rect 23308 31414 23336 31962
rect 23296 31408 23348 31414
rect 23296 31350 23348 31356
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 23400 31142 23428 32166
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 23020 29300 23072 29306
rect 23020 29242 23072 29248
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 22836 29232 22888 29238
rect 22836 29174 22888 29180
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22100 27542 22152 27548
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 22020 27062 22048 27270
rect 22008 27056 22060 27062
rect 22008 26998 22060 27004
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21744 25294 21772 26726
rect 22112 25294 22140 27542
rect 22296 27526 22416 27554
rect 22756 27538 22784 29106
rect 22744 27532 22796 27538
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22204 25498 22232 26250
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22112 24070 22140 24346
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 22112 23730 22140 24006
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20824 10690 20852 10950
rect 20824 10674 21036 10690
rect 20812 10668 21048 10674
rect 20864 10662 20996 10668
rect 20812 10610 20864 10616
rect 20996 10610 21048 10616
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19444 9110 19472 9522
rect 20548 9178 20576 10202
rect 20640 10130 20668 10542
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 10198 20760 10406
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20640 9722 20668 10066
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20732 9450 20760 10134
rect 20824 10062 20852 10610
rect 21560 10198 21588 21490
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 20602 21864 20878
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21914 20360 21970 20369
rect 21914 20295 21916 20304
rect 21968 20295 21970 20304
rect 21916 20266 21968 20272
rect 21928 19854 21956 20266
rect 21916 19848 21968 19854
rect 22112 19802 22140 23666
rect 21916 19790 21968 19796
rect 22020 19774 22140 19802
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21928 18766 21956 18906
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 22020 18290 22048 19774
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22112 18970 22140 19654
rect 22296 19378 22324 27526
rect 22744 27474 22796 27480
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 22388 26586 22416 27406
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22848 26450 22876 27406
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22572 25498 22600 25774
rect 23400 25770 23428 26930
rect 23388 25764 23440 25770
rect 23388 25706 23440 25712
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 23676 25294 23704 29242
rect 23768 28966 23796 31214
rect 23756 28960 23808 28966
rect 23756 28902 23808 28908
rect 23768 25498 23796 28902
rect 23860 26450 23888 34954
rect 25056 34610 25084 34954
rect 25608 34610 25636 36042
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26252 35154 26280 35430
rect 26240 35148 26292 35154
rect 26240 35090 26292 35096
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 24032 34536 24084 34542
rect 24032 34478 24084 34484
rect 24044 33658 24072 34478
rect 27264 34066 27292 36042
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 27712 35488 27764 35494
rect 27712 35430 27764 35436
rect 26332 34060 26384 34066
rect 26332 34002 26384 34008
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 24032 33652 24084 33658
rect 24032 33594 24084 33600
rect 25424 33522 25452 33934
rect 25596 33924 25648 33930
rect 25596 33866 25648 33872
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24872 32502 24900 32846
rect 25320 32836 25372 32842
rect 25320 32778 25372 32784
rect 25332 32570 25360 32778
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 31278 23980 32166
rect 25516 31482 25544 32370
rect 25608 32298 25636 33866
rect 25596 32292 25648 32298
rect 25596 32234 25648 32240
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 23940 31272 23992 31278
rect 23940 31214 23992 31220
rect 26240 31272 26292 31278
rect 26240 31214 26292 31220
rect 23952 30870 23980 31214
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 23940 30864 23992 30870
rect 23940 30806 23992 30812
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29306 24532 29582
rect 24308 29300 24360 29306
rect 24308 29242 24360 29248
rect 24492 29300 24544 29306
rect 24492 29242 24544 29248
rect 24320 29170 24348 29242
rect 24596 29186 24624 31078
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 25412 30796 25464 30802
rect 25412 30738 25464 30744
rect 25424 30190 25452 30738
rect 25412 30184 25464 30190
rect 25412 30126 25464 30132
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 25240 29714 25268 29990
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24504 29158 24624 29186
rect 23848 26444 23900 26450
rect 23848 26386 23900 26392
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23492 24818 23520 25162
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 23186 22968 23462
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22756 22098 22784 22986
rect 22744 22092 22796 22098
rect 23032 22094 23060 24754
rect 23584 24698 23612 25230
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23492 24682 23612 24698
rect 23480 24676 23612 24682
rect 23532 24670 23612 24676
rect 23480 24618 23532 24624
rect 23492 23594 23520 24618
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 22744 22034 22796 22040
rect 22940 22066 23060 22094
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22112 18426 22140 18770
rect 22296 18630 22324 19314
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22388 18766 22416 19110
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22020 17882 22048 18226
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21652 14890 21680 15030
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 21652 12442 21680 14826
rect 21744 14414 21772 15846
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 21928 14618 21956 14758
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21744 13326 21772 14350
rect 21928 13530 21956 14554
rect 22020 14074 22048 14894
rect 22388 14822 22416 15438
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21744 12986 21772 13262
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21928 12646 21956 13466
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22020 12918 22048 13262
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 22112 12782 22140 14418
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21652 12238 21680 12378
rect 22112 12306 22140 12718
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 22204 11218 22232 13126
rect 22284 12640 22336 12646
rect 22388 12628 22416 14758
rect 22480 14618 22508 21966
rect 22940 19446 22968 22066
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23308 20534 23336 20742
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22848 18970 22876 19110
rect 22836 18964 22888 18970
rect 22888 18924 22968 18952
rect 22836 18906 22888 18912
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22848 18358 22876 18634
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22848 17678 22876 18294
rect 22940 18086 22968 18924
rect 23032 18834 23060 19246
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 18290 23060 18770
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23124 18290 23152 18702
rect 23308 18698 23336 19314
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 22928 18080 22980 18086
rect 22928 18022 22980 18028
rect 22940 17882 22968 18022
rect 22928 17876 22980 17882
rect 22928 17818 22980 17824
rect 23032 17814 23060 18226
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23124 17678 23152 18226
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 22848 17338 22876 17614
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 23308 16182 23336 18634
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23492 16114 23520 23530
rect 23676 22094 23704 24822
rect 23768 24614 23796 25434
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23860 22710 23888 26386
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 23940 25968 23992 25974
rect 23940 25910 23992 25916
rect 23952 23186 23980 25910
rect 24412 25906 24440 26318
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24320 25498 24348 25774
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24504 25362 24532 29158
rect 25424 29034 25452 30126
rect 25516 30054 25544 30874
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25596 30660 25648 30666
rect 25596 30602 25648 30608
rect 25608 30326 25636 30602
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 25504 30048 25556 30054
rect 25504 29990 25556 29996
rect 25412 29028 25464 29034
rect 25412 28970 25464 28976
rect 25412 25832 25464 25838
rect 25412 25774 25464 25780
rect 24492 25356 24544 25362
rect 24492 25298 24544 25304
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 24044 24818 24072 25230
rect 24504 24886 24532 25298
rect 24492 24880 24544 24886
rect 24492 24822 24544 24828
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 25424 24682 25452 25774
rect 25412 24676 25464 24682
rect 25412 24618 25464 24624
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 24492 22568 24544 22574
rect 24492 22510 24544 22516
rect 23584 22066 23704 22094
rect 23584 16250 23612 22066
rect 24504 21554 24532 22510
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 25516 21078 25544 29990
rect 25608 29102 25636 30262
rect 25792 30258 25820 30670
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25596 25152 25648 25158
rect 25596 25094 25648 25100
rect 25504 21072 25556 21078
rect 25504 21014 25556 21020
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24412 19514 24440 20878
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 24400 19508 24452 19514
rect 24400 19450 24452 19456
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24320 18970 24348 19314
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24412 18426 24440 19314
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24780 18290 24808 18566
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23768 17202 23796 17478
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23768 16250 23796 16594
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22572 15026 22600 15982
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15502 23336 15846
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23492 15434 23520 16050
rect 23584 15570 23612 16186
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24688 15570 24716 15982
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23584 15094 23612 15506
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 14618 22600 14962
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22572 12850 22600 14554
rect 23400 14482 23428 14758
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23676 14414 23704 15438
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23860 13938 23888 15302
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 24412 13530 24440 14350
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22468 12640 22520 12646
rect 22388 12600 22468 12628
rect 22284 12582 22336 12588
rect 22468 12582 22520 12588
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21928 10198 21956 10542
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19444 6866 19472 7142
rect 20732 6866 20760 7822
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 20180 6390 20208 6666
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19076 5642 19104 6258
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 17972 4542 18092 4570
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17052 4282 17080 4422
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17236 4214 17264 4422
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 17972 3942 18000 4422
rect 18064 4282 18092 4542
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18984 4146 19012 5170
rect 19076 4758 19104 5578
rect 19168 5302 19196 6054
rect 20180 5710 20208 6326
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 19156 5296 19208 5302
rect 19156 5238 19208 5244
rect 19444 5166 19472 5646
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19996 5234 20024 5510
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4146 19288 4558
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 4282 19380 4490
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19444 4078 19472 4966
rect 20180 4826 20208 5646
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20536 5228 20588 5234
rect 20732 5216 20760 5510
rect 20824 5302 20852 9454
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 6458 20944 7686
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20916 5710 20944 6394
rect 21192 5914 21220 9862
rect 22112 7886 22140 10746
rect 22296 10062 22324 12582
rect 22480 12442 22508 12582
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22572 12238 22600 12786
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 10062 23152 12038
rect 23768 11762 23796 12582
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22848 9518 22876 9862
rect 22836 9512 22888 9518
rect 22836 9454 22888 9460
rect 22940 8566 22968 9862
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23388 9444 23440 9450
rect 23388 9386 23440 9392
rect 22928 8560 22980 8566
rect 22928 8502 22980 8508
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22112 6798 22140 7822
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22296 6458 22324 8366
rect 23400 8362 23428 9386
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23400 7342 23428 8298
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 22296 5370 22324 6394
rect 23124 5778 23152 7142
rect 23400 6866 23428 7278
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23216 6390 23244 6598
rect 23204 6384 23256 6390
rect 23204 6326 23256 6332
rect 23400 6254 23428 6802
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20588 5188 20760 5216
rect 20536 5170 20588 5176
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 4758 20300 5102
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17972 3738 18000 3878
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 20548 3466 20576 5170
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21284 4622 21312 4966
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 22112 4146 22140 4490
rect 22296 4282 22324 5306
rect 22572 4690 22600 5714
rect 22756 5166 22784 5714
rect 23124 5370 23152 5714
rect 23216 5710 23244 6054
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23308 5234 23336 5578
rect 23492 5302 23520 6598
rect 23584 5710 23612 6666
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22756 4622 22784 5102
rect 23584 4826 23612 5170
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 23676 4214 23704 9454
rect 24320 8498 24348 12582
rect 24688 12434 24716 15506
rect 24596 12406 24716 12434
rect 24596 10810 24624 12406
rect 25240 12238 25268 19858
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24584 10804 24636 10810
rect 24584 10746 24636 10752
rect 24596 10606 24624 10746
rect 24688 10742 24716 11086
rect 25056 10742 25084 12106
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 25056 9654 25084 10678
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 25332 9382 25360 11086
rect 25424 9654 25452 19722
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25516 14482 25544 15370
rect 25608 14482 25636 25094
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25700 22710 25728 22918
rect 25688 22704 25740 22710
rect 25688 22646 25740 22652
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25700 21894 25728 22034
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25700 9994 25728 21830
rect 25792 20874 25820 30194
rect 26252 30122 26280 31214
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 26068 27130 26096 27406
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26344 26994 26372 34002
rect 27724 33590 27752 35430
rect 28460 35290 28488 35634
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28356 35080 28408 35086
rect 28356 35022 28408 35028
rect 28368 34746 28396 35022
rect 28356 34740 28408 34746
rect 28356 34682 28408 34688
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 28552 33658 28580 34546
rect 28632 33924 28684 33930
rect 28632 33866 28684 33872
rect 28540 33652 28592 33658
rect 28540 33594 28592 33600
rect 28644 33590 28672 33866
rect 27712 33584 27764 33590
rect 27712 33526 27764 33532
rect 28632 33584 28684 33590
rect 28632 33526 28684 33532
rect 27724 32978 27752 33526
rect 28816 33516 28868 33522
rect 28816 33458 28868 33464
rect 28828 33318 28856 33458
rect 29000 33448 29052 33454
rect 29000 33390 29052 33396
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 28816 33312 28868 33318
rect 28816 33254 28868 33260
rect 28368 32978 28396 33254
rect 27712 32972 27764 32978
rect 27712 32914 27764 32920
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 26700 32836 26752 32842
rect 26700 32778 26752 32784
rect 27344 32836 27396 32842
rect 27344 32778 27396 32784
rect 26712 29714 26740 32778
rect 27356 31346 27384 32778
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 27620 31272 27672 31278
rect 27620 31214 27672 31220
rect 27632 30122 27660 31214
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 27620 30116 27672 30122
rect 27620 30058 27672 30064
rect 26700 29708 26752 29714
rect 26700 29650 26752 29656
rect 26332 26988 26384 26994
rect 26332 26930 26384 26936
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26252 26042 26280 26250
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26712 25974 26740 29650
rect 28276 29238 28304 30126
rect 28264 29232 28316 29238
rect 28264 29174 28316 29180
rect 28080 28484 28132 28490
rect 28080 28426 28132 28432
rect 27068 27532 27120 27538
rect 27068 27474 27120 27480
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 26988 27062 27016 27270
rect 26976 27056 27028 27062
rect 26976 26998 27028 27004
rect 26976 26444 27028 26450
rect 26976 26386 27028 26392
rect 26700 25968 26752 25974
rect 26700 25910 26752 25916
rect 26884 25968 26936 25974
rect 26884 25910 26936 25916
rect 26896 25158 26924 25910
rect 26884 25152 26936 25158
rect 26884 25094 26936 25100
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 26252 21010 26280 21898
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 26344 19786 26372 22442
rect 26436 22098 26464 23734
rect 26792 23520 26844 23526
rect 26792 23462 26844 23468
rect 26804 23118 26832 23462
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26896 22642 26924 25094
rect 26884 22636 26936 22642
rect 26884 22578 26936 22584
rect 26424 22092 26476 22098
rect 26988 22094 27016 26386
rect 27080 25838 27108 27474
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27356 26926 27384 27270
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 27172 25906 27200 26862
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 27080 25158 27108 25774
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27172 23322 27200 23666
rect 27160 23316 27212 23322
rect 27160 23258 27212 23264
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 26424 22034 26476 22040
rect 26896 22066 27016 22094
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26332 18896 26384 18902
rect 26332 18838 26384 18844
rect 26344 18426 26372 18838
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26528 17746 26556 18158
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26148 17128 26200 17134
rect 26148 17070 26200 17076
rect 26160 16182 26188 17070
rect 26148 16176 26200 16182
rect 26148 16118 26200 16124
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 12850 25912 13262
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25976 12306 26004 13806
rect 26896 13394 26924 22066
rect 27080 21554 27108 23054
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27080 21010 27108 21490
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 27264 19514 27292 19722
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 26988 18834 27016 19382
rect 26976 18828 27028 18834
rect 26976 18770 27028 18776
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27264 16794 27292 17138
rect 27252 16788 27304 16794
rect 27252 16730 27304 16736
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 26896 12646 26924 13330
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 25700 9761 25728 9930
rect 25686 9752 25742 9761
rect 25686 9687 25742 9696
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 24492 8560 24544 8566
rect 24492 8502 24544 8508
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24504 6866 24532 8502
rect 25332 7954 25360 9318
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23952 6458 23980 6734
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 24596 4622 24624 4966
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 23664 4208 23716 4214
rect 23664 4150 23716 4156
rect 24412 4146 24440 4422
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24872 4078 24900 7890
rect 25700 6186 25728 9687
rect 26436 9586 26464 10474
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 26160 8974 26188 9318
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 25976 7886 26004 8774
rect 26344 8362 26372 8774
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 26344 8090 26372 8298
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 26896 7478 26924 12582
rect 27356 12434 27384 26862
rect 27632 26858 27660 27338
rect 27620 26852 27672 26858
rect 27620 26794 27672 26800
rect 28092 26042 28120 28426
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28184 27674 28212 28018
rect 28172 27668 28224 27674
rect 28172 27610 28224 27616
rect 28368 27334 28396 32914
rect 29012 32366 29040 33390
rect 28632 32360 28684 32366
rect 28632 32302 28684 32308
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 28644 30802 28672 32302
rect 28632 30796 28684 30802
rect 28632 30738 28684 30744
rect 28632 27940 28684 27946
rect 28632 27882 28684 27888
rect 28644 27402 28672 27882
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 28356 27328 28408 27334
rect 28356 27270 28408 27276
rect 28080 26036 28132 26042
rect 28080 25978 28132 25984
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27816 24614 27844 25094
rect 27804 24608 27856 24614
rect 27804 24550 27856 24556
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 27540 22778 27568 23054
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27540 21622 27568 21830
rect 27724 21690 27752 21966
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27448 20398 27476 20742
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27448 18426 27476 20334
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27540 17610 27568 18158
rect 27724 17746 27752 18362
rect 27816 18290 27844 24550
rect 28816 24132 28868 24138
rect 28816 24074 28868 24080
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 27908 22778 27936 23054
rect 27896 22772 27948 22778
rect 27896 22714 27948 22720
rect 28172 22568 28224 22574
rect 28172 22510 28224 22516
rect 28184 20874 28212 22510
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 28276 20874 28304 21286
rect 28552 21146 28580 21490
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28264 20868 28316 20874
rect 28264 20810 28316 20816
rect 28276 20466 28304 20810
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 28828 19922 28856 24074
rect 29012 23866 29040 32302
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 29104 28762 29132 29106
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29196 28506 29224 37062
rect 29932 36922 29960 37198
rect 37648 37120 37700 37126
rect 37648 37062 37700 37068
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 30932 36168 30984 36174
rect 30932 36110 30984 36116
rect 30380 36100 30432 36106
rect 30380 36042 30432 36048
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29472 33658 29500 34546
rect 29460 33652 29512 33658
rect 29460 33594 29512 33600
rect 29564 33590 29592 35974
rect 30392 35834 30420 36042
rect 30380 35828 30432 35834
rect 30380 35770 30432 35776
rect 29644 35692 29696 35698
rect 29644 35634 29696 35640
rect 29656 34746 29684 35634
rect 30944 35630 30972 36110
rect 30932 35624 30984 35630
rect 30932 35566 30984 35572
rect 32588 35624 32640 35630
rect 32588 35566 32640 35572
rect 29644 34740 29696 34746
rect 29644 34682 29696 34688
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 29736 33856 29788 33862
rect 29736 33798 29788 33804
rect 30932 33856 30984 33862
rect 30932 33798 30984 33804
rect 31208 33856 31260 33862
rect 31208 33798 31260 33804
rect 29552 33584 29604 33590
rect 29552 33526 29604 33532
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29472 33386 29500 33458
rect 29460 33380 29512 33386
rect 29460 33322 29512 33328
rect 29368 30660 29420 30666
rect 29368 30602 29420 30608
rect 29276 30184 29328 30190
rect 29276 30126 29328 30132
rect 29288 29306 29316 30126
rect 29276 29300 29328 29306
rect 29276 29242 29328 29248
rect 29196 28478 29316 28506
rect 29288 28422 29316 28478
rect 29276 28416 29328 28422
rect 29276 28358 29328 28364
rect 29288 27334 29316 28358
rect 29276 27328 29328 27334
rect 29276 27270 29328 27276
rect 29288 26994 29316 27270
rect 29276 26988 29328 26994
rect 29276 26930 29328 26936
rect 29092 25764 29144 25770
rect 29092 25706 29144 25712
rect 29104 24954 29132 25706
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 29012 21962 29040 23802
rect 29104 23662 29132 24890
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 28816 19916 28868 19922
rect 28816 19858 28868 19864
rect 29092 19440 29144 19446
rect 29092 19382 29144 19388
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27712 17740 27764 17746
rect 27712 17682 27764 17688
rect 27528 17604 27580 17610
rect 27528 17546 27580 17552
rect 27540 17202 27568 17546
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27632 16590 27660 17478
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 13394 27568 14350
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27724 12918 27752 17682
rect 27816 17678 27844 18022
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 28644 14890 28672 19110
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28828 15026 28856 17614
rect 28920 15502 28948 18702
rect 29104 18426 29132 19382
rect 29092 18420 29144 18426
rect 29092 18362 29144 18368
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 29012 15706 29040 17206
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 29012 15094 29040 15642
rect 29104 15570 29132 18362
rect 29288 17882 29316 26930
rect 29380 26518 29408 30602
rect 29368 26512 29420 26518
rect 29368 26454 29420 26460
rect 29380 26042 29408 26454
rect 29368 26036 29420 26042
rect 29368 25978 29420 25984
rect 29380 25906 29408 25978
rect 29368 25900 29420 25906
rect 29368 25842 29420 25848
rect 29472 22642 29500 33322
rect 29564 32502 29592 33526
rect 29748 33454 29776 33798
rect 30944 33590 30972 33798
rect 31220 33674 31248 33798
rect 31128 33658 31248 33674
rect 31312 33658 31340 34546
rect 32036 34536 32088 34542
rect 32036 34478 32088 34484
rect 31116 33652 31248 33658
rect 31168 33646 31248 33652
rect 31116 33594 31168 33600
rect 30932 33584 30984 33590
rect 30984 33532 31064 33538
rect 30932 33526 31064 33532
rect 30748 33516 30800 33522
rect 30944 33510 31064 33526
rect 30748 33458 30800 33464
rect 29736 33448 29788 33454
rect 29736 33390 29788 33396
rect 30760 32774 30788 33458
rect 31036 32842 31064 33510
rect 31024 32836 31076 32842
rect 31024 32778 31076 32784
rect 30748 32768 30800 32774
rect 30748 32710 30800 32716
rect 29552 32496 29604 32502
rect 29552 32438 29604 32444
rect 30932 31884 30984 31890
rect 30932 31826 30984 31832
rect 30944 31346 30972 31826
rect 31036 31414 31064 32778
rect 31220 31958 31248 33646
rect 31300 33652 31352 33658
rect 31300 33594 31352 33600
rect 31576 32768 31628 32774
rect 31576 32710 31628 32716
rect 31208 31952 31260 31958
rect 31208 31894 31260 31900
rect 31588 31890 31616 32710
rect 32048 32366 32076 34478
rect 32312 34400 32364 34406
rect 32312 34342 32364 34348
rect 32324 33998 32352 34342
rect 32600 34066 32628 35566
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 32588 34060 32640 34066
rect 32588 34002 32640 34008
rect 32312 33992 32364 33998
rect 32312 33934 32364 33940
rect 32496 33380 32548 33386
rect 32496 33322 32548 33328
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32036 32360 32088 32366
rect 32036 32302 32088 32308
rect 31576 31884 31628 31890
rect 31576 31826 31628 31832
rect 31024 31408 31076 31414
rect 31024 31350 31076 31356
rect 31484 31408 31536 31414
rect 31484 31350 31536 31356
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 31392 31204 31444 31210
rect 31392 31146 31444 31152
rect 29644 30660 29696 30666
rect 29644 30602 29696 30608
rect 29656 30258 29684 30602
rect 31404 30326 31432 31146
rect 31496 31142 31524 31350
rect 31484 31136 31536 31142
rect 31484 31078 31536 31084
rect 31392 30320 31444 30326
rect 31392 30262 31444 30268
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30300 28150 30328 30194
rect 31404 28234 31432 30262
rect 31312 28206 31432 28234
rect 30288 28144 30340 28150
rect 30288 28086 30340 28092
rect 30300 26994 30328 28086
rect 30472 28076 30524 28082
rect 30472 28018 30524 28024
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30288 26988 30340 26994
rect 30288 26930 30340 26936
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30392 26450 30420 26726
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30104 25696 30156 25702
rect 30104 25638 30156 25644
rect 30116 25294 30144 25638
rect 30300 25498 30328 26318
rect 30392 26042 30420 26386
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 30288 25492 30340 25498
rect 30288 25434 30340 25440
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 29932 24206 29960 25230
rect 30196 24812 30248 24818
rect 30196 24754 30248 24760
rect 30208 24410 30236 24754
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 30484 24342 30512 28018
rect 30564 27056 30616 27062
rect 30564 26998 30616 27004
rect 30576 26586 30604 26998
rect 30944 26790 30972 28018
rect 30932 26784 30984 26790
rect 30932 26726 30984 26732
rect 30564 26580 30616 26586
rect 30564 26522 30616 26528
rect 31312 25974 31340 28206
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 31404 27674 31432 28018
rect 31392 27668 31444 27674
rect 31392 27610 31444 27616
rect 30564 25968 30616 25974
rect 30564 25910 30616 25916
rect 31300 25968 31352 25974
rect 31300 25910 31352 25916
rect 30472 24336 30524 24342
rect 30472 24278 30524 24284
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29840 23798 29868 24006
rect 29828 23792 29880 23798
rect 29828 23734 29880 23740
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29472 22098 29500 22578
rect 29460 22092 29512 22098
rect 29748 22094 29776 23598
rect 29748 22066 29868 22094
rect 29460 22034 29512 22040
rect 29552 20936 29604 20942
rect 29380 20896 29552 20924
rect 29380 20806 29408 20896
rect 29552 20878 29604 20884
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29380 19378 29408 20742
rect 29736 19780 29788 19786
rect 29736 19722 29788 19728
rect 29748 19514 29776 19722
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29380 18154 29408 19314
rect 29840 19310 29868 22066
rect 29932 21554 29960 24142
rect 30300 23866 30328 24142
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 30024 21486 30052 22578
rect 30484 22094 30512 24278
rect 30392 22066 30512 22094
rect 30392 22030 30420 22066
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 30104 21956 30156 21962
rect 30104 21898 30156 21904
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 30024 19666 30052 21422
rect 30116 20874 30144 21898
rect 30288 21480 30340 21486
rect 30288 21422 30340 21428
rect 30104 20868 30156 20874
rect 30104 20810 30156 20816
rect 30116 20534 30144 20810
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 29932 19638 30052 19666
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29368 18148 29420 18154
rect 29368 18090 29420 18096
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29288 17678 29316 17818
rect 29276 17672 29328 17678
rect 29276 17614 29328 17620
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29380 16046 29408 17070
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29380 15570 29408 15982
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28632 14884 28684 14890
rect 28632 14826 28684 14832
rect 28828 14618 28856 14962
rect 29380 14890 29408 15506
rect 29644 15360 29696 15366
rect 29644 15302 29696 15308
rect 28908 14884 28960 14890
rect 28908 14826 28960 14832
rect 29368 14884 29420 14890
rect 29368 14826 29420 14832
rect 28816 14612 28868 14618
rect 28816 14554 28868 14560
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 28092 13258 28120 14214
rect 28080 13252 28132 13258
rect 28080 13194 28132 13200
rect 27712 12912 27764 12918
rect 27712 12854 27764 12860
rect 27264 12406 27384 12434
rect 27264 12306 27292 12406
rect 27252 12300 27304 12306
rect 27252 12242 27304 12248
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 26988 10810 27016 11018
rect 26976 10804 27028 10810
rect 26976 10746 27028 10752
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27172 9722 27200 10610
rect 27264 10010 27292 12242
rect 27436 12164 27488 12170
rect 27436 12106 27488 12112
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 10130 27384 11630
rect 27448 11286 27476 12106
rect 27436 11280 27488 11286
rect 27436 11222 27488 11228
rect 27448 10810 27476 11222
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27448 10266 27476 10610
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27264 9982 27384 10010
rect 27160 9716 27212 9722
rect 27160 9658 27212 9664
rect 27356 9586 27384 9982
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26988 9178 27016 9454
rect 27356 9450 27384 9522
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 26976 9172 27028 9178
rect 26976 9114 27028 9120
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 27264 7206 27292 7278
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 25688 6180 25740 6186
rect 25688 6122 25740 6128
rect 25780 6180 25832 6186
rect 25780 6122 25832 6128
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25148 5370 25176 5510
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25792 4826 25820 6122
rect 25962 5264 26018 5273
rect 25962 5199 25964 5208
rect 26016 5199 26018 5208
rect 25964 5170 26016 5176
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24688 3534 24716 3878
rect 24872 3738 24900 4014
rect 25976 3738 26004 5170
rect 26884 5160 26936 5166
rect 27264 5137 27292 7142
rect 27356 6390 27384 9386
rect 27448 8974 27476 10202
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27540 8514 27568 9998
rect 28000 9994 28028 10406
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 27448 8486 27568 8514
rect 27448 7324 27476 8486
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27540 7478 27568 8366
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27448 7296 27568 7324
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27344 5296 27396 5302
rect 27344 5238 27396 5244
rect 26884 5102 26936 5108
rect 27250 5128 27306 5137
rect 26896 4826 26924 5102
rect 27250 5063 27306 5072
rect 26884 4820 26936 4826
rect 26884 4762 26936 4768
rect 27356 4690 27384 5238
rect 27540 5166 27568 7296
rect 28092 6390 28120 13194
rect 28816 12912 28868 12918
rect 28816 12854 28868 12860
rect 28828 11694 28856 12854
rect 28920 11898 28948 14826
rect 29656 14414 29684 15302
rect 29736 15088 29788 15094
rect 29736 15030 29788 15036
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29380 13870 29408 14350
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28828 11558 28856 11630
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28816 11552 28868 11558
rect 28816 11494 28868 11500
rect 28080 6384 28132 6390
rect 28080 6326 28132 6332
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27540 4690 27568 5102
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27632 4622 27660 5306
rect 28368 5030 28396 11494
rect 29104 10742 29132 12922
rect 29276 12776 29328 12782
rect 29276 12718 29328 12724
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 28998 9616 29054 9625
rect 28998 9551 29054 9560
rect 29012 9178 29040 9551
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 29104 8974 29132 10678
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 29012 8566 29040 8774
rect 29104 8634 29132 8910
rect 29092 8628 29144 8634
rect 29092 8570 29144 8576
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28460 4622 28488 4966
rect 29196 4622 29224 11698
rect 29288 11218 29316 12718
rect 29380 12434 29408 13806
rect 29748 12986 29776 15030
rect 29932 13938 29960 19638
rect 30116 19530 30144 20470
rect 30300 20398 30328 21422
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30300 19922 30328 20334
rect 30288 19916 30340 19922
rect 30288 19858 30340 19864
rect 30024 19502 30144 19530
rect 30392 19514 30420 20402
rect 30576 19718 30604 25910
rect 30932 24608 30984 24614
rect 30932 24550 30984 24556
rect 30944 24206 30972 24550
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 30852 23798 30880 24142
rect 30840 23792 30892 23798
rect 30840 23734 30892 23740
rect 31496 21146 31524 31078
rect 31484 21140 31536 21146
rect 31484 21082 31536 21088
rect 31024 20868 31076 20874
rect 31024 20810 31076 20816
rect 31036 20602 31064 20810
rect 31024 20596 31076 20602
rect 31024 20538 31076 20544
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 30380 19508 30432 19514
rect 30024 19378 30052 19502
rect 30380 19450 30432 19456
rect 30104 19440 30156 19446
rect 30104 19382 30156 19388
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 30012 19236 30064 19242
rect 30012 19178 30064 19184
rect 30024 18630 30052 19178
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 30024 15910 30052 18566
rect 30116 17746 30144 19382
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30104 17740 30156 17746
rect 30104 17682 30156 17688
rect 30012 15904 30064 15910
rect 30012 15846 30064 15852
rect 30024 15366 30052 15846
rect 30208 15570 30236 19246
rect 30576 18834 30604 19654
rect 31312 19378 31340 19654
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 30564 18828 30616 18834
rect 30564 18770 30616 18776
rect 31312 18698 31340 19314
rect 31588 18766 31616 31826
rect 32048 22778 32076 32302
rect 32416 31482 32444 32370
rect 32404 31476 32456 31482
rect 32404 31418 32456 31424
rect 32508 31346 32536 33322
rect 32600 32434 32628 34002
rect 35348 33924 35400 33930
rect 35348 33866 35400 33872
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32140 30938 32168 31282
rect 32128 30932 32180 30938
rect 32128 30874 32180 30880
rect 32416 30802 32444 31282
rect 32404 30796 32456 30802
rect 32404 30738 32456 30744
rect 32600 30258 32628 32370
rect 33048 32224 33100 32230
rect 33048 32166 33100 32172
rect 33060 31822 33088 32166
rect 33336 32026 33364 32370
rect 34428 32224 34480 32230
rect 34428 32166 34480 32172
rect 33324 32020 33376 32026
rect 33324 31962 33376 31968
rect 33048 31816 33100 31822
rect 33048 31758 33100 31764
rect 34440 31414 34468 32166
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35360 31482 35388 33866
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 34428 31408 34480 31414
rect 34428 31350 34480 31356
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34796 30320 34848 30326
rect 34796 30262 34848 30268
rect 32588 30252 32640 30258
rect 32588 30194 32640 30200
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 32324 28082 32352 28358
rect 34072 28218 34100 30194
rect 34808 29714 34836 30262
rect 35348 30048 35400 30054
rect 35348 29990 35400 29996
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34796 29708 34848 29714
rect 34796 29650 34848 29656
rect 34704 28960 34756 28966
rect 34704 28902 34756 28908
rect 34060 28212 34112 28218
rect 34060 28154 34112 28160
rect 34716 28150 34744 28902
rect 34808 28626 34836 29650
rect 35360 29238 35388 29990
rect 35348 29232 35400 29238
rect 35348 29174 35400 29180
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34704 28144 34756 28150
rect 34704 28086 34756 28092
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 34244 28076 34296 28082
rect 34244 28018 34296 28024
rect 32140 27402 32168 28018
rect 32324 27470 32352 28018
rect 34256 27674 34284 28018
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34428 27872 34480 27878
rect 34428 27814 34480 27820
rect 34244 27668 34296 27674
rect 34244 27610 34296 27616
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 34336 27464 34388 27470
rect 34336 27406 34388 27412
rect 32128 27396 32180 27402
rect 32128 27338 32180 27344
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32036 21888 32088 21894
rect 32036 21830 32088 21836
rect 32048 20942 32076 21830
rect 32140 21146 32168 27338
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 33336 27130 33364 27270
rect 33324 27124 33376 27130
rect 33324 27066 33376 27072
rect 33336 26234 33364 27066
rect 34348 26994 34376 27406
rect 34440 27130 34468 27814
rect 34532 27334 34560 27950
rect 34520 27328 34572 27334
rect 34520 27270 34572 27276
rect 34428 27124 34480 27130
rect 34428 27066 34480 27072
rect 33600 26988 33652 26994
rect 33600 26930 33652 26936
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 33612 26790 33640 26930
rect 33600 26784 33652 26790
rect 33600 26726 33652 26732
rect 33244 26206 33364 26234
rect 32496 24064 32548 24070
rect 32496 24006 32548 24012
rect 32508 23730 32536 24006
rect 32496 23724 32548 23730
rect 32496 23666 32548 23672
rect 32588 21344 32640 21350
rect 32588 21286 32640 21292
rect 32128 21140 32180 21146
rect 32128 21082 32180 21088
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 32048 18766 32076 19722
rect 32140 19514 32168 21082
rect 32312 21072 32364 21078
rect 32312 21014 32364 21020
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 32324 19378 32352 21014
rect 32600 19990 32628 21286
rect 32588 19984 32640 19990
rect 32588 19926 32640 19932
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32140 18970 32168 19314
rect 32128 18964 32180 18970
rect 32128 18906 32180 18912
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 31300 18692 31352 18698
rect 31300 18634 31352 18640
rect 30288 17604 30340 17610
rect 30288 17546 30340 17552
rect 30300 16658 30328 17546
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 31588 16250 31616 18702
rect 31668 18692 31720 18698
rect 31668 18634 31720 18640
rect 31680 17610 31708 18634
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32324 18290 32352 18566
rect 32312 18284 32364 18290
rect 32312 18226 32364 18232
rect 31668 17604 31720 17610
rect 31668 17546 31720 17552
rect 31208 16244 31260 16250
rect 31208 16186 31260 16192
rect 31576 16244 31628 16250
rect 31576 16186 31628 16192
rect 31116 15904 31168 15910
rect 31116 15846 31168 15852
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 31128 15502 31156 15846
rect 31220 15502 31248 16186
rect 32864 16108 32916 16114
rect 32864 16050 32916 16056
rect 32128 15904 32180 15910
rect 32128 15846 32180 15852
rect 32140 15706 32168 15846
rect 32128 15700 32180 15706
rect 32128 15642 32180 15648
rect 31116 15496 31168 15502
rect 31116 15438 31168 15444
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30012 15360 30064 15366
rect 30012 15302 30064 15308
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 29932 13530 29960 13874
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29380 12406 29500 12434
rect 29276 11212 29328 11218
rect 29276 11154 29328 11160
rect 29276 11076 29328 11082
rect 29276 11018 29328 11024
rect 29288 9994 29316 11018
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29276 9988 29328 9994
rect 29276 9930 29328 9936
rect 29288 9586 29316 9930
rect 29380 9654 29408 10610
rect 29472 10266 29500 12406
rect 29748 12306 29776 12922
rect 29736 12300 29788 12306
rect 29736 12242 29788 12248
rect 29748 11898 29776 12242
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 29564 11354 29592 11698
rect 29644 11620 29696 11626
rect 29644 11562 29696 11568
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29656 10742 29684 11562
rect 29748 10810 29776 11834
rect 29932 11830 29960 12106
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29644 10736 29696 10742
rect 29644 10678 29696 10684
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 29656 10198 29684 10678
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 29644 10192 29696 10198
rect 29644 10134 29696 10140
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 29368 9648 29420 9654
rect 29368 9590 29420 9596
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29472 9178 29500 9998
rect 29550 9616 29606 9625
rect 29550 9551 29552 9560
rect 29604 9551 29606 9560
rect 29552 9522 29604 9528
rect 29460 9172 29512 9178
rect 29460 9114 29512 9120
rect 29656 8498 29684 9998
rect 29644 8492 29696 8498
rect 29644 8434 29696 8440
rect 29748 5846 29776 10202
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29840 9722 29868 9998
rect 29828 9716 29880 9722
rect 29828 9658 29880 9664
rect 30024 8634 30052 15302
rect 30300 15094 30328 15370
rect 30288 15088 30340 15094
rect 30288 15030 30340 15036
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 30116 13870 30144 14758
rect 30484 14618 30512 14962
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 30116 11694 30144 13466
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30484 11830 30512 12582
rect 30472 11824 30524 11830
rect 30472 11766 30524 11772
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30104 11688 30156 11694
rect 30104 11630 30156 11636
rect 30300 11150 30328 11698
rect 30484 11354 30512 11766
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30208 9654 30236 10542
rect 30300 10130 30328 10746
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 30024 8362 30052 8570
rect 30300 8498 30328 9318
rect 30668 8906 30696 9862
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30656 8900 30708 8906
rect 30656 8842 30708 8848
rect 30484 8634 30512 8842
rect 30760 8634 30788 9930
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30012 8356 30064 8362
rect 30012 8298 30064 8304
rect 30024 7818 30052 8298
rect 30012 7812 30064 7818
rect 30012 7754 30064 7760
rect 30116 7478 30144 8434
rect 30484 7478 30512 8570
rect 30104 7472 30156 7478
rect 30104 7414 30156 7420
rect 30472 7472 30524 7478
rect 30472 7414 30524 7420
rect 30104 7336 30156 7342
rect 30104 7278 30156 7284
rect 29736 5840 29788 5846
rect 29736 5782 29788 5788
rect 30116 5710 30144 7278
rect 30484 6866 30512 7414
rect 31220 7410 31248 15438
rect 32220 15360 32272 15366
rect 32220 15302 32272 15308
rect 32232 15026 32260 15302
rect 32876 15162 32904 16050
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32600 12442 32628 14010
rect 32588 12436 32640 12442
rect 32588 12378 32640 12384
rect 32600 12238 32628 12378
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 33140 12232 33192 12238
rect 33140 12174 33192 12180
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32416 11218 32444 12038
rect 33152 11830 33180 12174
rect 33140 11824 33192 11830
rect 33140 11766 33192 11772
rect 32680 11552 32732 11558
rect 32680 11494 32732 11500
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32128 9920 32180 9926
rect 32128 9862 32180 9868
rect 32140 9654 32168 9862
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 32416 9450 32444 11154
rect 32404 9444 32456 9450
rect 32404 9386 32456 9392
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32600 8566 32628 9318
rect 32692 9042 32720 11494
rect 33244 10810 33272 26206
rect 33612 25770 33640 26726
rect 34348 25906 34376 26930
rect 34428 26920 34480 26926
rect 34532 26908 34560 27270
rect 34716 26994 34744 28086
rect 35360 28082 35388 29174
rect 35348 28076 35400 28082
rect 35348 28018 35400 28024
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34480 26880 34560 26908
rect 34428 26862 34480 26868
rect 34440 25906 34468 26862
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 34428 25900 34480 25906
rect 34428 25842 34480 25848
rect 34704 25900 34756 25906
rect 34704 25842 34756 25848
rect 33600 25764 33652 25770
rect 33600 25706 33652 25712
rect 34612 25764 34664 25770
rect 34612 25706 34664 25712
rect 34152 25696 34204 25702
rect 34152 25638 34204 25644
rect 34164 24206 34192 25638
rect 34152 24200 34204 24206
rect 34152 24142 34204 24148
rect 34520 23792 34572 23798
rect 34520 23734 34572 23740
rect 33876 23520 33928 23526
rect 33876 23462 33928 23468
rect 33888 22642 33916 23462
rect 34532 23118 34560 23734
rect 34520 23112 34572 23118
rect 34520 23054 34572 23060
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33888 21554 33916 22578
rect 33876 21548 33928 21554
rect 33876 21490 33928 21496
rect 34532 20942 34560 23054
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 33600 18624 33652 18630
rect 33600 18566 33652 18572
rect 33612 18426 33640 18566
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 34532 18358 34560 20878
rect 34520 18352 34572 18358
rect 34520 18294 34572 18300
rect 34520 17604 34572 17610
rect 34520 17546 34572 17552
rect 34532 16046 34560 17546
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 34072 14006 34100 15438
rect 34532 14414 34560 15982
rect 34624 15910 34652 25706
rect 34716 22710 34744 25842
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 24608 34848 24614
rect 34796 24550 34848 24556
rect 34808 24206 34836 24550
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34808 23662 34836 24142
rect 34888 24132 34940 24138
rect 34888 24074 34940 24080
rect 34900 23730 34928 24074
rect 34888 23724 34940 23730
rect 34888 23666 34940 23672
rect 34796 23656 34848 23662
rect 34796 23598 34848 23604
rect 34704 22704 34756 22710
rect 34704 22646 34756 22652
rect 34716 20466 34744 22646
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34716 19378 34744 19654
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34716 17202 34744 18226
rect 34808 18170 34836 23598
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35452 20466 35480 31078
rect 36452 29572 36504 29578
rect 36452 29514 36504 29520
rect 35808 29504 35860 29510
rect 35808 29446 35860 29452
rect 35820 29170 35848 29446
rect 36464 29306 36492 29514
rect 37372 29504 37424 29510
rect 37372 29446 37424 29452
rect 36452 29300 36504 29306
rect 36452 29242 36504 29248
rect 37384 29170 37412 29446
rect 35808 29164 35860 29170
rect 35808 29106 35860 29112
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 37372 29164 37424 29170
rect 37372 29106 37424 29112
rect 35624 28484 35676 28490
rect 35624 28426 35676 28432
rect 35532 28076 35584 28082
rect 35532 28018 35584 28024
rect 35544 27538 35572 28018
rect 35636 27674 35664 28426
rect 35624 27668 35676 27674
rect 35624 27610 35676 27616
rect 35532 27532 35584 27538
rect 35532 27474 35584 27480
rect 35544 26858 35572 27474
rect 35820 27470 35848 29106
rect 35900 29096 35952 29102
rect 35900 29038 35952 29044
rect 35912 28370 35940 29038
rect 36004 28762 36032 29106
rect 37004 29096 37056 29102
rect 37004 29038 37056 29044
rect 35992 28756 36044 28762
rect 35992 28698 36044 28704
rect 37016 28626 37044 29038
rect 37004 28620 37056 28626
rect 37004 28562 37056 28568
rect 36452 28552 36504 28558
rect 36452 28494 36504 28500
rect 35992 28416 36044 28422
rect 35912 28364 35992 28370
rect 35912 28358 36044 28364
rect 35912 28342 36032 28358
rect 35624 27464 35676 27470
rect 35624 27406 35676 27412
rect 35808 27464 35860 27470
rect 35808 27406 35860 27412
rect 35532 26852 35584 26858
rect 35532 26794 35584 26800
rect 35532 24064 35584 24070
rect 35532 24006 35584 24012
rect 35544 23798 35572 24006
rect 35532 23792 35584 23798
rect 35532 23734 35584 23740
rect 35636 23610 35664 27406
rect 35912 26994 35940 28342
rect 36464 28082 36492 28494
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 36268 27872 36320 27878
rect 36268 27814 36320 27820
rect 36280 27606 36308 27814
rect 36268 27600 36320 27606
rect 36268 27542 36320 27548
rect 36268 27396 36320 27402
rect 36268 27338 36320 27344
rect 35900 26988 35952 26994
rect 35900 26930 35952 26936
rect 35912 25906 35940 26930
rect 36280 26926 36308 27338
rect 36268 26920 36320 26926
rect 36268 26862 36320 26868
rect 35900 25900 35952 25906
rect 35900 25842 35952 25848
rect 36280 24818 36308 26862
rect 36084 24812 36136 24818
rect 36084 24754 36136 24760
rect 36268 24812 36320 24818
rect 36268 24754 36320 24760
rect 35900 24676 35952 24682
rect 35900 24618 35952 24624
rect 35716 24608 35768 24614
rect 35716 24550 35768 24556
rect 35728 24206 35756 24550
rect 35716 24200 35768 24206
rect 35716 24142 35768 24148
rect 35544 23582 35664 23610
rect 35440 20460 35492 20466
rect 35440 20402 35492 20408
rect 35544 20210 35572 23582
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 35636 23118 35664 23462
rect 35624 23112 35676 23118
rect 35624 23054 35676 23060
rect 35912 22778 35940 24618
rect 36096 24138 36124 24754
rect 36176 24336 36228 24342
rect 36176 24278 36228 24284
rect 36084 24132 36136 24138
rect 36084 24074 36136 24080
rect 35900 22772 35952 22778
rect 35900 22714 35952 22720
rect 36188 22166 36216 24278
rect 36280 24206 36308 24754
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 36820 24200 36872 24206
rect 36820 24142 36872 24148
rect 36728 23588 36780 23594
rect 36728 23530 36780 23536
rect 36176 22160 36228 22166
rect 36176 22102 36228 22108
rect 35716 21888 35768 21894
rect 35716 21830 35768 21836
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35452 20182 35572 20210
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35348 19780 35400 19786
rect 35348 19722 35400 19728
rect 35360 19514 35388 19722
rect 35348 19508 35400 19514
rect 35348 19450 35400 19456
rect 35452 19394 35480 20182
rect 35636 19990 35664 21286
rect 35728 20398 35756 21830
rect 36188 21622 36216 22102
rect 36360 22024 36412 22030
rect 36360 21966 36412 21972
rect 36268 21956 36320 21962
rect 36268 21898 36320 21904
rect 36176 21616 36228 21622
rect 36176 21558 36228 21564
rect 36280 21554 36308 21898
rect 36372 21690 36400 21966
rect 36740 21962 36768 23530
rect 36832 23322 36860 24142
rect 37016 24138 37044 28562
rect 37384 28558 37412 29106
rect 37372 28552 37424 28558
rect 37372 28494 37424 28500
rect 37372 24608 37424 24614
rect 37372 24550 37424 24556
rect 37004 24132 37056 24138
rect 37004 24074 37056 24080
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 36820 23316 36872 23322
rect 36820 23258 36872 23264
rect 36832 22030 36860 23258
rect 37188 22636 37240 22642
rect 37188 22578 37240 22584
rect 37200 22522 37228 22578
rect 37292 22522 37320 24006
rect 37384 23866 37412 24550
rect 37372 23860 37424 23866
rect 37372 23802 37424 23808
rect 37200 22494 37320 22522
rect 37292 22094 37320 22494
rect 37292 22066 37412 22094
rect 36820 22024 36872 22030
rect 36820 21966 36872 21972
rect 36728 21956 36780 21962
rect 36728 21898 36780 21904
rect 37384 21894 37412 22066
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 36360 21684 36412 21690
rect 36360 21626 36412 21632
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36084 20528 36136 20534
rect 36084 20470 36136 20476
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35624 19984 35676 19990
rect 35624 19926 35676 19932
rect 35716 19848 35768 19854
rect 35912 19836 35940 20198
rect 36096 19854 36124 20470
rect 36360 20392 36412 20398
rect 36360 20334 36412 20340
rect 36372 19854 36400 20334
rect 35768 19808 35940 19836
rect 35716 19790 35768 19796
rect 35716 19712 35768 19718
rect 35716 19654 35768 19660
rect 35532 19508 35584 19514
rect 35532 19450 35584 19456
rect 35360 19366 35480 19394
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35360 18290 35388 19366
rect 35440 19304 35492 19310
rect 35440 19246 35492 19252
rect 35452 18970 35480 19246
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 34808 18142 35480 18170
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 34624 15570 34652 15846
rect 34716 15586 34744 17138
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34808 15706 34836 17070
rect 35360 17066 35388 18022
rect 35348 17060 35400 17066
rect 35348 17002 35400 17008
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 34612 15564 34664 15570
rect 34716 15558 34836 15586
rect 34612 15506 34664 15512
rect 34624 15162 34652 15506
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34612 15156 34664 15162
rect 34612 15098 34664 15104
rect 34716 14618 34744 15438
rect 34704 14612 34756 14618
rect 34704 14554 34756 14560
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 34060 14000 34112 14006
rect 34060 13942 34112 13948
rect 34716 13326 34744 14554
rect 34808 14074 34836 15558
rect 35452 15450 35480 18142
rect 35544 17134 35572 19450
rect 35728 19378 35756 19654
rect 35716 19372 35768 19378
rect 35716 19314 35768 19320
rect 35624 18760 35676 18766
rect 35624 18702 35676 18708
rect 35636 18358 35664 18702
rect 35624 18352 35676 18358
rect 35624 18294 35676 18300
rect 35532 17128 35584 17134
rect 35532 17070 35584 17076
rect 35544 15570 35572 17070
rect 35636 16658 35664 18294
rect 35728 18290 35756 19314
rect 35808 18624 35860 18630
rect 35808 18566 35860 18572
rect 35716 18284 35768 18290
rect 35716 18226 35768 18232
rect 35820 18222 35848 18566
rect 35912 18426 35940 19808
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36360 19848 36412 19854
rect 36360 19790 36412 19796
rect 36096 19514 36124 19790
rect 36084 19508 36136 19514
rect 36084 19450 36136 19456
rect 36452 19440 36504 19446
rect 36452 19382 36504 19388
rect 36464 18766 36492 19382
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 35900 18420 35952 18426
rect 35900 18362 35952 18368
rect 36544 18284 36596 18290
rect 36544 18226 36596 18232
rect 37280 18284 37332 18290
rect 37280 18226 37332 18232
rect 35808 18216 35860 18222
rect 35808 18158 35860 18164
rect 35624 16652 35676 16658
rect 35624 16594 35676 16600
rect 35820 16454 35848 18158
rect 36556 17338 36584 18226
rect 37292 18086 37320 18226
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35912 16590 35940 16934
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 35808 16448 35860 16454
rect 35808 16390 35860 16396
rect 35820 16182 35848 16390
rect 35808 16176 35860 16182
rect 35808 16118 35860 16124
rect 35532 15564 35584 15570
rect 35532 15506 35584 15512
rect 35452 15422 35664 15450
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 35532 14408 35584 14414
rect 35532 14350 35584 14356
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 34704 13320 34756 13326
rect 34704 13262 34756 13268
rect 33428 12238 33456 13262
rect 34428 13252 34480 13258
rect 34428 13194 34480 13200
rect 34440 12782 34468 13194
rect 34808 12986 34836 14010
rect 35544 13870 35572 14350
rect 35440 13864 35492 13870
rect 35440 13806 35492 13812
rect 35532 13864 35584 13870
rect 35532 13806 35584 13812
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 35256 13184 35308 13190
rect 35256 13126 35308 13132
rect 34796 12980 34848 12986
rect 34796 12922 34848 12928
rect 35268 12850 35296 13126
rect 35452 12850 35480 13806
rect 35256 12844 35308 12850
rect 35256 12786 35308 12792
rect 35440 12844 35492 12850
rect 35440 12786 35492 12792
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 34428 12776 34480 12782
rect 34428 12718 34480 12724
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33428 11898 33456 12174
rect 33520 12170 33548 12718
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35452 12442 35480 12786
rect 35440 12436 35492 12442
rect 35440 12378 35492 12384
rect 33508 12164 33560 12170
rect 33508 12106 33560 12112
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33520 11694 33548 12106
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 33704 11830 33732 12038
rect 34428 11892 34480 11898
rect 34428 11834 34480 11840
rect 33692 11824 33744 11830
rect 33692 11766 33744 11772
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 34440 11354 34468 11834
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34428 11348 34480 11354
rect 34428 11290 34480 11296
rect 34888 11144 34940 11150
rect 34888 11086 34940 11092
rect 34152 11076 34204 11082
rect 34152 11018 34204 11024
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 33244 9518 33272 10746
rect 33232 9512 33284 9518
rect 33232 9454 33284 9460
rect 32680 9036 32732 9042
rect 32680 8978 32732 8984
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 30748 7404 30800 7410
rect 30748 7346 30800 7352
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 30760 7002 30788 7346
rect 30944 7206 30972 7346
rect 32692 7342 32720 8978
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 32680 7336 32732 7342
rect 32680 7278 32732 7284
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 33048 7200 33100 7206
rect 33048 7142 33100 7148
rect 30748 6996 30800 7002
rect 30748 6938 30800 6944
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 33060 6798 33088 7142
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 33048 6792 33100 6798
rect 33048 6734 33100 6740
rect 30392 5846 30420 6734
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 33048 6248 33100 6254
rect 33048 6190 33100 6196
rect 32864 5908 32916 5914
rect 32864 5850 32916 5856
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30116 5166 30144 5646
rect 30392 5166 30420 5782
rect 32220 5568 32272 5574
rect 32220 5510 32272 5516
rect 30840 5364 30892 5370
rect 30840 5306 30892 5312
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 29736 5024 29788 5030
rect 29736 4966 29788 4972
rect 29748 4622 29776 4966
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 28448 4616 28500 4622
rect 28448 4558 28500 4564
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 27632 4282 27660 4558
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 29736 4480 29788 4486
rect 29736 4422 29788 4428
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 28368 4214 28396 4422
rect 28356 4208 28408 4214
rect 28356 4150 28408 4156
rect 29748 4146 29776 4422
rect 30852 4282 30880 5306
rect 31944 5228 31996 5234
rect 31944 5170 31996 5176
rect 31956 4554 31984 5170
rect 32232 4622 32260 5510
rect 32876 4622 32904 5850
rect 33060 5658 33088 6190
rect 33152 5846 33180 6258
rect 33704 6186 33732 8366
rect 34060 7404 34112 7410
rect 34060 7346 34112 7352
rect 34072 6866 34100 7346
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 33876 6724 33928 6730
rect 33876 6666 33928 6672
rect 33888 6254 33916 6666
rect 34072 6662 34100 6802
rect 34164 6798 34192 11018
rect 34900 10810 34928 11086
rect 34888 10804 34940 10810
rect 34888 10746 34940 10752
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34624 8974 34652 9318
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34440 8430 34468 8842
rect 34428 8424 34480 8430
rect 34428 8366 34480 8372
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 34348 7410 34376 8298
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34348 7002 34376 7346
rect 34520 7200 34572 7206
rect 34520 7142 34572 7148
rect 34336 6996 34388 7002
rect 34336 6938 34388 6944
rect 34532 6934 34560 7142
rect 34520 6928 34572 6934
rect 34520 6870 34572 6876
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 33876 6248 33928 6254
rect 33876 6190 33928 6196
rect 33968 6248 34020 6254
rect 33968 6190 34020 6196
rect 33692 6180 33744 6186
rect 33692 6122 33744 6128
rect 33140 5840 33192 5846
rect 33140 5782 33192 5788
rect 33140 5704 33192 5710
rect 33060 5652 33140 5658
rect 33060 5646 33192 5652
rect 33232 5704 33284 5710
rect 33232 5646 33284 5652
rect 33060 5630 33180 5646
rect 33152 5166 33180 5630
rect 33244 5370 33272 5646
rect 33324 5568 33376 5574
rect 33324 5510 33376 5516
rect 33232 5364 33284 5370
rect 33232 5306 33284 5312
rect 33336 5234 33364 5510
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33140 5160 33192 5166
rect 33140 5102 33192 5108
rect 32220 4616 32272 4622
rect 32220 4558 32272 4564
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 31944 4548 31996 4554
rect 31944 4490 31996 4496
rect 30840 4276 30892 4282
rect 30840 4218 30892 4224
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29460 4072 29512 4078
rect 29460 4014 29512 4020
rect 29472 3738 29500 4014
rect 31956 3738 31984 4490
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 29460 3732 29512 3738
rect 29460 3674 29512 3680
rect 31944 3732 31996 3738
rect 31944 3674 31996 3680
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 24872 3194 24900 3674
rect 32140 3466 32168 4422
rect 32876 4282 32904 4558
rect 33336 4554 33364 5170
rect 33704 5098 33732 6122
rect 33876 6112 33928 6118
rect 33876 6054 33928 6060
rect 33888 5778 33916 6054
rect 33876 5772 33928 5778
rect 33876 5714 33928 5720
rect 33980 5370 34008 6190
rect 34072 6118 34100 6598
rect 34164 6322 34192 6734
rect 34152 6316 34204 6322
rect 34152 6258 34204 6264
rect 34060 6112 34112 6118
rect 34060 6054 34112 6060
rect 33968 5364 34020 5370
rect 33968 5306 34020 5312
rect 34532 5302 34560 6870
rect 34624 6866 34652 8910
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34624 5914 34652 6802
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34716 6390 34744 6598
rect 34704 6384 34756 6390
rect 34704 6326 34756 6332
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34520 5296 34572 5302
rect 34520 5238 34572 5244
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 33692 5092 33744 5098
rect 33692 5034 33744 5040
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 33428 4622 33456 4966
rect 34164 4826 34192 5170
rect 34152 4820 34204 4826
rect 34152 4762 34204 4768
rect 34808 4758 34836 10542
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 35360 9518 35388 12038
rect 35440 9580 35492 9586
rect 35440 9522 35492 9528
rect 35348 9512 35400 9518
rect 35348 9454 35400 9460
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 35452 9178 35480 9522
rect 35440 9172 35492 9178
rect 35440 9114 35492 9120
rect 35348 9036 35400 9042
rect 35348 8978 35400 8984
rect 34888 8968 34940 8974
rect 34888 8910 34940 8916
rect 34900 8634 34928 8910
rect 34888 8628 34940 8634
rect 34888 8570 34940 8576
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35164 6928 35216 6934
rect 35164 6870 35216 6876
rect 35176 6798 35204 6870
rect 35360 6798 35388 8978
rect 35544 8838 35572 13806
rect 35636 12434 35664 15422
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36464 15162 36492 15370
rect 36452 15156 36504 15162
rect 36452 15098 36504 15104
rect 36084 12640 36136 12646
rect 36084 12582 36136 12588
rect 35808 12436 35860 12442
rect 35636 12406 35756 12434
rect 35728 10606 35756 12406
rect 35808 12378 35860 12384
rect 35820 11082 35848 12378
rect 36096 12238 36124 12582
rect 36084 12232 36136 12238
rect 36084 12174 36136 12180
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 35808 11076 35860 11082
rect 35808 11018 35860 11024
rect 35820 10674 35848 11018
rect 35912 10742 35940 11086
rect 35900 10736 35952 10742
rect 35900 10678 35952 10684
rect 35808 10668 35860 10674
rect 35808 10610 35860 10616
rect 35716 10600 35768 10606
rect 35716 10542 35768 10548
rect 35912 9330 35940 10678
rect 35992 9376 36044 9382
rect 35912 9324 35992 9330
rect 35912 9318 36044 9324
rect 35912 9302 36032 9318
rect 35912 8974 35940 9302
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 35532 8832 35584 8838
rect 35532 8774 35584 8780
rect 35912 8498 35940 8910
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35164 6792 35216 6798
rect 35164 6734 35216 6740
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 34888 6724 34940 6730
rect 34888 6666 34940 6672
rect 34900 6458 34928 6666
rect 34888 6452 34940 6458
rect 34888 6394 34940 6400
rect 35820 6322 35848 6802
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 37292 5273 37320 18022
rect 37384 15706 37412 21830
rect 37660 20058 37688 37062
rect 38108 33992 38160 33998
rect 38106 33960 38108 33969
rect 38160 33960 38162 33969
rect 38106 33895 38162 33904
rect 38108 30048 38160 30054
rect 38108 29990 38160 29996
rect 38120 29889 38148 29990
rect 38106 29880 38162 29889
rect 38106 29815 38162 29824
rect 38016 26512 38068 26518
rect 38016 26454 38068 26460
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 37648 20052 37700 20058
rect 37648 19994 37700 20000
rect 37660 19854 37688 19994
rect 37648 19848 37700 19854
rect 37648 19790 37700 19796
rect 37660 18970 37688 19790
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37844 18426 37872 26318
rect 38028 25945 38056 26454
rect 38014 25936 38070 25945
rect 38014 25871 38070 25880
rect 38014 21992 38070 22001
rect 38014 21927 38070 21936
rect 38028 21894 38056 21927
rect 38016 21888 38068 21894
rect 38016 21830 38068 21836
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 38016 18080 38068 18086
rect 38016 18022 38068 18028
rect 38028 17921 38056 18022
rect 38014 17912 38070 17921
rect 38014 17847 38070 17856
rect 37372 15700 37424 15706
rect 37372 15642 37424 15648
rect 38016 14340 38068 14346
rect 38016 14282 38068 14288
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 37832 8356 37884 8362
rect 37832 8298 37884 8304
rect 37740 6656 37792 6662
rect 37740 6598 37792 6604
rect 37752 5642 37780 6598
rect 37844 6322 37872 8298
rect 37936 7274 37964 14214
rect 38028 13977 38056 14282
rect 38014 13968 38070 13977
rect 38014 13903 38070 13912
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38120 9897 38148 9998
rect 38106 9888 38162 9897
rect 38106 9823 38162 9832
rect 37924 7268 37976 7274
rect 37924 7210 37976 7216
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 38016 6112 38068 6118
rect 38016 6054 38068 6060
rect 38028 5953 38056 6054
rect 38014 5944 38070 5953
rect 38014 5879 38070 5888
rect 37740 5636 37792 5642
rect 37740 5578 37792 5584
rect 37278 5264 37334 5273
rect 37278 5199 37334 5208
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34796 4752 34848 4758
rect 34796 4694 34848 4700
rect 33416 4616 33468 4622
rect 33416 4558 33468 4564
rect 33324 4548 33376 4554
rect 33324 4490 33376 4496
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 32876 3534 32904 4218
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 32128 3460 32180 3466
rect 32128 3402 32180 3408
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 37752 2446 37780 5578
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 1601 1900 2314
rect 2792 2281 2820 2382
rect 2778 2272 2834 2281
rect 2778 2207 2834 2216
rect 1858 1592 1914 1601
rect 1858 1527 1914 1536
rect 3988 921 4016 2382
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 38028 2009 38056 2246
rect 38014 2000 38070 2009
rect 38014 1935 38070 1944
rect 3974 912 4030 921
rect 3974 847 4030 856
rect 1398 368 1454 377
rect 1398 303 1454 312
<< via2 >>
rect 3330 39616 3386 39672
rect 3238 38936 3294 38992
rect 3422 38256 3478 38312
rect 4066 37576 4122 37632
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3974 36896 4030 36952
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4066 36236 4122 36272
rect 4066 36216 4068 36236
rect 4068 36216 4120 36236
rect 4120 36216 4122 36236
rect 3422 35536 3478 35592
rect 3146 34856 3202 34912
rect 2870 34176 2926 34232
rect 1398 33532 1400 33552
rect 1400 33532 1452 33552
rect 1452 33532 1454 33552
rect 1398 33496 1454 33532
rect 1398 32136 1454 32192
rect 3238 31456 3294 31512
rect 1398 30812 1400 30832
rect 1400 30812 1452 30832
rect 1452 30812 1454 30832
rect 1398 30776 1454 30812
rect 1398 29416 1454 29472
rect 1398 28056 1454 28112
rect 1398 26696 1454 26752
rect 1398 25336 1454 25392
rect 1398 23976 1454 24032
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4618 32816 4674 32872
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 3882 30096 3938 30152
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 3790 28736 3846 28792
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27376 4122 27432
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 1398 22616 1454 22672
rect 1398 21256 1454 21312
rect 1398 19896 1454 19952
rect 3422 24656 3478 24712
rect 1398 18536 1454 18592
rect 1398 17176 1454 17232
rect 1398 15816 1454 15872
rect 1398 14456 1454 14512
rect 1398 13096 1454 13152
rect 1398 11736 1454 11792
rect 1398 10376 1454 10432
rect 1398 9052 1400 9072
rect 1400 9052 1452 9072
rect 1452 9052 1454 9072
rect 1398 9016 1454 9052
rect 1398 7656 1454 7712
rect 1398 6296 1454 6352
rect 1398 4936 1454 4992
rect 1398 3576 1454 3632
rect 3606 23296 3662 23352
rect 3422 21936 3478 21992
rect 3514 19216 3570 19272
rect 3422 17856 3478 17912
rect 3422 16496 3478 16552
rect 3422 15136 3478 15192
rect 3422 13776 3478 13832
rect 3238 12416 3294 12472
rect 3422 11056 3478 11112
rect 3422 9716 3478 9752
rect 3422 9696 3424 9716
rect 3424 9696 3476 9716
rect 3476 9696 3478 9716
rect 3422 8336 3478 8392
rect 3422 6976 3478 7032
rect 4526 26016 4582 26072
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 3974 20576 4030 20632
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3422 5616 3478 5672
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3422 2896 3478 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 9678 20304 9734 20360
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 38014 37848 38070 37904
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 14186 5072 14242 5128
rect 17222 5228 17278 5264
rect 17222 5208 17224 5228
rect 17224 5208 17276 5228
rect 17276 5208 17278 5228
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 21914 20324 21970 20360
rect 21914 20304 21916 20324
rect 21916 20304 21968 20324
rect 21968 20304 21970 20324
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 25686 9696 25742 9752
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 25962 5228 26018 5264
rect 25962 5208 25964 5228
rect 25964 5208 26016 5228
rect 26016 5208 26018 5228
rect 27250 5072 27306 5128
rect 28998 9560 29054 9616
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 29550 9580 29606 9616
rect 29550 9560 29552 9580
rect 29552 9560 29604 9580
rect 29604 9560 29606 9580
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 38106 33940 38108 33960
rect 38108 33940 38160 33960
rect 38160 33940 38162 33960
rect 38106 33904 38162 33940
rect 38106 29824 38162 29880
rect 38014 25880 38070 25936
rect 38014 21936 38070 21992
rect 38014 17856 38070 17912
rect 38014 13912 38070 13968
rect 38106 9832 38162 9888
rect 38014 5888 38070 5944
rect 37278 5208 37334 5264
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 2778 2216 2834 2272
rect 1858 1536 1914 1592
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38014 1944 38070 2000
rect 3974 856 4030 912
rect 1398 312 1454 368
<< metal3 >>
rect 0 39674 800 39704
rect 3325 39674 3391 39677
rect 0 39672 3391 39674
rect 0 39616 3330 39672
rect 3386 39616 3391 39672
rect 0 39614 3391 39616
rect 0 39584 800 39614
rect 3325 39611 3391 39614
rect 0 38994 800 39024
rect 3233 38994 3299 38997
rect 0 38992 3299 38994
rect 0 38936 3238 38992
rect 3294 38936 3299 38992
rect 0 38934 3299 38936
rect 0 38904 800 38934
rect 3233 38931 3299 38934
rect 0 38314 800 38344
rect 3417 38314 3483 38317
rect 0 38312 3483 38314
rect 0 38256 3422 38312
rect 3478 38256 3483 38312
rect 0 38254 3483 38256
rect 0 38224 800 38254
rect 3417 38251 3483 38254
rect 38009 37906 38075 37909
rect 39200 37906 40000 37936
rect 38009 37904 40000 37906
rect 38009 37848 38014 37904
rect 38070 37848 40000 37904
rect 38009 37846 40000 37848
rect 38009 37843 38075 37846
rect 39200 37816 40000 37846
rect 0 37634 800 37664
rect 4061 37634 4127 37637
rect 0 37632 4127 37634
rect 0 37576 4066 37632
rect 4122 37576 4127 37632
rect 0 37574 4127 37576
rect 0 37544 800 37574
rect 4061 37571 4127 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 0 36954 800 36984
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 3969 36954 4035 36957
rect 0 36952 4035 36954
rect 0 36896 3974 36952
rect 4030 36896 4035 36952
rect 0 36894 4035 36896
rect 0 36864 800 36894
rect 3969 36891 4035 36894
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36274 800 36304
rect 4061 36274 4127 36277
rect 0 36272 4127 36274
rect 0 36216 4066 36272
rect 4122 36216 4127 36272
rect 0 36214 4127 36216
rect 0 36184 800 36214
rect 4061 36211 4127 36214
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35594 800 35624
rect 3417 35594 3483 35597
rect 0 35592 3483 35594
rect 0 35536 3422 35592
rect 3478 35536 3483 35592
rect 0 35534 3483 35536
rect 0 35504 800 35534
rect 3417 35531 3483 35534
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34914 800 34944
rect 3141 34914 3207 34917
rect 0 34912 3207 34914
rect 0 34856 3146 34912
rect 3202 34856 3207 34912
rect 0 34854 3207 34856
rect 0 34824 800 34854
rect 3141 34851 3207 34854
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 0 34234 800 34264
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 2865 34234 2931 34237
rect 0 34232 2931 34234
rect 0 34176 2870 34232
rect 2926 34176 2931 34232
rect 0 34174 2931 34176
rect 0 34144 800 34174
rect 2865 34171 2931 34174
rect 38101 33962 38167 33965
rect 39200 33962 40000 33992
rect 38101 33960 40000 33962
rect 38101 33904 38106 33960
rect 38162 33904 40000 33960
rect 38101 33902 40000 33904
rect 38101 33899 38167 33902
rect 39200 33872 40000 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33554 800 33584
rect 1393 33554 1459 33557
rect 0 33552 1459 33554
rect 0 33496 1398 33552
rect 1454 33496 1459 33552
rect 0 33494 1459 33496
rect 0 33464 800 33494
rect 1393 33491 1459 33494
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32874 800 32904
rect 4613 32874 4679 32877
rect 0 32872 4679 32874
rect 0 32816 4618 32872
rect 4674 32816 4679 32872
rect 0 32814 4679 32816
rect 0 32784 800 32814
rect 4613 32811 4679 32814
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 0 32194 800 32224
rect 1393 32194 1459 32197
rect 0 32192 1459 32194
rect 0 32136 1398 32192
rect 1454 32136 1459 32192
rect 0 32134 1459 32136
rect 0 32104 800 32134
rect 1393 32131 1459 32134
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 0 31514 800 31544
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 3233 31514 3299 31517
rect 0 31512 3299 31514
rect 0 31456 3238 31512
rect 3294 31456 3299 31512
rect 0 31454 3299 31456
rect 0 31424 800 31454
rect 3233 31451 3299 31454
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30834 800 30864
rect 1393 30834 1459 30837
rect 0 30832 1459 30834
rect 0 30776 1398 30832
rect 1454 30776 1459 30832
rect 0 30774 1459 30776
rect 0 30744 800 30774
rect 1393 30771 1459 30774
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 30154 800 30184
rect 3877 30154 3943 30157
rect 0 30152 3943 30154
rect 0 30096 3882 30152
rect 3938 30096 3943 30152
rect 0 30094 3943 30096
rect 0 30064 800 30094
rect 3877 30091 3943 30094
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 38101 29882 38167 29885
rect 39200 29882 40000 29912
rect 38101 29880 40000 29882
rect 38101 29824 38106 29880
rect 38162 29824 40000 29880
rect 38101 29822 40000 29824
rect 38101 29819 38167 29822
rect 39200 29792 40000 29822
rect 0 29474 800 29504
rect 1393 29474 1459 29477
rect 0 29472 1459 29474
rect 0 29416 1398 29472
rect 1454 29416 1459 29472
rect 0 29414 1459 29416
rect 0 29384 800 29414
rect 1393 29411 1459 29414
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 3785 28794 3851 28797
rect 0 28792 3851 28794
rect 0 28736 3790 28792
rect 3846 28736 3851 28792
rect 0 28734 3851 28736
rect 0 28704 800 28734
rect 3785 28731 3851 28734
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 28114 800 28144
rect 1393 28114 1459 28117
rect 0 28112 1459 28114
rect 0 28056 1398 28112
rect 1454 28056 1459 28112
rect 0 28054 1459 28056
rect 0 28024 800 28054
rect 1393 28051 1459 28054
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27434 800 27464
rect 4061 27434 4127 27437
rect 0 27432 4127 27434
rect 0 27376 4066 27432
rect 4122 27376 4127 27432
rect 0 27374 4127 27376
rect 0 27344 800 27374
rect 4061 27371 4127 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 0 26754 800 26784
rect 1393 26754 1459 26757
rect 0 26752 1459 26754
rect 0 26696 1398 26752
rect 1454 26696 1459 26752
rect 0 26694 1459 26696
rect 0 26664 800 26694
rect 1393 26691 1459 26694
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 0 26074 800 26104
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 4521 26074 4587 26077
rect 0 26072 4587 26074
rect 0 26016 4526 26072
rect 4582 26016 4587 26072
rect 0 26014 4587 26016
rect 0 25984 800 26014
rect 4521 26011 4587 26014
rect 38009 25938 38075 25941
rect 39200 25938 40000 25968
rect 38009 25936 40000 25938
rect 38009 25880 38014 25936
rect 38070 25880 40000 25936
rect 38009 25878 40000 25880
rect 38009 25875 38075 25878
rect 39200 25848 40000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25394 800 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 800 25334
rect 1393 25331 1459 25334
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24714 800 24744
rect 3417 24714 3483 24717
rect 0 24712 3483 24714
rect 0 24656 3422 24712
rect 3478 24656 3483 24712
rect 0 24654 3483 24656
rect 0 24624 800 24654
rect 3417 24651 3483 24654
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 0 24034 800 24064
rect 1393 24034 1459 24037
rect 0 24032 1459 24034
rect 0 23976 1398 24032
rect 1454 23976 1459 24032
rect 0 23974 1459 23976
rect 0 23944 800 23974
rect 1393 23971 1459 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 4208 23424 4528 23425
rect 0 23354 800 23384
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 3601 23354 3667 23357
rect 0 23352 3667 23354
rect 0 23296 3606 23352
rect 3662 23296 3667 23352
rect 0 23294 3667 23296
rect 0 23264 800 23294
rect 3601 23291 3667 23294
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22674 800 22704
rect 1393 22674 1459 22677
rect 0 22672 1459 22674
rect 0 22616 1398 22672
rect 1454 22616 1459 22672
rect 0 22614 1459 22616
rect 0 22584 800 22614
rect 1393 22611 1459 22614
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21994 800 22024
rect 3417 21994 3483 21997
rect 0 21992 3483 21994
rect 0 21936 3422 21992
rect 3478 21936 3483 21992
rect 0 21934 3483 21936
rect 0 21904 800 21934
rect 3417 21931 3483 21934
rect 38009 21994 38075 21997
rect 39200 21994 40000 22024
rect 38009 21992 40000 21994
rect 38009 21936 38014 21992
rect 38070 21936 40000 21992
rect 38009 21934 40000 21936
rect 38009 21931 38075 21934
rect 39200 21904 40000 21934
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 0 21314 800 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 800 21254
rect 1393 21251 1459 21254
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 0 20634 800 20664
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 3969 20634 4035 20637
rect 0 20632 4035 20634
rect 0 20576 3974 20632
rect 4030 20576 4035 20632
rect 0 20574 4035 20576
rect 0 20544 800 20574
rect 3969 20571 4035 20574
rect 9673 20362 9739 20365
rect 21909 20362 21975 20365
rect 9673 20360 21975 20362
rect 9673 20304 9678 20360
rect 9734 20304 21914 20360
rect 21970 20304 21975 20360
rect 9673 20302 21975 20304
rect 9673 20299 9739 20302
rect 21909 20299 21975 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19954 800 19984
rect 1393 19954 1459 19957
rect 0 19952 1459 19954
rect 0 19896 1398 19952
rect 1454 19896 1459 19952
rect 0 19894 1459 19896
rect 0 19864 800 19894
rect 1393 19891 1459 19894
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19274 800 19304
rect 3509 19274 3575 19277
rect 0 19272 3575 19274
rect 0 19216 3514 19272
rect 3570 19216 3575 19272
rect 0 19214 3575 19216
rect 0 19184 800 19214
rect 3509 19211 3575 19214
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 0 18594 800 18624
rect 1393 18594 1459 18597
rect 0 18592 1459 18594
rect 0 18536 1398 18592
rect 1454 18536 1459 18592
rect 0 18534 1459 18536
rect 0 18504 800 18534
rect 1393 18531 1459 18534
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4208 17984 4528 17985
rect 0 17914 800 17944
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 3417 17914 3483 17917
rect 0 17912 3483 17914
rect 0 17856 3422 17912
rect 3478 17856 3483 17912
rect 0 17854 3483 17856
rect 0 17824 800 17854
rect 3417 17851 3483 17854
rect 38009 17914 38075 17917
rect 39200 17914 40000 17944
rect 38009 17912 40000 17914
rect 38009 17856 38014 17912
rect 38070 17856 40000 17912
rect 38009 17854 40000 17856
rect 38009 17851 38075 17854
rect 39200 17824 40000 17854
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17234 800 17264
rect 1393 17234 1459 17237
rect 0 17232 1459 17234
rect 0 17176 1398 17232
rect 1454 17176 1459 17232
rect 0 17174 1459 17176
rect 0 17144 800 17174
rect 1393 17171 1459 17174
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16554 800 16584
rect 3417 16554 3483 16557
rect 0 16552 3483 16554
rect 0 16496 3422 16552
rect 3478 16496 3483 16552
rect 0 16494 3483 16496
rect 0 16464 800 16494
rect 3417 16491 3483 16494
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 0 15874 800 15904
rect 1393 15874 1459 15877
rect 0 15872 1459 15874
rect 0 15816 1398 15872
rect 1454 15816 1459 15872
rect 0 15814 1459 15816
rect 0 15784 800 15814
rect 1393 15811 1459 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 0 15194 800 15224
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 3417 15194 3483 15197
rect 0 15192 3483 15194
rect 0 15136 3422 15192
rect 3478 15136 3483 15192
rect 0 15134 3483 15136
rect 0 15104 800 15134
rect 3417 15131 3483 15134
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 38009 13970 38075 13973
rect 39200 13970 40000 14000
rect 38009 13968 40000 13970
rect 38009 13912 38014 13968
rect 38070 13912 40000 13968
rect 38009 13910 40000 13912
rect 38009 13907 38075 13910
rect 39200 13880 40000 13910
rect 0 13834 800 13864
rect 3417 13834 3483 13837
rect 0 13832 3483 13834
rect 0 13776 3422 13832
rect 3478 13776 3483 13832
rect 0 13774 3483 13776
rect 0 13744 800 13774
rect 3417 13771 3483 13774
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4208 12544 4528 12545
rect 0 12474 800 12504
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 3233 12474 3299 12477
rect 0 12472 3299 12474
rect 0 12416 3238 12472
rect 3294 12416 3299 12472
rect 0 12414 3299 12416
rect 0 12384 800 12414
rect 3233 12411 3299 12414
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11794 800 11824
rect 1393 11794 1459 11797
rect 0 11792 1459 11794
rect 0 11736 1398 11792
rect 1454 11736 1459 11792
rect 0 11734 1459 11736
rect 0 11704 800 11734
rect 1393 11731 1459 11734
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 11114 800 11144
rect 3417 11114 3483 11117
rect 0 11112 3483 11114
rect 0 11056 3422 11112
rect 3478 11056 3483 11112
rect 0 11054 3483 11056
rect 0 11024 800 11054
rect 3417 11051 3483 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 38101 9890 38167 9893
rect 39200 9890 40000 9920
rect 38101 9888 40000 9890
rect 38101 9832 38106 9888
rect 38162 9832 40000 9888
rect 38101 9830 40000 9832
rect 38101 9827 38167 9830
rect 19568 9824 19888 9825
rect 0 9754 800 9784
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 39200 9800 40000 9830
rect 19568 9759 19888 9760
rect 3417 9754 3483 9757
rect 0 9752 3483 9754
rect 0 9696 3422 9752
rect 3478 9696 3483 9752
rect 0 9694 3483 9696
rect 0 9664 800 9694
rect 3417 9691 3483 9694
rect 25681 9754 25747 9757
rect 25681 9752 29010 9754
rect 25681 9696 25686 9752
rect 25742 9696 29010 9752
rect 25681 9694 29010 9696
rect 25681 9691 25747 9694
rect 28950 9621 29010 9694
rect 28950 9618 29059 9621
rect 29545 9618 29611 9621
rect 28950 9616 29611 9618
rect 28950 9560 28998 9616
rect 29054 9560 29550 9616
rect 29606 9560 29611 9616
rect 28950 9558 29611 9560
rect 28993 9555 29059 9558
rect 29545 9555 29611 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8394 800 8424
rect 3417 8394 3483 8397
rect 0 8392 3483 8394
rect 0 8336 3422 8392
rect 3478 8336 3483 8392
rect 0 8334 3483 8336
rect 0 8304 800 8334
rect 3417 8331 3483 8334
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 0 7714 800 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 4208 7104 4528 7105
rect 0 7034 800 7064
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 3417 7034 3483 7037
rect 0 7032 3483 7034
rect 0 6976 3422 7032
rect 3478 6976 3483 7032
rect 0 6974 3483 6976
rect 0 6944 800 6974
rect 3417 6971 3483 6974
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6354 800 6384
rect 1393 6354 1459 6357
rect 0 6352 1459 6354
rect 0 6296 1398 6352
rect 1454 6296 1459 6352
rect 0 6294 1459 6296
rect 0 6264 800 6294
rect 1393 6291 1459 6294
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 38009 5946 38075 5949
rect 39200 5946 40000 5976
rect 38009 5944 40000 5946
rect 38009 5888 38014 5944
rect 38070 5888 40000 5944
rect 38009 5886 40000 5888
rect 38009 5883 38075 5886
rect 39200 5856 40000 5886
rect 0 5674 800 5704
rect 3417 5674 3483 5677
rect 0 5672 3483 5674
rect 0 5616 3422 5672
rect 3478 5616 3483 5672
rect 0 5614 3483 5616
rect 0 5584 800 5614
rect 3417 5611 3483 5614
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 17217 5266 17283 5269
rect 6870 5264 17283 5266
rect 6870 5208 17222 5264
rect 17278 5208 17283 5264
rect 6870 5206 17283 5208
rect 0 4994 800 5024
rect 1393 4994 1459 4997
rect 0 4992 1459 4994
rect 0 4936 1398 4992
rect 1454 4936 1459 4992
rect 0 4934 1459 4936
rect 0 4904 800 4934
rect 1393 4931 1459 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 0 4314 800 4344
rect 6870 4314 6930 5206
rect 17217 5203 17283 5206
rect 25957 5266 26023 5269
rect 37273 5266 37339 5269
rect 25957 5264 37339 5266
rect 25957 5208 25962 5264
rect 26018 5208 37278 5264
rect 37334 5208 37339 5264
rect 25957 5206 37339 5208
rect 25957 5203 26023 5206
rect 37273 5203 37339 5206
rect 14181 5130 14247 5133
rect 27245 5130 27311 5133
rect 14181 5128 27311 5130
rect 14181 5072 14186 5128
rect 14242 5072 27250 5128
rect 27306 5072 27311 5128
rect 14181 5070 27311 5072
rect 14181 5067 14247 5070
rect 27245 5067 27311 5070
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4254 6930 4314
rect 0 4224 800 4254
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3634 800 3664
rect 1393 3634 1459 3637
rect 0 3632 1459 3634
rect 0 3576 1398 3632
rect 1454 3576 1459 3632
rect 0 3574 1459 3576
rect 0 3544 800 3574
rect 1393 3571 1459 3574
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2954 800 2984
rect 3417 2954 3483 2957
rect 0 2952 3483 2954
rect 0 2896 3422 2952
rect 3478 2896 3483 2952
rect 0 2894 3483 2896
rect 0 2864 800 2894
rect 3417 2891 3483 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 0 2274 800 2304
rect 2773 2274 2839 2277
rect 0 2272 2839 2274
rect 0 2216 2778 2272
rect 2834 2216 2839 2272
rect 0 2214 2839 2216
rect 0 2184 800 2214
rect 2773 2211 2839 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 38009 2002 38075 2005
rect 39200 2002 40000 2032
rect 38009 2000 40000 2002
rect 38009 1944 38014 2000
rect 38070 1944 40000 2000
rect 38009 1942 40000 1944
rect 38009 1939 38075 1942
rect 39200 1912 40000 1942
rect 0 1594 800 1624
rect 1853 1594 1919 1597
rect 0 1592 1919 1594
rect 0 1536 1858 1592
rect 1914 1536 1919 1592
rect 0 1534 1919 1536
rect 0 1504 800 1534
rect 1853 1531 1919 1534
rect 0 914 800 944
rect 3969 914 4035 917
rect 0 912 4035 914
rect 0 856 3974 912
rect 4030 856 4035 912
rect 0 854 4035 856
rect 0 824 800 854
rect 3969 851 4035 854
rect 0 370 800 400
rect 1393 370 1459 373
rect 0 368 1459 370
rect 0 312 1398 368
rect 1454 312 1459 368
rect 0 310 1459 312
rect 0 280 800 310
rect 1393 307 1459 310
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1644511149
transform 1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1644511149
transform -1 0 23460 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1644511149
transform -1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1644511149
transform 1 0 20148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__C
timestamp 1644511149
transform -1 0 22264 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__D
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A
timestamp 1644511149
transform 1 0 32292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__D
timestamp 1644511149
transform 1 0 21620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1644511149
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 1644511149
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__C
timestamp 1644511149
transform 1 0 17848 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__C
timestamp 1644511149
transform 1 0 16468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__D
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__C
timestamp 1644511149
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__D
timestamp 1644511149
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1644511149
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1644511149
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1644511149
transform 1 0 6164 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1644511149
transform -1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__C
timestamp 1644511149
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__D
timestamp 1644511149
transform -1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C
timestamp 1644511149
transform -1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1644511149
transform -1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1644511149
transform -1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1644511149
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1644511149
transform -1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A
timestamp 1644511149
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1644511149
transform 1 0 5704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1644511149
transform 1 0 5060 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1644511149
transform 1 0 5336 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1644511149
transform 1 0 5704 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1644511149
transform 1 0 6992 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1644511149
transform -1 0 7452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1644511149
transform 1 0 8004 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1644511149
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1644511149
transform -1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1644511149
transform -1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1644511149
transform 1 0 20976 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__C
timestamp 1644511149
transform 1 0 23920 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1644511149
transform -1 0 24932 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__C
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__C
timestamp 1644511149
transform 1 0 19780 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1644511149
transform 1 0 17572 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1644511149
transform 1 0 21160 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1644511149
transform -1 0 23736 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__C
timestamp 1644511149
transform 1 0 24656 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1644511149
transform -1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__D
timestamp 1644511149
transform -1 0 23920 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__D
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__D
timestamp 1644511149
transform 1 0 22540 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1644511149
transform 1 0 6808 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__D
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__D
timestamp 1644511149
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1644511149
transform -1 0 5244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1644511149
transform 1 0 8464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1644511149
transform -1 0 4784 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__D
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__D
timestamp 1644511149
transform 1 0 5612 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__D
timestamp 1644511149
transform 1 0 6256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__D
timestamp 1644511149
transform 1 0 20240 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__D
timestamp 1644511149
transform 1 0 20148 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__D
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__D
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__C
timestamp 1644511149
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__S
timestamp 1644511149
transform -1 0 34408 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1644511149
transform -1 0 35512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B
timestamp 1644511149
transform -1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__C
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A2
timestamp 1644511149
transform -1 0 34684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__C1
timestamp 1644511149
transform 1 0 34500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1644511149
transform 1 0 19320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__B
timestamp 1644511149
transform -1 0 20056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__C
timestamp 1644511149
transform -1 0 20148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1644511149
transform 1 0 31464 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B2
timestamp 1644511149
transform 1 0 31924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B1
timestamp 1644511149
transform -1 0 29072 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B2
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__B1
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__B2
timestamp 1644511149
transform -1 0 29716 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__B1
timestamp 1644511149
transform -1 0 30544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__B2
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B2
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__B2
timestamp 1644511149
transform -1 0 27600 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__B2
timestamp 1644511149
transform 1 0 28612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A0
timestamp 1644511149
transform 1 0 32660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__S
timestamp 1644511149
transform -1 0 33396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1644511149
transform -1 0 32936 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__S
timestamp 1644511149
transform -1 0 34224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1644511149
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B1
timestamp 1644511149
transform 1 0 33856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__C
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1644511149
transform 1 0 28336 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A0
timestamp 1644511149
transform -1 0 31372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A0
timestamp 1644511149
transform 1 0 29348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1644511149
transform 1 0 29808 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A0
timestamp 1644511149
transform -1 0 28980 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__S
timestamp 1644511149
transform 1 0 26404 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1644511149
transform -1 0 25668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A0
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A0
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A1
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A
timestamp 1644511149
transform 1 0 31464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A0
timestamp 1644511149
transform 1 0 26772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__S
timestamp 1644511149
transform 1 0 27324 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A
timestamp 1644511149
transform 1 0 28888 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A0
timestamp 1644511149
transform 1 0 28244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__S
timestamp 1644511149
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__A
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A0
timestamp 1644511149
transform 1 0 29440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1644511149
transform 1 0 29992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A
timestamp 1644511149
transform 1 0 33580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B1
timestamp 1644511149
transform -1 0 37444 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A
timestamp 1644511149
transform 1 0 34132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A
timestamp 1644511149
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1644511149
transform -1 0 34960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__C1
timestamp 1644511149
transform -1 0 35788 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1644511149
transform 1 0 33488 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1644511149
transform -1 0 33488 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__B1
timestamp 1644511149
transform 1 0 36064 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A3
timestamp 1644511149
transform 1 0 33580 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A
timestamp 1644511149
transform 1 0 33672 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A1
timestamp 1644511149
transform -1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B_N
timestamp 1644511149
transform -1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__C
timestamp 1644511149
transform -1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B2
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B2
timestamp 1644511149
transform 1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B2
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1644511149
transform -1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B2
timestamp 1644511149
transform 1 0 15088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A
timestamp 1644511149
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B2
timestamp 1644511149
transform -1 0 14260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A
timestamp 1644511149
transform 1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__B2
timestamp 1644511149
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1644511149
transform -1 0 10948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B2
timestamp 1644511149
transform -1 0 12696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1644511149
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B2
timestamp 1644511149
transform 1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A0
timestamp 1644511149
transform 1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A0
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A1
timestamp 1644511149
transform -1 0 24104 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1644511149
transform 1 0 25208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A
timestamp 1644511149
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B
timestamp 1644511149
transform 1 0 21712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__C
timestamp 1644511149
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__C1
timestamp 1644511149
transform 1 0 34500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A
timestamp 1644511149
transform 1 0 20516 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B
timestamp 1644511149
transform -1 0 20608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__C
timestamp 1644511149
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1644511149
transform 1 0 30452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__C1
timestamp 1644511149
transform -1 0 32660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1644511149
transform 1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B1
timestamp 1644511149
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1644511149
transform 1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1
timestamp 1644511149
transform 1 0 29992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A1
timestamp 1644511149
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B1
timestamp 1644511149
transform -1 0 27048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__C1
timestamp 1644511149
transform -1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1644511149
transform 1 0 29532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1644511149
transform 1 0 28888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A
timestamp 1644511149
transform 1 0 30176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A
timestamp 1644511149
transform -1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B
timestamp 1644511149
transform -1 0 20608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__C
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__B1
timestamp 1644511149
transform 1 0 33764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A
timestamp 1644511149
transform 1 0 31464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__CLK
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__CLK
timestamp 1644511149
transform 1 0 28796 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__CLK
timestamp 1644511149
transform 1 0 28888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 1644511149
transform 1 0 23644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__CLK
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 1644511149
transform 1 0 14168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__CLK
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__CLK
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 1644511149
transform -1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__CLK
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__CLK
timestamp 1644511149
transform -1 0 24564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__CLK
timestamp 1644511149
transform 1 0 35420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__CLK
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__CLK
timestamp 1644511149
transform -1 0 25300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__CLK
timestamp 1644511149
transform 1 0 28980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__CLK
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__CLK
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__CLK
timestamp 1644511149
transform 1 0 29716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__CLK
timestamp 1644511149
transform 1 0 30544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__CLK
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__CLK
timestamp 1644511149
transform 1 0 30084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__CLK
timestamp 1644511149
transform 1 0 34776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__CLK
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__CLK
timestamp 1644511149
transform 1 0 32568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__CLK
timestamp 1644511149
transform 1 0 31004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A
timestamp 1644511149
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1644511149
transform 1 0 21896 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 2208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 1564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 2208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 2208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 2208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 2208 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 2208 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 2208 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 2208 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 1564 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 2208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 1564 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 2208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 2208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 29992 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 37444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 37536 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1644511149
transform 1 0 37260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1644511149
transform -1 0 37444 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18
timestamp 1644511149
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_38 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_12
timestamp 1644511149
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_16 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_20
timestamp 1644511149
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_255
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_267
timestamp 1644511149
transform 1 0 25668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_58
timestamp 1644511149
transform 1 0 6440 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_107
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_119
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_143
timestamp 1644511149
transform 1 0 14260 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_155
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_167
timestamp 1644511149
transform 1 0 16468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_272
timestamp 1644511149
transform 1 0 26128 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_284
timestamp 1644511149
transform 1 0 27232 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_311
timestamp 1644511149
transform 1 0 29716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_317
timestamp 1644511149
transform 1 0 30268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_327
timestamp 1644511149
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_347
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1644511149
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_16
timestamp 1644511149
transform 1 0 2576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1644511149
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1644511149
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_115
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp 1644511149
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_158
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1644511149
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_195
timestamp 1644511149
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_241
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_247
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_268
timestamp 1644511149
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_287
timestamp 1644511149
transform 1 0 27508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1644511149
transform 1 0 29072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_324
timestamp 1644511149
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_341
timestamp 1644511149
transform 1 0 32476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_344
timestamp 1644511149
transform 1 0 32752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_356
timestamp 1644511149
transform 1 0 33856 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_368
timestamp 1644511149
transform 1 0 34960 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_380
timestamp 1644511149
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1644511149
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1644511149
transform 1 0 6808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_74
timestamp 1644511149
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1644511149
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1644511149
transform 1 0 9108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1644511149
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1644511149
transform 1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_113
timestamp 1644511149
transform 1 0 11500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_125
timestamp 1644511149
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1644511149
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1644511149
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1644511149
transform 1 0 18032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_213
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_222
timestamp 1644511149
transform 1 0 21528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1644511149
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1644511149
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_264
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_276
timestamp 1644511149
transform 1 0 26496 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_298
timestamp 1644511149
transform 1 0 28520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_312
timestamp 1644511149
transform 1 0 29808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_318
timestamp 1644511149
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_332
timestamp 1644511149
transform 1 0 31648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_339
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_343
timestamp 1644511149
transform 1 0 32660 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_12
timestamp 1644511149
transform 1 0 2208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1644511149
transform 1 0 2944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1644511149
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1644511149
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 1644511149
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1644511149
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_120
timestamp 1644511149
transform 1 0 12144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1644511149
transform 1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp 1644511149
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1644511149
transform 1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_155
timestamp 1644511149
transform 1 0 15364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1644511149
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1644511149
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_182
timestamp 1644511149
transform 1 0 17848 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_204
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_210
timestamp 1644511149
transform 1 0 20424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_248
timestamp 1644511149
transform 1 0 23920 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1644511149
transform 1 0 25484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_290
timestamp 1644511149
transform 1 0 27784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_302
timestamp 1644511149
transform 1 0 28888 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_311
timestamp 1644511149
transform 1 0 29716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_323
timestamp 1644511149
transform 1 0 30820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_343
timestamp 1644511149
transform 1 0 32660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_347
timestamp 1644511149
transform 1 0 33028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_355
timestamp 1644511149
transform 1 0 33764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_362
timestamp 1644511149
transform 1 0 34408 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_374
timestamp 1644511149
transform 1 0 35512 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_386
timestamp 1644511149
transform 1 0 36616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1644511149
transform 1 0 4416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_43
timestamp 1644511149
transform 1 0 5060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_55
timestamp 1644511149
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_67
timestamp 1644511149
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_106
timestamp 1644511149
transform 1 0 10856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_114
timestamp 1644511149
transform 1 0 11592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1644511149
transform 1 0 14352 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp 1644511149
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_166
timestamp 1644511149
transform 1 0 16376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1644511149
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1644511149
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_203
timestamp 1644511149
transform 1 0 19780 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_211
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_219
timestamp 1644511149
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_231
timestamp 1644511149
transform 1 0 22356 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_235
timestamp 1644511149
transform 1 0 22724 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_318
timestamp 1644511149
transform 1 0 30360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_330
timestamp 1644511149
transform 1 0 31464 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_342
timestamp 1644511149
transform 1 0 32568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_351
timestamp 1644511149
transform 1 0 33396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_367
timestamp 1644511149
transform 1 0 34868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_379
timestamp 1644511149
transform 1 0 35972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_391
timestamp 1644511149
transform 1 0 37076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1644511149
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1644511149
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1644511149
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1644511149
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1644511149
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp 1644511149
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1644511149
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_183
timestamp 1644511149
transform 1 0 17940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_191
timestamp 1644511149
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_198
timestamp 1644511149
transform 1 0 19320 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_210
timestamp 1644511149
transform 1 0 20424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_213
timestamp 1644511149
transform 1 0 20700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1644511149
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp 1644511149
transform 1 0 23644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_250
timestamp 1644511149
transform 1 0 24104 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_262
timestamp 1644511149
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1644511149
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_289
timestamp 1644511149
transform 1 0 27692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_301
timestamp 1644511149
transform 1 0 28796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_313
timestamp 1644511149
transform 1 0 29900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1644511149
transform 1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1644511149
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_345
timestamp 1644511149
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_359
timestamp 1644511149
transform 1 0 34132 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1644511149
transform 1 0 35972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1644511149
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_12
timestamp 1644511149
transform 1 0 2208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_35
timestamp 1644511149
transform 1 0 4324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_45
timestamp 1644511149
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_57
timestamp 1644511149
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_69
timestamp 1644511149
transform 1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1644511149
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_88
timestamp 1644511149
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp 1644511149
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_113
timestamp 1644511149
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_125
timestamp 1644511149
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1644511149
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1644511149
transform 1 0 14720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1644511149
transform 1 0 15272 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1644511149
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_218
timestamp 1644511149
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_230
timestamp 1644511149
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_236
timestamp 1644511149
transform 1 0 22816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1644511149
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_255
timestamp 1644511149
transform 1 0 24564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_267
timestamp 1644511149
transform 1 0 25668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_279
timestamp 1644511149
transform 1 0 26772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_291
timestamp 1644511149
transform 1 0 27876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1644511149
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_315
timestamp 1644511149
transform 1 0 30084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_319
timestamp 1644511149
transform 1 0 30452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_331
timestamp 1644511149
transform 1 0 31556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_343
timestamp 1644511149
transform 1 0 32660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_355
timestamp 1644511149
transform 1 0 33764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1644511149
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_379
timestamp 1644511149
transform 1 0 35972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_400
timestamp 1644511149
transform 1 0 37904 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1644511149
transform 1 0 38456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_28
timestamp 1644511149
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_59
timestamp 1644511149
transform 1 0 6532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_71
timestamp 1644511149
transform 1 0 7636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1644511149
transform 1 0 8280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_82
timestamp 1644511149
transform 1 0 8648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_85
timestamp 1644511149
transform 1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_91
timestamp 1644511149
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1644511149
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1644511149
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1644511149
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_143
timestamp 1644511149
transform 1 0 14260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_155
timestamp 1644511149
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_198
timestamp 1644511149
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_210
timestamp 1644511149
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1644511149
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_233
timestamp 1644511149
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1644511149
transform 1 0 23644 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_251
timestamp 1644511149
transform 1 0 24196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_263
timestamp 1644511149
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1644511149
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_313
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_316
timestamp 1644511149
transform 1 0 30176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1644511149
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_357
timestamp 1644511149
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_362
timestamp 1644511149
transform 1 0 34408 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_374
timestamp 1644511149
transform 1 0 35512 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_386
timestamp 1644511149
transform 1 0 36616 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_12
timestamp 1644511149
transform 1 0 2208 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_50
timestamp 1644511149
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_58
timestamp 1644511149
transform 1 0 6440 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1644511149
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_69
timestamp 1644511149
transform 1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1644511149
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_91
timestamp 1644511149
transform 1 0 9476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1644511149
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_107
timestamp 1644511149
transform 1 0 10948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_118
timestamp 1644511149
transform 1 0 11960 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1644511149
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1644511149
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1644511149
transform 1 0 14352 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1644511149
transform 1 0 15456 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_171
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_183
timestamp 1644511149
transform 1 0 17940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_217
timestamp 1644511149
transform 1 0 21068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_223
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_235
timestamp 1644511149
transform 1 0 22724 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_259
timestamp 1644511149
transform 1 0 24932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1644511149
transform 1 0 26864 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_292
timestamp 1644511149
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_23
timestamp 1644511149
transform 1 0 3220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_29
timestamp 1644511149
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1644511149
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1644511149
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_80
timestamp 1644511149
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1644511149
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_96
timestamp 1644511149
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1644511149
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1644511149
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_173
timestamp 1644511149
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_177
timestamp 1644511149
transform 1 0 17388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1644511149
transform 1 0 19596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1644511149
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_229
timestamp 1644511149
transform 1 0 22172 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_251
timestamp 1644511149
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_263
timestamp 1644511149
transform 1 0 25300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_301
timestamp 1644511149
transform 1 0 28796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_311
timestamp 1644511149
transform 1 0 29716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_323
timestamp 1644511149
transform 1 0 30820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_366
timestamp 1644511149
transform 1 0 34776 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_378
timestamp 1644511149
transform 1 0 35880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1644511149
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_396
timestamp 1644511149
transform 1 0 37536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_404
timestamp 1644511149
transform 1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_5
timestamp 1644511149
transform 1 0 1564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1644511149
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1644511149
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1644511149
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_49
timestamp 1644511149
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1644511149
transform 1 0 6716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1644511149
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1644511149
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_169
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_181
timestamp 1644511149
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1644511149
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_199
timestamp 1644511149
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_207
timestamp 1644511149
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_212
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1644511149
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1644511149
transform 1 0 27048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_294
timestamp 1644511149
transform 1 0 28152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_326
timestamp 1644511149
transform 1 0 31096 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_338
timestamp 1644511149
transform 1 0 32200 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_350
timestamp 1644511149
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1644511149
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_373
timestamp 1644511149
transform 1 0 35420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1644511149
transform 1 0 36524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_397
timestamp 1644511149
transform 1 0 37628 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1644511149
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_6
timestamp 1644511149
transform 1 0 1656 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_36
timestamp 1644511149
transform 1 0 4416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1644511149
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_59
timestamp 1644511149
transform 1 0 6532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_67
timestamp 1644511149
transform 1 0 7268 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1644511149
transform 1 0 7544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1644511149
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1644511149
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_142
timestamp 1644511149
transform 1 0 14168 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_150
timestamp 1644511149
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_154
timestamp 1644511149
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1644511149
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_206
timestamp 1644511149
transform 1 0 20056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_212
timestamp 1644511149
transform 1 0 20608 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1644511149
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1644511149
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_255
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_263
timestamp 1644511149
transform 1 0 25300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1644511149
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_287
timestamp 1644511149
transform 1 0 27508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_299
timestamp 1644511149
transform 1 0 28612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1644511149
transform 1 0 29716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_320
timestamp 1644511149
transform 1 0 30544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1644511149
transform 1 0 32660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_355
timestamp 1644511149
transform 1 0 33764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_363
timestamp 1644511149
transform 1 0 34500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_368
timestamp 1644511149
transform 1 0 34960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1644511149
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1644511149
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_61
timestamp 1644511149
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1644511149
transform 1 0 7452 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1644511149
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1644511149
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1644511149
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1644511149
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1644511149
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_168
timestamp 1644511149
transform 1 0 16560 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_179
timestamp 1644511149
transform 1 0 17572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_187
timestamp 1644511149
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1644511149
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1644511149
transform 1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_220
timestamp 1644511149
transform 1 0 21344 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_226
timestamp 1644511149
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_240
timestamp 1644511149
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1644511149
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_296
timestamp 1644511149
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_318
timestamp 1644511149
transform 1 0 30360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_338
timestamp 1644511149
transform 1 0 32200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_350
timestamp 1644511149
transform 1 0 33304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1644511149
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_397
timestamp 1644511149
transform 1 0 37628 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_12
timestamp 1644511149
transform 1 0 2208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_20
timestamp 1644511149
transform 1 0 2944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_43
timestamp 1644511149
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1644511149
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1644511149
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_67
timestamp 1644511149
transform 1 0 7268 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 1644511149
transform 1 0 7820 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_76
timestamp 1644511149
transform 1 0 8096 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_88
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1644511149
transform 1 0 10304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1644511149
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1644511149
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_138
timestamp 1644511149
transform 1 0 13800 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_150
timestamp 1644511149
transform 1 0 14904 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1644511149
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1644511149
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_213
timestamp 1644511149
transform 1 0 20700 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_259
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_287
timestamp 1644511149
transform 1 0 27508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1644511149
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_311
timestamp 1644511149
transform 1 0 29716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_319
timestamp 1644511149
transform 1 0 30452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_322
timestamp 1644511149
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1644511149
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_355
timestamp 1644511149
transform 1 0 33764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_365
timestamp 1644511149
transform 1 0 34684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_372
timestamp 1644511149
transform 1 0 35328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1644511149
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_35
timestamp 1644511149
transform 1 0 4324 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1644511149
transform 1 0 5060 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1644511149
transform 1 0 5796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_59
timestamp 1644511149
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1644511149
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_72
timestamp 1644511149
transform 1 0 7728 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_106
timestamp 1644511149
transform 1 0 10856 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_122
timestamp 1644511149
transform 1 0 12328 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1644511149
transform 1 0 14352 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_152
timestamp 1644511149
transform 1 0 15088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1644511149
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_200
timestamp 1644511149
transform 1 0 19504 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1644511149
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_210
timestamp 1644511149
transform 1 0 20424 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_213
timestamp 1644511149
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1644511149
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1644511149
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1644511149
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_263
timestamp 1644511149
transform 1 0 25300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_283
timestamp 1644511149
transform 1 0 27140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_295
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1644511149
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_318
timestamp 1644511149
transform 1 0 30360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_372
timestamp 1644511149
transform 1 0 35328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_381
timestamp 1644511149
transform 1 0 36156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_393
timestamp 1644511149
transform 1 0 37260 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1644511149
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_61
timestamp 1644511149
transform 1 0 6716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1644511149
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_80
timestamp 1644511149
transform 1 0 8464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_86
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1644511149
transform 1 0 12420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_183
timestamp 1644511149
transform 1 0 17940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_195
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_207
timestamp 1644511149
transform 1 0 20148 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1644511149
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_303
timestamp 1644511149
transform 1 0 28980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_314
timestamp 1644511149
transform 1 0 29992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_320
timestamp 1644511149
transform 1 0 30544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_326
timestamp 1644511149
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1644511149
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_345
timestamp 1644511149
transform 1 0 32844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_351
timestamp 1644511149
transform 1 0 33396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_371
timestamp 1644511149
transform 1 0 35236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1644511149
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_12
timestamp 1644511149
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_20
timestamp 1644511149
transform 1 0 2944 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_35
timestamp 1644511149
transform 1 0 4324 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1644511149
transform 1 0 4968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_54
timestamp 1644511149
transform 1 0 6072 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_57
timestamp 1644511149
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_69
timestamp 1644511149
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1644511149
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1644511149
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_116
timestamp 1644511149
transform 1 0 11776 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_120
timestamp 1644511149
transform 1 0 12144 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1644511149
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1644511149
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_143
timestamp 1644511149
transform 1 0 14260 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_155
timestamp 1644511149
transform 1 0 15364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1644511149
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_171
timestamp 1644511149
transform 1 0 16836 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1644511149
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1644511149
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_235
timestamp 1644511149
transform 1 0 22724 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1644511149
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1644511149
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_328
timestamp 1644511149
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_340
timestamp 1644511149
transform 1 0 32384 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_343
timestamp 1644511149
transform 1 0 32660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1644511149
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_375
timestamp 1644511149
transform 1 0 35604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_395
timestamp 1644511149
transform 1 0 37444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1644511149
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1644511149
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1644511149
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_136
timestamp 1644511149
transform 1 0 13616 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_148
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1644511149
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 1644511149
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_206
timestamp 1644511149
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1644511149
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_232
timestamp 1644511149
transform 1 0 22448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_236
timestamp 1644511149
transform 1 0 22816 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1644511149
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1644511149
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1644511149
transform 1 0 25484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1644511149
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_307
timestamp 1644511149
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_313
timestamp 1644511149
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1644511149
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1644511149
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_365
timestamp 1644511149
transform 1 0 34684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_377
timestamp 1644511149
transform 1 0 35788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1644511149
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp 1644511149
transform 1 0 1656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_12
timestamp 1644511149
transform 1 0 2208 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1644511149
transform 1 0 4048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1644511149
transform 1 0 4692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_46
timestamp 1644511149
transform 1 0 5336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_52
timestamp 1644511149
transform 1 0 5888 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_64
timestamp 1644511149
transform 1 0 6992 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1644511149
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_183
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1644511149
transform 1 0 20240 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1644511149
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_230
timestamp 1644511149
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 1644511149
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1644511149
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1644511149
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_329
timestamp 1644511149
transform 1 0 31372 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_341
timestamp 1644511149
transform 1 0 32476 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_353
timestamp 1644511149
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1644511149
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_369
timestamp 1644511149
transform 1 0 35052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_381
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_393
timestamp 1644511149
transform 1 0 37260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1644511149
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1644511149
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1644511149
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1644511149
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1644511149
transform 1 0 13156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_138
timestamp 1644511149
transform 1 0 13800 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_146
timestamp 1644511149
transform 1 0 14536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_150
timestamp 1644511149
transform 1 0 14904 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1644511149
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_179
timestamp 1644511149
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_191
timestamp 1644511149
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_203
timestamp 1644511149
transform 1 0 19780 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1644511149
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_254
timestamp 1644511149
transform 1 0 24472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1644511149
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_313
timestamp 1644511149
transform 1 0 29900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1644511149
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_324
timestamp 1644511149
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_344
timestamp 1644511149
transform 1 0 32752 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_377
timestamp 1644511149
transform 1 0 35788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_389
timestamp 1644511149
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1644511149
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_35
timestamp 1644511149
transform 1 0 4324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_47
timestamp 1644511149
transform 1 0 5428 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_59
timestamp 1644511149
transform 1 0 6532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1644511149
transform 1 0 7636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_76
timestamp 1644511149
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_88
timestamp 1644511149
transform 1 0 9200 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_100
timestamp 1644511149
transform 1 0 10304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_112
timestamp 1644511149
transform 1 0 11408 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1644511149
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_155
timestamp 1644511149
transform 1 0 15364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_167
timestamp 1644511149
transform 1 0 16468 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1644511149
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_207
timestamp 1644511149
transform 1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1644511149
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1644511149
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1644511149
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_263
timestamp 1644511149
transform 1 0 25300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_295
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1644511149
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_368
timestamp 1644511149
transform 1 0 34960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_374
timestamp 1644511149
transform 1 0 35512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_386
timestamp 1644511149
transform 1 0 36616 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_392
timestamp 1644511149
transform 1 0 37168 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_395
timestamp 1644511149
transform 1 0 37444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_6
timestamp 1644511149
transform 1 0 1656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_20
timestamp 1644511149
transform 1 0 2944 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_42
timestamp 1644511149
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1644511149
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1644511149
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_75
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1644511149
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1644511149
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_134
timestamp 1644511149
transform 1 0 13432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1644511149
transform 1 0 14352 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_202
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_210
timestamp 1644511149
transform 1 0 20424 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1644511149
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1644511149
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1644511149
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_303
timestamp 1644511149
transform 1 0 28980 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_323
timestamp 1644511149
transform 1 0 30820 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_342
timestamp 1644511149
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_354
timestamp 1644511149
transform 1 0 33672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_362
timestamp 1644511149
transform 1 0 34408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_365
timestamp 1644511149
transform 1 0 34684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_376
timestamp 1644511149
transform 1 0 35696 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_50
timestamp 1644511149
transform 1 0 5704 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_62
timestamp 1644511149
transform 1 0 6808 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1644511149
transform 1 0 7268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1644511149
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1644511149
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_88
timestamp 1644511149
transform 1 0 9200 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_100
timestamp 1644511149
transform 1 0 10304 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_185
timestamp 1644511149
transform 1 0 18124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_220
timestamp 1644511149
transform 1 0 21344 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_319
timestamp 1644511149
transform 1 0 30452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_332
timestamp 1644511149
transform 1 0 31648 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_338
timestamp 1644511149
transform 1 0 32200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_341
timestamp 1644511149
transform 1 0 32476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_355
timestamp 1644511149
transform 1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_369
timestamp 1644511149
transform 1 0 35052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_379
timestamp 1644511149
transform 1 0 35972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_400
timestamp 1644511149
transform 1 0 37904 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1644511149
transform 1 0 38456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_16
timestamp 1644511149
transform 1 0 2576 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1644511149
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1644511149
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_92
timestamp 1644511149
transform 1 0 9568 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1644511149
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_122
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_131
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1644511149
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_195
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_203
timestamp 1644511149
transform 1 0 19780 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1644511149
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_228
timestamp 1644511149
transform 1 0 22080 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_234
timestamp 1644511149
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_247
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_253
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1644511149
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_310
timestamp 1644511149
transform 1 0 29624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_318
timestamp 1644511149
transform 1 0 30360 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_323
timestamp 1644511149
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_339
timestamp 1644511149
transform 1 0 32292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_348
timestamp 1644511149
transform 1 0 33120 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_377
timestamp 1644511149
transform 1 0 35788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1644511149
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1644511149
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_66
timestamp 1644511149
transform 1 0 7176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1644511149
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1644511149
transform 1 0 9108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1644511149
transform 1 0 10212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1644511149
transform 1 0 11316 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_123
timestamp 1644511149
transform 1 0 12420 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1644511149
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_148
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_160
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_180
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1644511149
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1644511149
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_281
timestamp 1644511149
transform 1 0 26956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_288
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1644511149
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_373
timestamp 1644511149
transform 1 0 35420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_391
timestamp 1644511149
transform 1 0 37076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp 1644511149
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_68
timestamp 1644511149
transform 1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1644511149
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_84
timestamp 1644511149
transform 1 0 8832 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_96
timestamp 1644511149
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_143
timestamp 1644511149
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_202
timestamp 1644511149
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1644511149
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1644511149
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_235
timestamp 1644511149
transform 1 0 22724 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_243
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_256
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_268
timestamp 1644511149
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_297
timestamp 1644511149
transform 1 0 28428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_303
timestamp 1644511149
transform 1 0 28980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_309
timestamp 1644511149
transform 1 0 29532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_316
timestamp 1644511149
transform 1 0 30176 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1644511149
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_365
timestamp 1644511149
transform 1 0 34684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_377
timestamp 1644511149
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_12
timestamp 1644511149
transform 1 0 2208 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_61
timestamp 1644511149
transform 1 0 6716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_64
timestamp 1644511149
transform 1 0 6992 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_68
timestamp 1644511149
transform 1 0 7360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_75
timestamp 1644511149
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_106
timestamp 1644511149
transform 1 0 10856 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_118
timestamp 1644511149
transform 1 0 11960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_125
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1644511149
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_180
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1644511149
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_226
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1644511149
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1644511149
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_311
timestamp 1644511149
transform 1 0 29716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_336
timestamp 1644511149
transform 1 0 32016 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_348
timestamp 1644511149
transform 1 0 33120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1644511149
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_40
timestamp 1644511149
transform 1 0 4784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1644511149
transform 1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1644511149
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_60
timestamp 1644511149
transform 1 0 6624 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1644511149
transform 1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1644511149
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_89
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1644511149
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1644511149
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1644511149
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_121
timestamp 1644511149
transform 1 0 12236 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_133
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_141
timestamp 1644511149
transform 1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_177
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1644511149
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1644511149
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_229
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_235
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_248
timestamp 1644511149
transform 1 0 23920 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_267
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_291
timestamp 1644511149
transform 1 0 27876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_309
timestamp 1644511149
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_321
timestamp 1644511149
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1644511149
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_354
timestamp 1644511149
transform 1 0 33672 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_366
timestamp 1644511149
transform 1 0 34776 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_380
timestamp 1644511149
transform 1 0 36064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_384
timestamp 1644511149
transform 1 0 36432 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1644511149
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_395
timestamp 1644511149
transform 1 0 37444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_12
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_38
timestamp 1644511149
transform 1 0 4600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_50
timestamp 1644511149
transform 1 0 5704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1644511149
transform 1 0 6440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_63
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_70
timestamp 1644511149
transform 1 0 7544 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1644511149
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_101
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_126
timestamp 1644511149
transform 1 0 12696 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1644511149
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1644511149
transform 1 0 14628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_169
timestamp 1644511149
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_207
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_219
timestamp 1644511149
transform 1 0 21252 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_223
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_243
timestamp 1644511149
transform 1 0 23460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_290
timestamp 1644511149
transform 1 0 27784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1644511149
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_319
timestamp 1644511149
transform 1 0 30452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_332
timestamp 1644511149
transform 1 0 31648 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1644511149
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1644511149
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_374
timestamp 1644511149
transform 1 0 35512 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_382
timestamp 1644511149
transform 1 0 36248 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_399
timestamp 1644511149
transform 1 0 37812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_59
timestamp 1644511149
transform 1 0 6532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_71
timestamp 1644511149
transform 1 0 7636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1644511149
transform 1 0 8740 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_97
timestamp 1644511149
transform 1 0 10028 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_102
timestamp 1644511149
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1644511149
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_117
timestamp 1644511149
transform 1 0 11868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_138
timestamp 1644511149
transform 1 0 13800 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_143
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_184
timestamp 1644511149
transform 1 0 18032 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_232
timestamp 1644511149
transform 1 0 22448 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_242
timestamp 1644511149
transform 1 0 23368 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_250
timestamp 1644511149
transform 1 0 24104 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_262
timestamp 1644511149
transform 1 0 25208 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1644511149
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_301
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_312
timestamp 1644511149
transform 1 0 29808 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1644511149
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_346
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_354
timestamp 1644511149
transform 1 0 33672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_358
timestamp 1644511149
transform 1 0 34040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_366
timestamp 1644511149
transform 1 0 34776 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_35
timestamp 1644511149
transform 1 0 4324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_60
timestamp 1644511149
transform 1 0 6624 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_72
timestamp 1644511149
transform 1 0 7728 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 1644511149
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_166
timestamp 1644511149
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 1644511149
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_217
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_287
timestamp 1644511149
transform 1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_293
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1644511149
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_322
timestamp 1644511149
transform 1 0 30728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_326
timestamp 1644511149
transform 1 0 31096 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_379
timestamp 1644511149
transform 1 0 35972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_386
timestamp 1644511149
transform 1 0 36616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1644511149
transform 1 0 37260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_399
timestamp 1644511149
transform 1 0 37812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_6
timestamp 1644511149
transform 1 0 1656 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1644511149
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_31
timestamp 1644511149
transform 1 0 3956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1644511149
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1644511149
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1644511149
transform 1 0 7912 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1644511149
transform 1 0 9016 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_98
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_148
timestamp 1644511149
transform 1 0 14720 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_175
timestamp 1644511149
transform 1 0 17204 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_187
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_191
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_194
timestamp 1644511149
transform 1 0 18952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_202
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1644511149
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1644511149
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_228
timestamp 1644511149
transform 1 0 22080 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1644511149
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1644511149
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1644511149
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_313
timestamp 1644511149
transform 1 0 29900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_367
timestamp 1644511149
transform 1 0 34868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_374
timestamp 1644511149
transform 1 0 35512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_386
timestamp 1644511149
transform 1 0 36616 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_5
timestamp 1644511149
transform 1 0 1564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_13
timestamp 1644511149
transform 1 0 2300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1644511149
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_50
timestamp 1644511149
transform 1 0 5704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_58
timestamp 1644511149
transform 1 0 6440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_143
timestamp 1644511149
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_175
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_240
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_275
timestamp 1644511149
transform 1 0 26404 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_283
timestamp 1644511149
transform 1 0 27140 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_299
timestamp 1644511149
transform 1 0 28612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_313
timestamp 1644511149
transform 1 0 29900 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_319
timestamp 1644511149
transform 1 0 30452 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_336
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1644511149
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_12
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_24
timestamp 1644511149
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_36
timestamp 1644511149
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_48
timestamp 1644511149
transform 1 0 5520 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1644511149
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_63
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1644511149
transform 1 0 7544 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1644511149
transform 1 0 8648 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1644511149
transform 1 0 9752 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_106
timestamp 1644511149
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_120
timestamp 1644511149
transform 1 0 12144 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_132
timestamp 1644511149
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_142
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_153
timestamp 1644511149
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1644511149
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_177
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_189
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_201
timestamp 1644511149
transform 1 0 19596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_235
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_247
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_259
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_297
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_306
timestamp 1644511149
transform 1 0 29256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_324
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_344
timestamp 1644511149
transform 1 0 32752 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_356
timestamp 1644511149
transform 1 0 33856 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_368
timestamp 1644511149
transform 1 0 34960 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_376
timestamp 1644511149
transform 1 0 35696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1644511149
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_61
timestamp 1644511149
transform 1 0 6716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1644511149
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_104
timestamp 1644511149
transform 1 0 10672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_112
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_116
timestamp 1644511149
transform 1 0 11776 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_124
timestamp 1644511149
transform 1 0 12512 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_185
timestamp 1644511149
transform 1 0 18124 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_200
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_208
timestamp 1644511149
transform 1 0 20240 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1644511149
transform 1 0 20884 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_231
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_276
timestamp 1644511149
transform 1 0 26496 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_284
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_290
timestamp 1644511149
transform 1 0 27784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_317
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_329
timestamp 1644511149
transform 1 0 31372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_338
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_350
timestamp 1644511149
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_373
timestamp 1644511149
transform 1 0 35420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_385
timestamp 1644511149
transform 1 0 36524 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_395
timestamp 1644511149
transform 1 0 37444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_45
timestamp 1644511149
transform 1 0 5244 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_63
timestamp 1644511149
transform 1 0 6900 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_92
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_104
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_206
timestamp 1644511149
transform 1 0 20056 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1644511149
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_233
timestamp 1644511149
transform 1 0 22540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1644511149
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_269
timestamp 1644511149
transform 1 0 25852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_288
timestamp 1644511149
transform 1 0 27600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_300
timestamp 1644511149
transform 1 0 28704 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_312
timestamp 1644511149
transform 1 0 29808 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1644511149
transform 1 0 30728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1644511149
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_359
timestamp 1644511149
transform 1 0 34132 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_371
timestamp 1644511149
transform 1 0 35236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1644511149
transform 1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1644511149
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_12
timestamp 1644511149
transform 1 0 2208 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_18
timestamp 1644511149
transform 1 0 2760 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1644511149
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_32
timestamp 1644511149
transform 1 0 4048 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_40
timestamp 1644511149
transform 1 0 4784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1644511149
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_52
timestamp 1644511149
transform 1 0 5888 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1644511149
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_66
timestamp 1644511149
transform 1 0 7176 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_70
timestamp 1644511149
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_88
timestamp 1644511149
transform 1 0 9200 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_100
timestamp 1644511149
transform 1 0 10304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_112
timestamp 1644511149
transform 1 0 11408 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_118
timestamp 1644511149
transform 1 0 11960 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_154
timestamp 1644511149
transform 1 0 15272 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_283
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_292
timestamp 1644511149
transform 1 0 27968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_373
timestamp 1644511149
transform 1 0 35420 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_390
timestamp 1644511149
transform 1 0 36984 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_402
timestamp 1644511149
transform 1 0 38088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1644511149
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_60
timestamp 1644511149
transform 1 0 6624 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_87
timestamp 1644511149
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1644511149
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1644511149
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_155
timestamp 1644511149
transform 1 0 15364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_175
timestamp 1644511149
transform 1 0 17204 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_187
timestamp 1644511149
transform 1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_211
timestamp 1644511149
transform 1 0 20516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_240
timestamp 1644511149
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_264
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_284
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_296
timestamp 1644511149
transform 1 0 28336 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_302
timestamp 1644511149
transform 1 0 28888 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_318
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1644511149
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_354
timestamp 1644511149
transform 1 0 33672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_358
timestamp 1644511149
transform 1 0 34040 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_368
timestamp 1644511149
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1644511149
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_396
timestamp 1644511149
transform 1 0 37536 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_404
timestamp 1644511149
transform 1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_6
timestamp 1644511149
transform 1 0 1656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_12
timestamp 1644511149
transform 1 0 2208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_70
timestamp 1644511149
transform 1 0 7544 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1644511149
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_128
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_148
timestamp 1644511149
transform 1 0 14720 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_167
timestamp 1644511149
transform 1 0 16468 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1644511149
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_200
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_212
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_224
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_297
timestamp 1644511149
transform 1 0 28428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_340
timestamp 1644511149
transform 1 0 32384 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_346
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_350
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_356
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_371
timestamp 1644511149
transform 1 0 35236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_382
timestamp 1644511149
transform 1 0 36248 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_38
timestamp 1644511149
transform 1 0 4600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_46
timestamp 1644511149
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1644511149
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1644511149
transform 1 0 8648 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1644511149
transform 1 0 9752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1644511149
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_136
timestamp 1644511149
transform 1 0 13616 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1644511149
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1644511149
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1644511149
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1644511149
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_245
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_252
timestamp 1644511149
transform 1 0 24288 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1644511149
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_306
timestamp 1644511149
transform 1 0 29256 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_318
timestamp 1644511149
transform 1 0 30360 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_323
timestamp 1644511149
transform 1 0 30820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_365
timestamp 1644511149
transform 1 0 34684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_368
timestamp 1644511149
transform 1 0 34960 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_383
timestamp 1644511149
transform 1 0 36340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_10
timestamp 1644511149
transform 1 0 2024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp 1644511149
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_35
timestamp 1644511149
transform 1 0 4324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1644511149
transform 1 0 4968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1644511149
transform 1 0 6072 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_66
timestamp 1644511149
transform 1 0 7176 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1644511149
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1644511149
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_95
timestamp 1644511149
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_107
timestamp 1644511149
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_119
timestamp 1644511149
transform 1 0 12052 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_131
timestamp 1644511149
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_158
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_170
timestamp 1644511149
transform 1 0 16744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1644511149
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1644511149
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_234
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_271
timestamp 1644511149
transform 1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_281
timestamp 1644511149
transform 1 0 26956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_287
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_318
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_330
timestamp 1644511149
transform 1 0 31464 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_342
timestamp 1644511149
transform 1 0 32568 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1644511149
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1644511149
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_6
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_12
timestamp 1644511149
transform 1 0 2208 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_18
timestamp 1644511149
transform 1 0 2760 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_22
timestamp 1644511149
transform 1 0 3128 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_32
timestamp 1644511149
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_44
timestamp 1644511149
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_63
timestamp 1644511149
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_66
timestamp 1644511149
transform 1 0 7176 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_72
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_79
timestamp 1644511149
transform 1 0 8372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1644511149
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_140
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_148
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_153
timestamp 1644511149
transform 1 0 15180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_204
timestamp 1644511149
transform 1 0 19872 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1644511149
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_260
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_290
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_296
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_304
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_309
timestamp 1644511149
transform 1 0 29532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_322
timestamp 1644511149
transform 1 0 30728 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1644511149
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_355
timestamp 1644511149
transform 1 0 33764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_366
timestamp 1644511149
transform 1 0 34776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_50
timestamp 1644511149
transform 1 0 5704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_64
timestamp 1644511149
transform 1 0 6992 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_72
timestamp 1644511149
transform 1 0 7728 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1644511149
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_106
timestamp 1644511149
transform 1 0 10856 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_118
timestamp 1644511149
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_122
timestamp 1644511149
transform 1 0 12328 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1644511149
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_155
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_167
timestamp 1644511149
transform 1 0 16468 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_183
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_205
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_219
timestamp 1644511149
transform 1 0 21252 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_256
timestamp 1644511149
transform 1 0 24656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_268
timestamp 1644511149
transform 1 0 25760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_293
timestamp 1644511149
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1644511149
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_320
timestamp 1644511149
transform 1 0 30544 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_332
timestamp 1644511149
transform 1 0 31648 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_344
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1644511149
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_397
timestamp 1644511149
transform 1 0 37628 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1644511149
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_12
timestamp 1644511149
transform 1 0 2208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_24
timestamp 1644511149
transform 1 0 3312 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1644511149
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1644511149
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 1644511149
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_83
timestamp 1644511149
transform 1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_91
timestamp 1644511149
transform 1 0 9476 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1644511149
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1644511149
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_159
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_210
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_246
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_258
timestamp 1644511149
transform 1 0 24840 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_264
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_302
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_312
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_354
timestamp 1644511149
transform 1 0 33672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_369
timestamp 1644511149
transform 1 0 35052 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_375
timestamp 1644511149
transform 1 0 35604 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1644511149
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_35
timestamp 1644511149
transform 1 0 4324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_42
timestamp 1644511149
transform 1 0 4968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_48
timestamp 1644511149
transform 1 0 5520 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_60
timestamp 1644511149
transform 1 0 6624 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_66
timestamp 1644511149
transform 1 0 7176 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_70
timestamp 1644511149
transform 1 0 7544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1644511149
transform 1 0 9660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1644511149
transform 1 0 11868 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_129
timestamp 1644511149
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1644511149
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_147
timestamp 1644511149
transform 1 0 14628 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_159
timestamp 1644511149
transform 1 0 15732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_163
timestamp 1644511149
transform 1 0 16100 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_174
timestamp 1644511149
transform 1 0 17112 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1644511149
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_205
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_212
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_218
timestamp 1644511149
transform 1 0 21160 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_225
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_239
timestamp 1644511149
transform 1 0 23092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_273
timestamp 1644511149
transform 1 0 26220 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_297
timestamp 1644511149
transform 1 0 28428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1644511149
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_314
timestamp 1644511149
transform 1 0 29992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_326
timestamp 1644511149
transform 1 0 31096 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_332
timestamp 1644511149
transform 1 0 31648 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_344
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_352
timestamp 1644511149
transform 1 0 33488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_369
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_376
timestamp 1644511149
transform 1 0 35696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_382
timestamp 1644511149
transform 1 0 36248 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_394
timestamp 1644511149
transform 1 0 37352 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1644511149
transform 1 0 38456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_34
timestamp 1644511149
transform 1 0 4232 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_46
timestamp 1644511149
transform 1 0 5336 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1644511149
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_73
timestamp 1644511149
transform 1 0 7820 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_80
timestamp 1644511149
transform 1 0 8464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_86
timestamp 1644511149
transform 1 0 9016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_91
timestamp 1644511149
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1644511149
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_143
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_155
timestamp 1644511149
transform 1 0 15364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_175
timestamp 1644511149
transform 1 0 17204 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_187
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_199
timestamp 1644511149
transform 1 0 19412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1644511149
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_228
timestamp 1644511149
transform 1 0 22080 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_240
timestamp 1644511149
transform 1 0 23184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_252
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_264
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_287
timestamp 1644511149
transform 1 0 27508 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_304
timestamp 1644511149
transform 1 0 29072 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_316
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_321
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_342
timestamp 1644511149
transform 1 0 32568 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_354
timestamp 1644511149
transform 1 0 33672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_364
timestamp 1644511149
transform 1 0 34592 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_378
timestamp 1644511149
transform 1 0 35880 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_387
timestamp 1644511149
transform 1 0 36708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_6
timestamp 1644511149
transform 1 0 1656 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_12
timestamp 1644511149
transform 1 0 2208 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_20
timestamp 1644511149
transform 1 0 2944 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_35
timestamp 1644511149
transform 1 0 4324 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_47
timestamp 1644511149
transform 1 0 5428 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_59
timestamp 1644511149
transform 1 0 6532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_71
timestamp 1644511149
transform 1 0 7636 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_88
timestamp 1644511149
transform 1 0 9200 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_100
timestamp 1644511149
transform 1 0 10304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_112
timestamp 1644511149
transform 1 0 11408 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_124
timestamp 1644511149
transform 1 0 12512 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_151
timestamp 1644511149
transform 1 0 14996 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_169
timestamp 1644511149
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_211
timestamp 1644511149
transform 1 0 20516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_223
timestamp 1644511149
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1644511149
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_298
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_387
timestamp 1644511149
transform 1 0 36708 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_395
timestamp 1644511149
transform 1 0 37444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_9
timestamp 1644511149
transform 1 0 1932 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_20
timestamp 1644511149
transform 1 0 2944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1644511149
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1644511149
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1644511149
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_142
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_156
timestamp 1644511149
transform 1 0 15456 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1644511149
transform 1 0 16928 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_184
timestamp 1644511149
transform 1 0 18032 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_190
timestamp 1644511149
transform 1 0 18584 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_212
timestamp 1644511149
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_228
timestamp 1644511149
transform 1 0 22080 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_238
timestamp 1644511149
transform 1 0 23000 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_246
timestamp 1644511149
transform 1 0 23736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_255
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_267
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_301
timestamp 1644511149
transform 1 0 28796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_307
timestamp 1644511149
transform 1 0 29348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_319
timestamp 1644511149
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1644511149
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_365
timestamp 1644511149
transform 1 0 34684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_12
timestamp 1644511149
transform 1 0 2208 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_20
timestamp 1644511149
transform 1 0 2944 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_50
timestamp 1644511149
transform 1 0 5704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_58
timestamp 1644511149
transform 1 0 6440 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_63
timestamp 1644511149
transform 1 0 6900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_69
timestamp 1644511149
transform 1 0 7452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 1644511149
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_88
timestamp 1644511149
transform 1 0 9200 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_95
timestamp 1644511149
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_107
timestamp 1644511149
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_122
timestamp 1644511149
transform 1 0 12328 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_151
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_163
timestamp 1644511149
transform 1 0 16100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_200
timestamp 1644511149
transform 1 0 19504 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_240
timestamp 1644511149
transform 1 0 23184 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1644511149
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1644511149
transform 1 0 24840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_295
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_373
timestamp 1644511149
transform 1 0 35420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_399
timestamp 1644511149
transform 1 0 37812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_14
timestamp 1644511149
transform 1 0 2392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_46
timestamp 1644511149
transform 1 0 5336 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_68
timestamp 1644511149
transform 1 0 7360 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_74
timestamp 1644511149
transform 1 0 7912 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1644511149
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_146
timestamp 1644511149
transform 1 0 14536 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1644511149
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_172
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_178
timestamp 1644511149
transform 1 0 17480 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_200
timestamp 1644511149
transform 1 0 19504 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_212
timestamp 1644511149
transform 1 0 20608 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_235
timestamp 1644511149
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_247
timestamp 1644511149
transform 1 0 23828 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_287
timestamp 1644511149
transform 1 0 27508 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_330
timestamp 1644511149
transform 1 0 31464 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_371
timestamp 1644511149
transform 1 0 35236 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_383
timestamp 1644511149
transform 1 0 36340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_399
timestamp 1644511149
transform 1 0 37812 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_5
timestamp 1644511149
transform 1 0 1564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_17
timestamp 1644511149
transform 1 0 2668 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1644511149
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_49
timestamp 1644511149
transform 1 0 5612 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_58
timestamp 1644511149
transform 1 0 6440 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_70
timestamp 1644511149
transform 1 0 7544 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1644511149
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_106
timestamp 1644511149
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_118
timestamp 1644511149
transform 1 0 11960 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_129
timestamp 1644511149
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1644511149
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_183
timestamp 1644511149
transform 1 0 17940 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_219
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_237
timestamp 1644511149
transform 1 0 22908 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1644511149
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_272
timestamp 1644511149
transform 1 0 26128 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_284
timestamp 1644511149
transform 1 0 27232 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_295
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_330
timestamp 1644511149
transform 1 0 31464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_334
timestamp 1644511149
transform 1 0 31832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1644511149
transform 1 0 32108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1644511149
transform 1 0 33212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1644511149
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_6
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_22
timestamp 1644511149
transform 1 0 3128 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_34
timestamp 1644511149
transform 1 0 4232 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_46
timestamp 1644511149
transform 1 0 5336 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_60
timestamp 1644511149
transform 1 0 6624 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_66
timestamp 1644511149
transform 1 0 7176 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_71
timestamp 1644511149
transform 1 0 7636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_77
timestamp 1644511149
transform 1 0 8188 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_88
timestamp 1644511149
transform 1 0 9200 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_100
timestamp 1644511149
transform 1 0 10304 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_119
timestamp 1644511149
transform 1 0 12052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_123
timestamp 1644511149
transform 1 0 12420 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_129
timestamp 1644511149
transform 1 0 12972 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1644511149
transform 1 0 14996 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1644511149
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_201
timestamp 1644511149
transform 1 0 19596 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1644511149
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_253
timestamp 1644511149
transform 1 0 24380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_259
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_291
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_303
timestamp 1644511149
transform 1 0 28980 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_311
timestamp 1644511149
transform 1 0 29716 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_322
timestamp 1644511149
transform 1 0 30728 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_344
timestamp 1644511149
transform 1 0 32752 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_356
timestamp 1644511149
transform 1 0 33856 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1644511149
transform 1 0 34408 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_375
timestamp 1644511149
transform 1 0 35604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_387
timestamp 1644511149
transform 1 0 36708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_45
timestamp 1644511149
transform 1 0 5244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_70
timestamp 1644511149
transform 1 0 7544 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1644511149
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1644511149
transform 1 0 14352 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_156
timestamp 1644511149
transform 1 0 15456 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_203
timestamp 1644511149
transform 1 0 19780 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_218
timestamp 1644511149
transform 1 0 21160 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_226
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_231
timestamp 1644511149
transform 1 0 22356 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_350
timestamp 1644511149
transform 1 0 33304 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1644511149
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_12
timestamp 1644511149
transform 1 0 2208 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_24
timestamp 1644511149
transform 1 0 3312 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_36
timestamp 1644511149
transform 1 0 4416 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_40
timestamp 1644511149
transform 1 0 4784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1644511149
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_83
timestamp 1644511149
transform 1 0 8740 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_95
timestamp 1644511149
transform 1 0 9844 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_107
timestamp 1644511149
transform 1 0 10948 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_121
timestamp 1644511149
transform 1 0 12236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_144
timestamp 1644511149
transform 1 0 14352 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_158
timestamp 1644511149
transform 1 0 15640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1644511149
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_175
timestamp 1644511149
transform 1 0 17204 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_190
timestamp 1644511149
transform 1 0 18584 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_197
timestamp 1644511149
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_204
timestamp 1644511149
transform 1 0 19872 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1644511149
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_230
timestamp 1644511149
transform 1 0 22264 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_244
timestamp 1644511149
transform 1 0 23552 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_250
timestamp 1644511149
transform 1 0 24104 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_266
timestamp 1644511149
transform 1 0 25576 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_318
timestamp 1644511149
transform 1 0 30360 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_330
timestamp 1644511149
transform 1 0 31464 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_342
timestamp 1644511149
transform 1 0 32568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_346
timestamp 1644511149
transform 1 0 32936 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_363
timestamp 1644511149
transform 1 0 34500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_375
timestamp 1644511149
transform 1 0 35604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1644511149
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_38
timestamp 1644511149
transform 1 0 4600 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_46
timestamp 1644511149
transform 1 0 5336 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_52
timestamp 1644511149
transform 1 0 5888 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_64
timestamp 1644511149
transform 1 0 6992 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_72
timestamp 1644511149
transform 1 0 7728 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_91
timestamp 1644511149
transform 1 0 9476 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_103
timestamp 1644511149
transform 1 0 10580 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_115
timestamp 1644511149
transform 1 0 11684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_123
timestamp 1644511149
transform 1 0 12420 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_127
timestamp 1644511149
transform 1 0 12788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_151
timestamp 1644511149
transform 1 0 14996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_157
timestamp 1644511149
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_164
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1644511149
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_206
timestamp 1644511149
transform 1 0 20056 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_213
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_257
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_279
timestamp 1644511149
transform 1 0 26772 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_315
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_319
timestamp 1644511149
transform 1 0 30452 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_322
timestamp 1644511149
transform 1 0 30728 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_334
timestamp 1644511149
transform 1 0 31832 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_346
timestamp 1644511149
transform 1 0 32936 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_358
timestamp 1644511149
transform 1 0 34040 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_5
timestamp 1644511149
transform 1 0 1564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_35
timestamp 1644511149
transform 1 0 4324 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_45
timestamp 1644511149
transform 1 0 5244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_85
timestamp 1644511149
transform 1 0 8924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_89
timestamp 1644511149
transform 1 0 9292 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_101
timestamp 1644511149
transform 1 0 10396 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_109
timestamp 1644511149
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_121
timestamp 1644511149
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_144
timestamp 1644511149
transform 1 0 14352 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 1644511149
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1644511149
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_188
timestamp 1644511149
transform 1 0 18400 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_200
timestamp 1644511149
transform 1 0 19504 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_213
timestamp 1644511149
transform 1 0 20700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1644511149
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_240
timestamp 1644511149
transform 1 0 23184 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_252
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_267
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_302
timestamp 1644511149
transform 1 0 28888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_313
timestamp 1644511149
transform 1 0 29900 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_321
timestamp 1644511149
transform 1 0 30636 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_14
timestamp 1644511149
transform 1 0 2392 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_32
timestamp 1644511149
transform 1 0 4048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_42
timestamp 1644511149
transform 1 0 4968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_52
timestamp 1644511149
transform 1 0 5888 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_58
timestamp 1644511149
transform 1 0 6440 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_70
timestamp 1644511149
transform 1 0 7544 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1644511149
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_88
timestamp 1644511149
transform 1 0 9200 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_95
timestamp 1644511149
transform 1 0 9844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_107
timestamp 1644511149
transform 1 0 10948 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_119
timestamp 1644511149
transform 1 0 12052 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_123
timestamp 1644511149
transform 1 0 12420 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_127
timestamp 1644511149
transform 1 0 12788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_157
timestamp 1644511149
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_164
timestamp 1644511149
transform 1 0 16192 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_176
timestamp 1644511149
transform 1 0 17296 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_184
timestamp 1644511149
transform 1 0 18032 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_191
timestamp 1644511149
transform 1 0 18676 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_261
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_285
timestamp 1644511149
transform 1 0 27324 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_297
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_311
timestamp 1644511149
transform 1 0 29716 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_317
timestamp 1644511149
transform 1 0 30268 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_320
timestamp 1644511149
transform 1 0 30544 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_326
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_355
timestamp 1644511149
transform 1 0 33764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_393
timestamp 1644511149
transform 1 0 37260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_396
timestamp 1644511149
transform 1 0 37536 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_23
timestamp 1644511149
transform 1 0 3220 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_35
timestamp 1644511149
transform 1 0 4324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_45
timestamp 1644511149
transform 1 0 5244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_65
timestamp 1644511149
transform 1 0 7084 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_71
timestamp 1644511149
transform 1 0 7636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_82
timestamp 1644511149
transform 1 0 8648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1644511149
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_136
timestamp 1644511149
transform 1 0 13616 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_150
timestamp 1644511149
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_154
timestamp 1644511149
transform 1 0 15272 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_158
timestamp 1644511149
transform 1 0 15640 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1644511149
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1644511149
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1644511149
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_243
timestamp 1644511149
transform 1 0 23460 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_254
timestamp 1644511149
transform 1 0 24472 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_268
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1644511149
transform 1 0 28796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_311
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_323
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_331
timestamp 1644511149
transform 1 0 31556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_340
timestamp 1644511149
transform 1 0 32384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_352
timestamp 1644511149
transform 1 0 33488 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_364
timestamp 1644511149
transform 1 0 34592 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_376
timestamp 1644511149
transform 1 0 35696 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_11
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_34
timestamp 1644511149
transform 1 0 4232 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_59
timestamp 1644511149
transform 1 0 6532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_67
timestamp 1644511149
transform 1 0 7268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_71
timestamp 1644511149
transform 1 0 7636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_106
timestamp 1644511149
transform 1 0 10856 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_114
timestamp 1644511149
transform 1 0 11592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1644511149
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_151
timestamp 1644511149
transform 1 0 14996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_155
timestamp 1644511149
transform 1 0 15364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_181
timestamp 1644511149
transform 1 0 17756 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_225
timestamp 1644511149
transform 1 0 21804 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_232
timestamp 1644511149
transform 1 0 22448 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1644511149
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_274
timestamp 1644511149
transform 1 0 26312 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_286
timestamp 1644511149
transform 1 0 27416 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_294
timestamp 1644511149
transform 1 0 28152 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_298
timestamp 1644511149
transform 1 0 28520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1644511149
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_38
timestamp 1644511149
transform 1 0 4600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1644511149
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1644511149
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_65
timestamp 1644511149
transform 1 0 7084 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_88
timestamp 1644511149
transform 1 0 9200 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_100
timestamp 1644511149
transform 1 0 10304 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_104
timestamp 1644511149
transform 1 0 10672 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1644511149
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_155
timestamp 1644511149
transform 1 0 15364 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_159
timestamp 1644511149
transform 1 0 15732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_191
timestamp 1644511149
transform 1 0 18676 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_235
timestamp 1644511149
transform 1 0 22724 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_264
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_271
timestamp 1644511149
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_312
timestamp 1644511149
transform 1 0 29808 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_324
timestamp 1644511149
transform 1 0 30912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1644511149
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_36
timestamp 1644511149
transform 1 0 4416 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_61
timestamp 1644511149
transform 1 0 6716 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_73
timestamp 1644511149
transform 1 0 7820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1644511149
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_106
timestamp 1644511149
transform 1 0 10856 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_114
timestamp 1644511149
transform 1 0 11592 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_120
timestamp 1644511149
transform 1 0 12144 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_129
timestamp 1644511149
transform 1 0 12972 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_162
timestamp 1644511149
transform 1 0 16008 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_170
timestamp 1644511149
transform 1 0 16744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_215
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1644511149
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_244
timestamp 1644511149
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_256
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_285
timestamp 1644511149
transform 1 0 27324 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_297
timestamp 1644511149
transform 1 0 28428 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1644511149
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1644511149
transform 1 0 32108 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1644511149
transform 1 0 33212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_361
timestamp 1644511149
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_38
timestamp 1644511149
transform 1 0 4600 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1644511149
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1644511149
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_87
timestamp 1644511149
transform 1 0 9108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_152
timestamp 1644511149
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_178
timestamp 1644511149
transform 1 0 17480 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_190
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_202
timestamp 1644511149
transform 1 0 19688 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_250
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_262
timestamp 1644511149
transform 1 0 25208 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_268
timestamp 1644511149
transform 1 0 25760 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_311
timestamp 1644511149
transform 1 0 29716 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_326
timestamp 1644511149
transform 1 0 31096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1644511149
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_173
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_185
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_229
timestamp 1644511149
transform 1 0 22172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_313
timestamp 1644511149
transform 1 0 29900 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_318
timestamp 1644511149
transform 1 0 30360 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_330
timestamp 1644511149
transform 1 0 31464 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1644511149
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0687_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0688_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0689_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18768 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0690_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0692_
timestamp 1644511149
transform 1 0 5152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0693_
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0694_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0695_
timestamp 1644511149
transform 1 0 22080 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0696_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0697_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0698_
timestamp 1644511149
transform 1 0 2392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0699_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3312 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0700_
timestamp 1644511149
transform 1 0 20056 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0701_
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1644511149
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0703_
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0704_
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0705_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0706_
timestamp 1644511149
transform -1 0 3312 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0707_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0708_
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1644511149
transform -1 0 22080 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0710_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0711_
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0712_
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0713_
timestamp 1644511149
transform 1 0 25576 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 1644511149
transform -1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0715_
timestamp 1644511149
transform -1 0 21344 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0716_
timestamp 1644511149
transform 1 0 21712 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0717_
timestamp 1644511149
transform 1 0 22448 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0718_
timestamp 1644511149
transform 1 0 21896 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0719_
timestamp 1644511149
transform -1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0720_
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0721_
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0722_
timestamp 1644511149
transform 1 0 21712 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0723_
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0724_
timestamp 1644511149
transform 1 0 14260 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0725_
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0726_
timestamp 1644511149
transform 1 0 20792 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0727_
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0728_
timestamp 1644511149
transform -1 0 20884 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0729_
timestamp 1644511149
transform -1 0 20240 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0730_
timestamp 1644511149
transform -1 0 16376 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0732_
timestamp 1644511149
transform -1 0 16192 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0733_
timestamp 1644511149
transform -1 0 15088 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0734_
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1644511149
transform -1 0 15824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0736_
timestamp 1644511149
transform -1 0 14996 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0738_
timestamp 1644511149
transform -1 0 14720 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0739_
timestamp 1644511149
transform -1 0 14076 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0740_
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0742_
timestamp 1644511149
transform -1 0 13432 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1644511149
transform 1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0744_
timestamp 1644511149
transform -1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0745_
timestamp 1644511149
transform -1 0 11868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0746_
timestamp 1644511149
transform 1 0 14536 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 1644511149
transform 1 0 14996 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0748_
timestamp 1644511149
transform -1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0749_
timestamp 1644511149
transform 1 0 11500 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0750_
timestamp 1644511149
transform -1 0 13248 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1644511149
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0753_
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0755_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0756_
timestamp 1644511149
transform 1 0 3036 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0757_
timestamp 1644511149
transform 1 0 18584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0758_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0759_
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0760_
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0761_
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0762_
timestamp 1644511149
transform -1 0 19688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0763_
timestamp 1644511149
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1644511149
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0765_
timestamp 1644511149
transform 1 0 3128 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0766_
timestamp 1644511149
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0767_
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0768_
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0769_
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0770_
timestamp 1644511149
transform -1 0 33120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0771_
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0772_
timestamp 1644511149
transform -1 0 14444 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0773_
timestamp 1644511149
transform -1 0 13616 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 1644511149
transform 1 0 15088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0775_
timestamp 1644511149
transform -1 0 14628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 1644511149
transform 1 0 12604 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0777_
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1644511149
transform -1 0 16284 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0779_
timestamp 1644511149
transform 1 0 14904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1644511149
transform 1 0 14168 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0781_
timestamp 1644511149
transform 1 0 15088 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1644511149
transform -1 0 17112 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0783_
timestamp 1644511149
transform 1 0 15088 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 1644511149
transform -1 0 17756 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0785_
timestamp 1644511149
transform -1 0 14536 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0786_
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0787_
timestamp 1644511149
transform 1 0 16192 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0788_
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0789_
timestamp 1644511149
transform -1 0 14628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0790_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0791_
timestamp 1644511149
transform -1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0792_
timestamp 1644511149
transform -1 0 13616 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0793_
timestamp 1644511149
transform -1 0 15088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0795_
timestamp 1644511149
transform -1 0 14260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0796_
timestamp 1644511149
transform -1 0 13616 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0797_
timestamp 1644511149
transform 1 0 15364 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0798_
timestamp 1644511149
transform -1 0 13616 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0799_
timestamp 1644511149
transform 1 0 14996 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0800_
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1644511149
transform -1 0 16928 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0802_
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0803_
timestamp 1644511149
transform 1 0 14904 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 1644511149
transform -1 0 15640 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0805_
timestamp 1644511149
transform -1 0 14996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0806_
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0807_
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0808_
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0809_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0810_
timestamp 1644511149
transform -1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0811_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0812_
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0813_
timestamp 1644511149
transform 1 0 22172 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0814_
timestamp 1644511149
transform 1 0 22908 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0815_
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0816_
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0817_
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0818_
timestamp 1644511149
transform -1 0 18492 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0819_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 1644511149
transform -1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0821_
timestamp 1644511149
transform 1 0 15640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0822_
timestamp 1644511149
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0823_
timestamp 1644511149
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1644511149
transform -1 0 7452 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0825_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 1644511149
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0827_
timestamp 1644511149
transform 1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0828_
timestamp 1644511149
transform 1 0 11040 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0829_
timestamp 1644511149
transform -1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0830_
timestamp 1644511149
transform -1 0 7728 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0832_
timestamp 1644511149
transform 1 0 10580 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0833_
timestamp 1644511149
transform -1 0 7268 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0834_
timestamp 1644511149
transform 1 0 7728 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0835_
timestamp 1644511149
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0836_
timestamp 1644511149
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0837_
timestamp 1644511149
transform -1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0838_
timestamp 1644511149
transform 1 0 7912 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0839_
timestamp 1644511149
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0840_
timestamp 1644511149
transform -1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0841_
timestamp 1644511149
transform -1 0 5612 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0842_
timestamp 1644511149
transform -1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0843_
timestamp 1644511149
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0844_
timestamp 1644511149
transform 1 0 4508 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0845_
timestamp 1644511149
transform -1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1644511149
transform -1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0847_
timestamp 1644511149
transform 1 0 4784 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0848_
timestamp 1644511149
transform -1 0 4324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0850_
timestamp 1644511149
transform -1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1644511149
transform -1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0852_
timestamp 1644511149
transform -1 0 4232 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 1644511149
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0854_
timestamp 1644511149
transform 1 0 4416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1644511149
transform 1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0856_
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 1644511149
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0858_
timestamp 1644511149
transform -1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0859_
timestamp 1644511149
transform -1 0 4324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1644511149
transform -1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0861_
timestamp 1644511149
transform -1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0862_
timestamp 1644511149
transform -1 0 4324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0863_
timestamp 1644511149
transform -1 0 3312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0864_
timestamp 1644511149
transform -1 0 3956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 1644511149
transform -1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0866_
timestamp 1644511149
transform -1 0 3864 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0867_
timestamp 1644511149
transform -1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0868_
timestamp 1644511149
transform 1 0 4416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1644511149
transform 1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0870_
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0871_
timestamp 1644511149
transform 1 0 4692 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1644511149
transform 1 0 5060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0873_
timestamp 1644511149
transform -1 0 4048 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 1644511149
transform -1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0875_
timestamp 1644511149
transform -1 0 6992 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0876_
timestamp 1644511149
transform -1 0 4232 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 1644511149
transform -1 0 3312 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0878_
timestamp 1644511149
transform -1 0 4324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0879_
timestamp 1644511149
transform -1 0 2944 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1644511149
transform -1 0 4324 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1644511149
transform -1 0 3312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0882_
timestamp 1644511149
transform -1 0 6900 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0883_
timestamp 1644511149
transform -1 0 7360 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0884_
timestamp 1644511149
transform 1 0 5888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0885_
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1644511149
transform -1 0 7636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0887_
timestamp 1644511149
transform 1 0 6900 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1644511149
transform -1 0 7636 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0889_
timestamp 1644511149
transform -1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0890_
timestamp 1644511149
transform -1 0 9476 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1644511149
transform -1 0 9200 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0892_
timestamp 1644511149
transform 1 0 7912 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1644511149
transform -1 0 8648 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0894_
timestamp 1644511149
transform 1 0 8188 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1644511149
transform 1 0 9568 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1644511149
transform -1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1644511149
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0900_
timestamp 1644511149
transform 1 0 21620 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1644511149
transform -1 0 22448 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0902_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7912 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0904_
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0905_
timestamp 1644511149
transform 1 0 23552 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0906_
timestamp 1644511149
transform 1 0 23000 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1644511149
transform -1 0 24932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0908_
timestamp 1644511149
transform 1 0 23828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0910_
timestamp 1644511149
transform 1 0 21620 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0911_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0912_
timestamp 1644511149
transform 1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 1644511149
transform 1 0 19596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0914_
timestamp 1644511149
transform -1 0 19780 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1644511149
transform 1 0 18308 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1644511149
transform -1 0 17204 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0918_
timestamp 1644511149
transform -1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0919_
timestamp 1644511149
transform -1 0 15640 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0920_
timestamp 1644511149
transform -1 0 16192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0921_
timestamp 1644511149
transform -1 0 14996 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0922_
timestamp 1644511149
transform -1 0 17112 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0923_
timestamp 1644511149
transform -1 0 15640 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0924_
timestamp 1644511149
transform -1 0 16192 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0925_
timestamp 1644511149
transform -1 0 14904 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0926_
timestamp 1644511149
transform -1 0 20056 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0927_
timestamp 1644511149
transform -1 0 20700 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0928_
timestamp 1644511149
transform 1 0 18124 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 1644511149
transform -1 0 17664 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 1644511149
transform -1 0 20700 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1644511149
transform -1 0 20792 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0932_
timestamp 1644511149
transform -1 0 19964 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0933_
timestamp 1644511149
transform 1 0 19044 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0934_
timestamp 1644511149
transform -1 0 20884 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1644511149
transform -1 0 18768 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0936_
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0938_
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1644511149
transform -1 0 22724 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0940_
timestamp 1644511149
transform 1 0 22724 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0941_
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0942_
timestamp 1644511149
transform 1 0 22632 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0943_
timestamp 1644511149
transform 1 0 24840 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0944_
timestamp 1644511149
transform -1 0 22080 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1644511149
transform 1 0 22908 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0946_
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1644511149
transform -1 0 24840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0948_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0949_
timestamp 1644511149
transform 1 0 25668 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0950_
timestamp 1644511149
transform 1 0 23368 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1644511149
transform -1 0 25024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0953_
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1644511149
transform -1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1644511149
transform -1 0 21712 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1644511149
transform -1 0 22172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0957_
timestamp 1644511149
transform 1 0 22816 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0958_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0959_
timestamp 1644511149
transform 1 0 22908 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1644511149
transform -1 0 24564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0961_
timestamp 1644511149
transform -1 0 10488 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0962_
timestamp 1644511149
transform -1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0963_
timestamp 1644511149
transform 1 0 22816 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1644511149
transform -1 0 25208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0965_
timestamp 1644511149
transform 1 0 21988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0966_
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0967_
timestamp 1644511149
transform 1 0 22724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0968_
timestamp 1644511149
transform 1 0 23736 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0969_
timestamp 1644511149
transform -1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1644511149
transform -1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0971_
timestamp 1644511149
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1644511149
transform -1 0 7544 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1644511149
transform -1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0974_
timestamp 1644511149
transform 1 0 7544 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0975_
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0976_
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1644511149
transform 1 0 7636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0979_
timestamp 1644511149
transform 1 0 6808 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1644511149
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0981_
timestamp 1644511149
transform 1 0 6624 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1644511149
transform -1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0983_
timestamp 1644511149
transform 1 0 7452 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1644511149
transform -1 0 8648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1644511149
transform -1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1644511149
transform 1 0 5612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0988_
timestamp 1644511149
transform -1 0 6900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1644511149
transform 1 0 5428 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0990_
timestamp 1644511149
transform 1 0 6164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1644511149
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0993_
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1644511149
transform -1 0 7544 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0995_
timestamp 1644511149
transform 1 0 6256 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1644511149
transform 1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0997_
timestamp 1644511149
transform -1 0 5888 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1644511149
transform -1 0 7452 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1644511149
transform -1 0 7544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1644511149
transform -1 0 8096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1002_
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1644511149
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1004_
timestamp 1644511149
transform 1 0 7820 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1644511149
transform 1 0 9844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1006_
timestamp 1644511149
transform 1 0 7820 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1007_
timestamp 1644511149
transform 1 0 7912 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1644511149
transform -1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1644511149
transform 1 0 7912 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1644511149
transform -1 0 9200 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1644511149
transform 1 0 7912 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform -1 0 8464 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1644511149
transform 1 0 4968 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1644511149
transform 1 0 5520 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1644511149
transform -1 0 5428 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1016_
timestamp 1644511149
transform -1 0 5244 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1018_
timestamp 1644511149
transform -1 0 4600 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1019_
timestamp 1644511149
transform -1 0 4324 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1644511149
transform -1 0 9476 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1021_
timestamp 1644511149
transform 1 0 4416 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1023_
timestamp 1644511149
transform -1 0 5244 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1644511149
transform -1 0 4232 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1025_
timestamp 1644511149
transform -1 0 5888 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1026_
timestamp 1644511149
transform -1 0 3312 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1027_
timestamp 1644511149
transform 1 0 9108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1644511149
transform 1 0 9292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1029_
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1644511149
transform -1 0 21988 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1031_
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1644511149
transform 1 0 22172 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1033_
timestamp 1644511149
transform 1 0 21252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1644511149
transform -1 0 22632 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1035_
timestamp 1644511149
transform -1 0 20608 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1036_
timestamp 1644511149
transform -1 0 20516 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1037_
timestamp 1644511149
transform 1 0 22448 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1038_
timestamp 1644511149
transform 1 0 28244 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1039_
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1040_
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1041_
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1042_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1043_
timestamp 1644511149
transform 1 0 25576 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1044_
timestamp 1644511149
transform 1 0 27324 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1045_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1046_
timestamp 1644511149
transform 1 0 29808 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1047_
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1048_
timestamp 1644511149
transform 1 0 17848 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1049_
timestamp 1644511149
transform 1 0 20884 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1050_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1051_
timestamp 1644511149
transform 1 0 20240 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1644511149
transform -1 0 22080 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1053_
timestamp 1644511149
transform -1 0 17572 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1644511149
transform -1 0 16836 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1056_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1057_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1644511149
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1059_
timestamp 1644511149
transform -1 0 17388 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1644511149
transform -1 0 16192 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1644511149
transform -1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1062_
timestamp 1644511149
transform 1 0 13156 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1063_
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1644511149
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1065_
timestamp 1644511149
transform -1 0 13616 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1644511149
transform 1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1067_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1068_
timestamp 1644511149
transform -1 0 15364 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1069_
timestamp 1644511149
transform -1 0 12788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1070_
timestamp 1644511149
transform -1 0 12328 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1071_
timestamp 1644511149
transform -1 0 12696 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1644511149
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1073_
timestamp 1644511149
transform -1 0 13616 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1644511149
transform -1 0 12420 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1075_
timestamp 1644511149
transform -1 0 13800 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1076_
timestamp 1644511149
transform -1 0 13432 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1077_
timestamp 1644511149
transform -1 0 14352 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1079_
timestamp 1644511149
transform -1 0 18768 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1644511149
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1081_
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform -1 0 19504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1083_
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1084_
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1085_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29624 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1644511149
transform -1 0 36800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1087_
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1644511149
transform -1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1089_
timestamp 1644511149
transform 1 0 33764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1090_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35696 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 36340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1092_
timestamp 1644511149
transform -1 0 35604 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1093_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35512 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1094_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1096_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1097_
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1098_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1644511149
transform -1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1100_
timestamp 1644511149
transform 1 0 29900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1644511149
transform 1 0 32384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1102_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1103_
timestamp 1644511149
transform -1 0 30728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1104_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34868 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1105_
timestamp 1644511149
transform -1 0 30268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform -1 0 32752 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _1107_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1108_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19504 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _1109_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20240 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1110_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1111_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1112_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1113_
timestamp 1644511149
transform -1 0 33304 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1114_
timestamp 1644511149
transform -1 0 28888 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1115_
timestamp 1644511149
transform -1 0 28796 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1644511149
transform -1 0 28520 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1117_
timestamp 1644511149
transform -1 0 29900 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1118_
timestamp 1644511149
transform 1 0 29256 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1119_
timestamp 1644511149
transform -1 0 29808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1120_
timestamp 1644511149
transform 1 0 30728 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1121_
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1644511149
transform -1 0 32384 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1123_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1124_
timestamp 1644511149
transform -1 0 27968 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1126_
timestamp 1644511149
transform 1 0 29992 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1127_
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1128_
timestamp 1644511149
transform -1 0 29256 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1130_
timestamp 1644511149
transform 1 0 20700 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1131_
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1644511149
transform -1 0 32292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1134_
timestamp 1644511149
transform -1 0 31648 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1135_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1136_
timestamp 1644511149
transform -1 0 35512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 1644511149
transform 1 0 35144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1138_
timestamp 1644511149
transform 1 0 35880 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1139_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36984 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1140_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1141_
timestamp 1644511149
transform 1 0 28612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1142_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34408 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1143_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1144_
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1145_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1146_
timestamp 1644511149
transform 1 0 28888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1147_
timestamp 1644511149
transform 1 0 30360 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1644511149
transform 1 0 30176 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1150_
timestamp 1644511149
transform 1 0 29900 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1151_
timestamp 1644511149
transform 1 0 29900 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1152_
timestamp 1644511149
transform -1 0 30544 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1153_
timestamp 1644511149
transform 1 0 29256 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1154_
timestamp 1644511149
transform 1 0 26956 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1155_
timestamp 1644511149
transform -1 0 26496 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1156_
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1157_
timestamp 1644511149
transform -1 0 30360 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1644511149
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1160_
timestamp 1644511149
transform 1 0 30544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1161_
timestamp 1644511149
transform -1 0 31648 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1644511149
transform -1 0 35696 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1164_
timestamp 1644511149
transform -1 0 27784 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1644511149
transform -1 0 29348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1167_
timestamp 1644511149
transform -1 0 27876 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1168_
timestamp 1644511149
transform 1 0 28612 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1644511149
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1170_
timestamp 1644511149
transform 1 0 29624 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1644511149
transform -1 0 30636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1173_
timestamp 1644511149
transform 1 0 34132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1174_
timestamp 1644511149
transform 1 0 35696 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1644511149
transform -1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1177_
timestamp 1644511149
transform 1 0 31372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1178_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31648 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _1179_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35420 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1180_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35604 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1181_
timestamp 1644511149
transform -1 0 34960 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1644511149
transform -1 0 36340 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1184_
timestamp 1644511149
transform 1 0 35696 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1185_
timestamp 1644511149
transform -1 0 35236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1186_
timestamp 1644511149
transform 1 0 34960 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 1644511149
transform -1 0 35052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1188_
timestamp 1644511149
transform -1 0 37444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1189_
timestamp 1644511149
transform -1 0 36524 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1644511149
transform 1 0 34040 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1191_
timestamp 1644511149
transform 1 0 33856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1192_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34040 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1193_
timestamp 1644511149
transform -1 0 36708 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1194_
timestamp 1644511149
transform -1 0 35696 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1195_
timestamp 1644511149
transform -1 0 35420 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1196_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34132 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1644511149
transform -1 0 33304 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1644511149
transform -1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1199_
timestamp 1644511149
transform 1 0 22816 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1201_
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _1202_
timestamp 1644511149
transform -1 0 20056 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1644511149
transform 1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1204_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1205_
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1206_
timestamp 1644511149
transform -1 0 23000 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1208_
timestamp 1644511149
transform -1 0 17296 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1209_
timestamp 1644511149
transform 1 0 16744 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1211_
timestamp 1644511149
transform -1 0 16376 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1644511149
transform -1 0 16192 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1644511149
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1214_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1215_
timestamp 1644511149
transform -1 0 14996 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1216_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1217_
timestamp 1644511149
transform -1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1218_
timestamp 1644511149
transform -1 0 13708 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1219_
timestamp 1644511149
transform -1 0 13432 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1220_
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1221_
timestamp 1644511149
transform -1 0 10948 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1222_
timestamp 1644511149
transform -1 0 10580 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1644511149
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1224_
timestamp 1644511149
transform -1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1225_
timestamp 1644511149
transform -1 0 9936 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1644511149
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1227_
timestamp 1644511149
transform -1 0 20516 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1228_
timestamp 1644511149
transform -1 0 19872 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1229_
timestamp 1644511149
transform -1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1644511149
transform -1 0 22908 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1231_
timestamp 1644511149
transform -1 0 23644 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1644511149
transform 1 0 26864 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1644511149
transform 1 0 24656 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 1644511149
transform -1 0 23736 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1235_
timestamp 1644511149
transform 1 0 23276 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1644511149
transform -1 0 24840 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1644511149
transform -1 0 24656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1238_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1239_
timestamp 1644511149
transform 1 0 29348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1644511149
transform -1 0 35052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1241_
timestamp 1644511149
transform -1 0 35788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1242_
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1243_
timestamp 1644511149
transform 1 0 30636 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1244_
timestamp 1644511149
transform -1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1245_
timestamp 1644511149
transform 1 0 27968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1246_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1247_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 1644511149
transform 1 0 29256 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1249_
timestamp 1644511149
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1250_
timestamp 1644511149
transform -1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1644511149
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1644511149
transform 1 0 30176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1253_
timestamp 1644511149
transform -1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1254_
timestamp 1644511149
transform 1 0 25944 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1255_
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1256_
timestamp 1644511149
transform -1 0 29992 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1257_
timestamp 1644511149
transform -1 0 29992 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1644511149
transform 1 0 30084 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1644511149
transform -1 0 30820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1644511149
transform 1 0 34132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1644511149
transform -1 0 36156 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1262_
timestamp 1644511149
transform -1 0 35328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1263_
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1264_
timestamp 1644511149
transform -1 0 34132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1265_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28980 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1644511149
transform -1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1267_
timestamp 1644511149
transform 1 0 30084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 1644511149
transform -1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1269_
timestamp 1644511149
transform 1 0 33856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1270_
timestamp 1644511149
transform -1 0 34776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1271_
timestamp 1644511149
transform -1 0 35420 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1272_
timestamp 1644511149
transform 1 0 20792 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 1644511149
transform -1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1644511149
transform -1 0 34408 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1275_
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1276_
timestamp 1644511149
transform 1 0 33396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1644511149
transform -1 0 33028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1278_
timestamp 1644511149
transform 1 0 32752 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1279_
timestamp 1644511149
transform -1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1280_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35604 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1644511149
transform 1 0 33028 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1644511149
transform -1 0 29164 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1644511149
transform -1 0 31004 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1644511149
transform -1 0 32660 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1644511149
transform -1 0 27140 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1644511149
transform 1 0 32200 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1644511149
transform 1 0 36340 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1644511149
transform 1 0 30544 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1644511149
transform 1 0 27600 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1292_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1293_
timestamp 1644511149
transform 1 0 36340 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1294_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1644511149
transform -1 0 30820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1644511149
transform 1 0 35512 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1644511149
transform 1 0 35328 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1644511149
transform 1 0 36340 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1644511149
transform 1 0 33764 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1644511149
transform 1 0 35236 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1644511149
transform 1 0 32200 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1644511149
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1644511149
transform 1 0 12696 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1644511149
transform 1 0 12144 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1644511149
transform -1 0 9752 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1311_
timestamp 1644511149
transform 1 0 24564 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1644511149
transform 1 0 35972 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1644511149
transform 1 0 33764 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1644511149
transform 1 0 25668 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1315_
timestamp 1644511149
transform -1 0 31096 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1316_
timestamp 1644511149
transform 1 0 36340 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1317_
timestamp 1644511149
transform 1 0 25300 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1644511149
transform 1 0 30728 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1644511149
transform -1 0 29072 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1644511149
transform 1 0 29440 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1644511149
transform 1 0 35328 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1644511149
transform -1 0 35972 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1644511149
transform 1 0 32752 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1644511149
transform 1 0 31556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1326__36 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1327__37
timestamp 1644511149
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1328__38
timestamp 1644511149
transform 1 0 13524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1329__39
timestamp 1644511149
transform -1 0 12972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1330__40
timestamp 1644511149
transform -1 0 10672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1331__41
timestamp 1644511149
transform -1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1332__42
timestamp 1644511149
transform 1 0 10028 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1333__43
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1334__44
timestamp 1644511149
transform -1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1335__45
timestamp 1644511149
transform -1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1336__46
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1337__47
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1338__48
timestamp 1644511149
transform -1 0 17940 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1339__49
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1340__50
timestamp 1644511149
transform 1 0 12512 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1341__51
timestamp 1644511149
transform 1 0 12512 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1342__52
timestamp 1644511149
transform 1 0 11868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1343__53
timestamp 1644511149
transform -1 0 18400 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1344__54
timestamp 1644511149
transform 1 0 17204 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1345__55
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1346__56
timestamp 1644511149
transform 1 0 20976 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1347__57
timestamp 1644511149
transform -1 0 24656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1348__58
timestamp 1644511149
transform -1 0 25760 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1349__59
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1350__60
timestamp 1644511149
transform -1 0 8004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1351__61
timestamp 1644511149
transform -1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1352__62
timestamp 1644511149
transform 1 0 6992 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1353__63
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1354__64
timestamp 1644511149
transform -1 0 9292 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1355__65
timestamp 1644511149
transform -1 0 4968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1356__66
timestamp 1644511149
transform 1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1357__67
timestamp 1644511149
transform -1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1358__68
timestamp 1644511149
transform -1 0 7544 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1359__69
timestamp 1644511149
transform -1 0 3128 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1360__70
timestamp 1644511149
transform -1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1361__71
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1362__72
timestamp 1644511149
transform -1 0 9844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1363__73
timestamp 1644511149
transform -1 0 9200 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1364__74
timestamp 1644511149
transform 1 0 8280 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1365__75
timestamp 1644511149
transform -1 0 2760 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1366__76
timestamp 1644511149
transform -1 0 3036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1367__77
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1368__78
timestamp 1644511149
transform 1 0 4140 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1369__79
timestamp 1644511149
transform -1 0 5244 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1370__80
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1371__81
timestamp 1644511149
transform -1 0 23092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1372__82
timestamp 1644511149
transform -1 0 22080 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1373__83
timestamp 1644511149
transform -1 0 24656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1374__84
timestamp 1644511149
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1375__85
timestamp 1644511149
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1376__86
timestamp 1644511149
transform -1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1377__87
timestamp 1644511149
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1378__88
timestamp 1644511149
transform -1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1379__89
timestamp 1644511149
transform -1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1380__90
timestamp 1644511149
transform 1 0 2760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1381__91
timestamp 1644511149
transform -1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1382__92
timestamp 1644511149
transform -1 0 5152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1383__93
timestamp 1644511149
transform -1 0 3128 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1384__94
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1385__95
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1386__96
timestamp 1644511149
transform 1 0 2024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1387__97
timestamp 1644511149
transform -1 0 3036 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1388__98
timestamp 1644511149
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1389__99
timestamp 1644511149
transform -1 0 5888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1390__100
timestamp 1644511149
transform -1 0 7636 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1391__101
timestamp 1644511149
transform -1 0 9292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1392__102
timestamp 1644511149
transform 1 0 8832 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1393__103
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1394__104
timestamp 1644511149
transform -1 0 22540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1395__105
timestamp 1644511149
transform 1 0 25760 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1396__106
timestamp 1644511149
transform -1 0 25668 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1397__107
timestamp 1644511149
transform -1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1398__108
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1399__109
timestamp 1644511149
transform -1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1400__110
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1401__111
timestamp 1644511149
transform -1 0 12604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1402__112
timestamp 1644511149
transform 1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1403__113
timestamp 1644511149
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1404__114
timestamp 1644511149
transform -1 0 10672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1405__115
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1406__116
timestamp 1644511149
transform -1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1407__117
timestamp 1644511149
transform -1 0 17204 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1408__118
timestamp 1644511149
transform -1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1409__119
timestamp 1644511149
transform -1 0 18308 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1410__120
timestamp 1644511149
transform -1 0 17204 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1411__121
timestamp 1644511149
transform 1 0 12696 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1412__122
timestamp 1644511149
transform 1 0 12052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1413__123
timestamp 1644511149
transform 1 0 12144 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1414__124
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1415__125
timestamp 1644511149
transform -1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1416__126
timestamp 1644511149
transform -1 0 15732 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1417__127
timestamp 1644511149
transform 1 0 12696 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1418__128
timestamp 1644511149
transform -1 0 17020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1419__129
timestamp 1644511149
transform -1 0 18492 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1420__130
timestamp 1644511149
transform -1 0 12328 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1421__131
timestamp 1644511149
transform -1 0 23184 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1422__132
timestamp 1644511149
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1423__133
timestamp 1644511149
transform 1 0 37904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1424__134
timestamp 1644511149
transform 1 0 37904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1425_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33856 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1426_
timestamp 1644511149
transform -1 0 31464 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1427_
timestamp 1644511149
transform 1 0 27140 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1428_
timestamp 1644511149
transform 1 0 28428 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1429_
timestamp 1644511149
transform 1 0 30728 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1430_
timestamp 1644511149
transform -1 0 24748 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1431_
timestamp 1644511149
transform -1 0 24748 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1432_
timestamp 1644511149
transform -1 0 26588 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1433_
timestamp 1644511149
transform 1 0 17204 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1434_
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1435_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1436_
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1437_
timestamp 1644511149
transform 1 0 10396 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1438_
timestamp 1644511149
transform 1 0 9108 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1439_
timestamp 1644511149
transform -1 0 11776 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1440_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1441_
timestamp 1644511149
transform 1 0 11684 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1442_
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1443_
timestamp 1644511149
transform -1 0 20516 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1444_
timestamp 1644511149
transform -1 0 22540 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1445_
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1446_
timestamp 1644511149
transform -1 0 14996 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1447_
timestamp 1644511149
transform -1 0 14352 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1448_
timestamp 1644511149
transform -1 0 14352 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1449_
timestamp 1644511149
transform -1 0 13708 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1450_
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1451_
timestamp 1644511149
transform -1 0 18768 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1452_
timestamp 1644511149
transform -1 0 16008 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1453_
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1454_
timestamp 1644511149
transform 1 0 23460 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1455_
timestamp 1644511149
transform 1 0 25392 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1456_
timestamp 1644511149
transform 1 0 25208 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1457_
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1458_
timestamp 1644511149
transform -1 0 28060 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1459_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1460_
timestamp 1644511149
transform -1 0 26496 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1461_
timestamp 1644511149
transform -1 0 27232 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1462_
timestamp 1644511149
transform -1 0 27508 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1463_
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1464_
timestamp 1644511149
transform -1 0 26404 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1465_
timestamp 1644511149
transform 1 0 7728 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1466_
timestamp 1644511149
transform 1 0 8464 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1467_
timestamp 1644511149
transform 1 0 7636 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1468_
timestamp 1644511149
transform 1 0 7728 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1469_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1470_
timestamp 1644511149
transform 1 0 4692 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1471_
timestamp 1644511149
transform 1 0 6532 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1472_
timestamp 1644511149
transform 1 0 7636 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1473_
timestamp 1644511149
transform 1 0 7176 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1474_
timestamp 1644511149
transform 1 0 2760 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1475_
timestamp 1644511149
transform 1 0 8924 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1476_
timestamp 1644511149
transform -1 0 10856 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1477_
timestamp 1644511149
transform 1 0 8832 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1478_
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1479_
timestamp 1644511149
transform 1 0 8924 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1480_
timestamp 1644511149
transform 1 0 2392 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1481_
timestamp 1644511149
transform 1 0 2668 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1482_
timestamp 1644511149
transform -1 0 20608 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1483_
timestamp 1644511149
transform 1 0 4784 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1484_
timestamp 1644511149
transform 1 0 4600 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1485_
timestamp 1644511149
transform 1 0 2668 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1486_
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1487_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1488_
timestamp 1644511149
transform -1 0 24288 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1489_
timestamp 1644511149
transform 1 0 22264 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1490_
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1491_
timestamp 1644511149
transform 1 0 16560 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1492_
timestamp 1644511149
transform -1 0 14260 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1493_
timestamp 1644511149
transform -1 0 13616 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1494_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1495_
timestamp 1644511149
transform -1 0 10580 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1496_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1497_
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1498_
timestamp 1644511149
transform 1 0 4508 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1499_
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1500_
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1501_
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1502_
timestamp 1644511149
transform 1 0 3956 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1503_
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1504_
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1505_
timestamp 1644511149
transform -1 0 4968 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1506_
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1507_
timestamp 1644511149
transform 1 0 2668 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1508_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1509_
timestamp 1644511149
transform 1 0 3312 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1510_
timestamp 1644511149
transform 1 0 2760 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1511_
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1512_
timestamp 1644511149
transform 1 0 5612 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1513_
timestamp 1644511149
transform 1 0 7268 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1514_
timestamp 1644511149
transform 1 0 9016 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1515_
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1516_
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1517_
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1518_
timestamp 1644511149
transform -1 0 26312 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1519_
timestamp 1644511149
transform 1 0 25392 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1520_
timestamp 1644511149
transform 1 0 24840 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1521_
timestamp 1644511149
transform 1 0 33856 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1522_
timestamp 1644511149
transform -1 0 28796 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1523_
timestamp 1644511149
transform 1 0 25760 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1524_
timestamp 1644511149
transform -1 0 27600 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1525_
timestamp 1644511149
transform -1 0 29164 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1526_
timestamp 1644511149
transform 1 0 22632 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1527_
timestamp 1644511149
transform -1 0 29348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1644511149
transform -1 0 24932 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1644511149
transform -1 0 20056 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1644511149
transform 1 0 13892 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1644511149
transform 1 0 12328 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1644511149
transform 1 0 10764 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1644511149
transform -1 0 12144 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1644511149
transform 1 0 11592 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1644511149
transform 1 0 16836 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1644511149
transform 1 0 17664 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1644511149
transform 1 0 17940 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1644511149
transform -1 0 14536 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1644511149
transform -1 0 13616 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1644511149
transform -1 0 13616 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1644511149
transform 1 0 16652 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1644511149
transform 1 0 15456 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1644511149
transform 1 0 13156 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1644511149
transform 1 0 16744 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1644511149
transform 1 0 12052 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform -1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 28704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform -1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform 1 0 28612 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform -1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform 1 0 31832 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform -1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform -1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform -1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1644511149
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1644511149
transform -1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 37904 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1644511149
transform 1 0 37812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1644511149
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1644511149
transform 1 0 37812 0 1 36992
box -38 -48 406 592
<< labels >>
rlabel metal2 s 9954 39200 10010 40000 6 clk
port 0 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 peripheralBus_address[0]
port 1 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 peripheralBus_address[10]
port 2 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 peripheralBus_address[11]
port 3 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 peripheralBus_address[12]
port 4 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 peripheralBus_address[13]
port 5 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 peripheralBus_address[14]
port 6 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 peripheralBus_address[15]
port 7 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 peripheralBus_address[16]
port 8 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 peripheralBus_address[17]
port 9 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 peripheralBus_address[18]
port 10 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 peripheralBus_address[19]
port 11 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 peripheralBus_address[1]
port 12 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 peripheralBus_address[20]
port 13 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 peripheralBus_address[21]
port 14 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 peripheralBus_address[22]
port 15 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 peripheralBus_address[23]
port 16 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 peripheralBus_address[2]
port 17 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 peripheralBus_address[3]
port 18 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 peripheralBus_address[4]
port 19 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 peripheralBus_address[5]
port 20 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 peripheralBus_address[6]
port 21 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 peripheralBus_address[7]
port 22 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 peripheralBus_address[8]
port 23 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 peripheralBus_address[9]
port 24 nsew signal input
rlabel metal3 s 0 280 800 400 6 peripheralBus_busy
port 25 nsew signal tristate
rlabel metal3 s 0 2864 800 2984 6 peripheralBus_data[0]
port 26 nsew signal bidirectional
rlabel metal3 s 0 16464 800 16584 6 peripheralBus_data[10]
port 27 nsew signal bidirectional
rlabel metal3 s 0 17824 800 17944 6 peripheralBus_data[11]
port 28 nsew signal bidirectional
rlabel metal3 s 0 19184 800 19304 6 peripheralBus_data[12]
port 29 nsew signal bidirectional
rlabel metal3 s 0 20544 800 20664 6 peripheralBus_data[13]
port 30 nsew signal bidirectional
rlabel metal3 s 0 21904 800 22024 6 peripheralBus_data[14]
port 31 nsew signal bidirectional
rlabel metal3 s 0 23264 800 23384 6 peripheralBus_data[15]
port 32 nsew signal bidirectional
rlabel metal3 s 0 24624 800 24744 6 peripheralBus_data[16]
port 33 nsew signal bidirectional
rlabel metal3 s 0 25984 800 26104 6 peripheralBus_data[17]
port 34 nsew signal bidirectional
rlabel metal3 s 0 27344 800 27464 6 peripheralBus_data[18]
port 35 nsew signal bidirectional
rlabel metal3 s 0 28704 800 28824 6 peripheralBus_data[19]
port 36 nsew signal bidirectional
rlabel metal3 s 0 4224 800 4344 6 peripheralBus_data[1]
port 37 nsew signal bidirectional
rlabel metal3 s 0 30064 800 30184 6 peripheralBus_data[20]
port 38 nsew signal bidirectional
rlabel metal3 s 0 31424 800 31544 6 peripheralBus_data[21]
port 39 nsew signal bidirectional
rlabel metal3 s 0 32784 800 32904 6 peripheralBus_data[22]
port 40 nsew signal bidirectional
rlabel metal3 s 0 34144 800 34264 6 peripheralBus_data[23]
port 41 nsew signal bidirectional
rlabel metal3 s 0 34824 800 34944 6 peripheralBus_data[24]
port 42 nsew signal bidirectional
rlabel metal3 s 0 35504 800 35624 6 peripheralBus_data[25]
port 43 nsew signal bidirectional
rlabel metal3 s 0 36184 800 36304 6 peripheralBus_data[26]
port 44 nsew signal bidirectional
rlabel metal3 s 0 36864 800 36984 6 peripheralBus_data[27]
port 45 nsew signal bidirectional
rlabel metal3 s 0 37544 800 37664 6 peripheralBus_data[28]
port 46 nsew signal bidirectional
rlabel metal3 s 0 38224 800 38344 6 peripheralBus_data[29]
port 47 nsew signal bidirectional
rlabel metal3 s 0 5584 800 5704 6 peripheralBus_data[2]
port 48 nsew signal bidirectional
rlabel metal3 s 0 38904 800 39024 6 peripheralBus_data[30]
port 49 nsew signal bidirectional
rlabel metal3 s 0 39584 800 39704 6 peripheralBus_data[31]
port 50 nsew signal bidirectional
rlabel metal3 s 0 6944 800 7064 6 peripheralBus_data[3]
port 51 nsew signal bidirectional
rlabel metal3 s 0 8304 800 8424 6 peripheralBus_data[4]
port 52 nsew signal bidirectional
rlabel metal3 s 0 9664 800 9784 6 peripheralBus_data[5]
port 53 nsew signal bidirectional
rlabel metal3 s 0 11024 800 11144 6 peripheralBus_data[6]
port 54 nsew signal bidirectional
rlabel metal3 s 0 12384 800 12504 6 peripheralBus_data[7]
port 55 nsew signal bidirectional
rlabel metal3 s 0 13744 800 13864 6 peripheralBus_data[8]
port 56 nsew signal bidirectional
rlabel metal3 s 0 15104 800 15224 6 peripheralBus_data[9]
port 57 nsew signal bidirectional
rlabel metal3 s 0 824 800 944 6 peripheralBus_oe
port 58 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 peripheralBus_we
port 59 nsew signal input
rlabel metal2 s 29918 39200 29974 40000 6 rst
port 60 nsew signal input
rlabel metal3 s 39200 1912 40000 2032 6 spi_clk[0]
port 61 nsew signal tristate
rlabel metal3 s 39200 21904 40000 22024 6 spi_clk[1]
port 62 nsew signal tristate
rlabel metal3 s 39200 5856 40000 5976 6 spi_cs[0]
port 63 nsew signal tristate
rlabel metal3 s 39200 25848 40000 25968 6 spi_cs[1]
port 64 nsew signal tristate
rlabel metal3 s 39200 9800 40000 9920 6 spi_en[0]
port 65 nsew signal tristate
rlabel metal3 s 39200 29792 40000 29912 6 spi_en[1]
port 66 nsew signal tristate
rlabel metal3 s 39200 13880 40000 14000 6 spi_miso[0]
port 67 nsew signal input
rlabel metal3 s 39200 33872 40000 33992 6 spi_miso[1]
port 68 nsew signal input
rlabel metal3 s 39200 17824 40000 17944 6 spi_mosi[0]
port 69 nsew signal tristate
rlabel metal3 s 39200 37816 40000 37936 6 spi_mosi[1]
port 70 nsew signal tristate
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 71 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 71 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 72 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
