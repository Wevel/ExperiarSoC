VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 800.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 796.000 4.050 800.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 796.000 82.710 800.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 796.000 90.530 800.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 796.000 98.350 800.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 796.000 106.630 800.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 796.000 114.450 800.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 796.000 122.270 800.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 796.000 130.090 800.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 796.000 137.910 800.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 796.000 145.730 800.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 796.000 154.010 800.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 796.000 11.870 800.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 796.000 161.830 800.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 796.000 169.650 800.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 796.000 177.470 800.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 796.000 185.290 800.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 796.000 193.110 800.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 796.000 200.930 800.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 796.000 209.210 800.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 796.000 217.030 800.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 796.000 224.850 800.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 796.000 232.670 800.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 796.000 19.690 800.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 796.000 240.490 800.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 796.000 248.310 800.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 796.000 256.590 800.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 796.000 264.410 800.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 796.000 272.230 800.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 796.000 280.050 800.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 796.000 287.870 800.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 796.000 295.690 800.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 796.000 27.510 800.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 796.000 35.330 800.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 796.000 43.150 800.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 796.000 50.970 800.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 796.000 59.250 800.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 796.000 67.070 800.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 796.000 74.890 800.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 796.000 303.970 800.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 796.000 382.630 800.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 796.000 390.450 800.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 796.000 398.270 800.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 796.000 406.550 800.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 796.000 414.370 800.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 796.000 422.190 800.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 796.000 430.010 800.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 796.000 437.830 800.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 796.000 445.650 800.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 796.000 453.930 800.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 796.000 311.790 800.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 796.000 461.750 800.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 796.000 469.570 800.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 796.000 477.390 800.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 796.000 485.210 800.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 796.000 493.030 800.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 796.000 500.850 800.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 796.000 509.130 800.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 796.000 516.950 800.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 796.000 524.770 800.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 796.000 532.590 800.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 796.000 319.610 800.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 796.000 540.410 800.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 796.000 548.230 800.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 796.000 556.510 800.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 796.000 564.330 800.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 796.000 572.150 800.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 796.000 579.970 800.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 796.000 587.790 800.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 796.000 595.610 800.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 796.000 327.430 800.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 796.000 335.250 800.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 796.000 343.070 800.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 796.000 350.890 800.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 796.000 359.170 800.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 796.000 366.990 800.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 796.000 374.810 800.000 ;
    END
  END io_out[9]
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 333.240 600.000 333.840 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 466.520 600.000 467.120 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 599.800 600.000 600.400 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 733.080 600.000 733.680 ;
    END
  END jtag_tms
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 66.680 600.000 67.280 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 199.960 600.000 200.560 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 4.000 787.400 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.720 4.000 715.320 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 788.885 ;
      LAYER met1 ;
        RECT 5.130 6.840 595.630 789.780 ;
      LAYER met2 ;
        RECT 5.160 795.720 11.310 796.690 ;
        RECT 12.150 795.720 19.130 796.690 ;
        RECT 19.970 795.720 26.950 796.690 ;
        RECT 27.790 795.720 34.770 796.690 ;
        RECT 35.610 795.720 42.590 796.690 ;
        RECT 43.430 795.720 50.410 796.690 ;
        RECT 51.250 795.720 58.690 796.690 ;
        RECT 59.530 795.720 66.510 796.690 ;
        RECT 67.350 795.720 74.330 796.690 ;
        RECT 75.170 795.720 82.150 796.690 ;
        RECT 82.990 795.720 89.970 796.690 ;
        RECT 90.810 795.720 97.790 796.690 ;
        RECT 98.630 795.720 106.070 796.690 ;
        RECT 106.910 795.720 113.890 796.690 ;
        RECT 114.730 795.720 121.710 796.690 ;
        RECT 122.550 795.720 129.530 796.690 ;
        RECT 130.370 795.720 137.350 796.690 ;
        RECT 138.190 795.720 145.170 796.690 ;
        RECT 146.010 795.720 153.450 796.690 ;
        RECT 154.290 795.720 161.270 796.690 ;
        RECT 162.110 795.720 169.090 796.690 ;
        RECT 169.930 795.720 176.910 796.690 ;
        RECT 177.750 795.720 184.730 796.690 ;
        RECT 185.570 795.720 192.550 796.690 ;
        RECT 193.390 795.720 200.370 796.690 ;
        RECT 201.210 795.720 208.650 796.690 ;
        RECT 209.490 795.720 216.470 796.690 ;
        RECT 217.310 795.720 224.290 796.690 ;
        RECT 225.130 795.720 232.110 796.690 ;
        RECT 232.950 795.720 239.930 796.690 ;
        RECT 240.770 795.720 247.750 796.690 ;
        RECT 248.590 795.720 256.030 796.690 ;
        RECT 256.870 795.720 263.850 796.690 ;
        RECT 264.690 795.720 271.670 796.690 ;
        RECT 272.510 795.720 279.490 796.690 ;
        RECT 280.330 795.720 287.310 796.690 ;
        RECT 288.150 795.720 295.130 796.690 ;
        RECT 295.970 795.720 303.410 796.690 ;
        RECT 304.250 795.720 311.230 796.690 ;
        RECT 312.070 795.720 319.050 796.690 ;
        RECT 319.890 795.720 326.870 796.690 ;
        RECT 327.710 795.720 334.690 796.690 ;
        RECT 335.530 795.720 342.510 796.690 ;
        RECT 343.350 795.720 350.330 796.690 ;
        RECT 351.170 795.720 358.610 796.690 ;
        RECT 359.450 795.720 366.430 796.690 ;
        RECT 367.270 795.720 374.250 796.690 ;
        RECT 375.090 795.720 382.070 796.690 ;
        RECT 382.910 795.720 389.890 796.690 ;
        RECT 390.730 795.720 397.710 796.690 ;
        RECT 398.550 795.720 405.990 796.690 ;
        RECT 406.830 795.720 413.810 796.690 ;
        RECT 414.650 795.720 421.630 796.690 ;
        RECT 422.470 795.720 429.450 796.690 ;
        RECT 430.290 795.720 437.270 796.690 ;
        RECT 438.110 795.720 445.090 796.690 ;
        RECT 445.930 795.720 453.370 796.690 ;
        RECT 454.210 795.720 461.190 796.690 ;
        RECT 462.030 795.720 469.010 796.690 ;
        RECT 469.850 795.720 476.830 796.690 ;
        RECT 477.670 795.720 484.650 796.690 ;
        RECT 485.490 795.720 492.470 796.690 ;
        RECT 493.310 795.720 500.290 796.690 ;
        RECT 501.130 795.720 508.570 796.690 ;
        RECT 509.410 795.720 516.390 796.690 ;
        RECT 517.230 795.720 524.210 796.690 ;
        RECT 525.050 795.720 532.030 796.690 ;
        RECT 532.870 795.720 539.850 796.690 ;
        RECT 540.690 795.720 547.670 796.690 ;
        RECT 548.510 795.720 555.950 796.690 ;
        RECT 556.790 795.720 563.770 796.690 ;
        RECT 564.610 795.720 571.590 796.690 ;
        RECT 572.430 795.720 579.410 796.690 ;
        RECT 580.250 795.720 587.230 796.690 ;
        RECT 588.070 795.720 595.050 796.690 ;
        RECT 5.160 4.280 595.600 795.720 ;
        RECT 5.710 3.555 15.450 4.280 ;
        RECT 16.290 3.555 26.030 4.280 ;
        RECT 26.870 3.555 36.610 4.280 ;
        RECT 37.450 3.555 47.650 4.280 ;
        RECT 48.490 3.555 58.230 4.280 ;
        RECT 59.070 3.555 68.810 4.280 ;
        RECT 69.650 3.555 79.850 4.280 ;
        RECT 80.690 3.555 90.430 4.280 ;
        RECT 91.270 3.555 101.010 4.280 ;
        RECT 101.850 3.555 111.590 4.280 ;
        RECT 112.430 3.555 122.630 4.280 ;
        RECT 123.470 3.555 133.210 4.280 ;
        RECT 134.050 3.555 143.790 4.280 ;
        RECT 144.630 3.555 154.830 4.280 ;
        RECT 155.670 3.555 165.410 4.280 ;
        RECT 166.250 3.555 175.990 4.280 ;
        RECT 176.830 3.555 186.570 4.280 ;
        RECT 187.410 3.555 197.610 4.280 ;
        RECT 198.450 3.555 208.190 4.280 ;
        RECT 209.030 3.555 218.770 4.280 ;
        RECT 219.610 3.555 229.810 4.280 ;
        RECT 230.650 3.555 240.390 4.280 ;
        RECT 241.230 3.555 250.970 4.280 ;
        RECT 251.810 3.555 261.550 4.280 ;
        RECT 262.390 3.555 272.590 4.280 ;
        RECT 273.430 3.555 283.170 4.280 ;
        RECT 284.010 3.555 293.750 4.280 ;
        RECT 294.590 3.555 304.790 4.280 ;
        RECT 305.630 3.555 315.370 4.280 ;
        RECT 316.210 3.555 325.950 4.280 ;
        RECT 326.790 3.555 336.530 4.280 ;
        RECT 337.370 3.555 347.570 4.280 ;
        RECT 348.410 3.555 358.150 4.280 ;
        RECT 358.990 3.555 368.730 4.280 ;
        RECT 369.570 3.555 379.770 4.280 ;
        RECT 380.610 3.555 390.350 4.280 ;
        RECT 391.190 3.555 400.930 4.280 ;
        RECT 401.770 3.555 411.510 4.280 ;
        RECT 412.350 3.555 422.550 4.280 ;
        RECT 423.390 3.555 433.130 4.280 ;
        RECT 433.970 3.555 443.710 4.280 ;
        RECT 444.550 3.555 454.750 4.280 ;
        RECT 455.590 3.555 465.330 4.280 ;
        RECT 466.170 3.555 475.910 4.280 ;
        RECT 476.750 3.555 486.490 4.280 ;
        RECT 487.330 3.555 497.530 4.280 ;
        RECT 498.370 3.555 508.110 4.280 ;
        RECT 508.950 3.555 518.690 4.280 ;
        RECT 519.530 3.555 529.730 4.280 ;
        RECT 530.570 3.555 540.310 4.280 ;
        RECT 541.150 3.555 550.890 4.280 ;
        RECT 551.730 3.555 561.470 4.280 ;
        RECT 562.310 3.555 572.510 4.280 ;
        RECT 573.350 3.555 583.090 4.280 ;
        RECT 583.930 3.555 593.670 4.280 ;
        RECT 594.510 3.555 595.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 794.560 596.000 795.425 ;
        RECT 4.000 787.800 596.000 794.560 ;
        RECT 4.400 786.400 596.000 787.800 ;
        RECT 4.000 779.640 596.000 786.400 ;
        RECT 4.400 778.240 596.000 779.640 ;
        RECT 4.000 771.480 596.000 778.240 ;
        RECT 4.400 770.080 596.000 771.480 ;
        RECT 4.000 764.000 596.000 770.080 ;
        RECT 4.400 762.600 596.000 764.000 ;
        RECT 4.000 755.840 596.000 762.600 ;
        RECT 4.400 754.440 596.000 755.840 ;
        RECT 4.000 747.680 596.000 754.440 ;
        RECT 4.400 746.280 596.000 747.680 ;
        RECT 4.000 739.520 596.000 746.280 ;
        RECT 4.400 738.120 596.000 739.520 ;
        RECT 4.000 734.080 596.000 738.120 ;
        RECT 4.000 732.680 595.600 734.080 ;
        RECT 4.000 732.040 596.000 732.680 ;
        RECT 4.400 730.640 596.000 732.040 ;
        RECT 4.000 723.880 596.000 730.640 ;
        RECT 4.400 722.480 596.000 723.880 ;
        RECT 4.000 715.720 596.000 722.480 ;
        RECT 4.400 714.320 596.000 715.720 ;
        RECT 4.000 707.560 596.000 714.320 ;
        RECT 4.400 706.160 596.000 707.560 ;
        RECT 4.000 700.080 596.000 706.160 ;
        RECT 4.400 698.680 596.000 700.080 ;
        RECT 4.000 691.920 596.000 698.680 ;
        RECT 4.400 690.520 596.000 691.920 ;
        RECT 4.000 683.760 596.000 690.520 ;
        RECT 4.400 682.360 596.000 683.760 ;
        RECT 4.000 675.600 596.000 682.360 ;
        RECT 4.400 674.200 596.000 675.600 ;
        RECT 4.000 668.120 596.000 674.200 ;
        RECT 4.400 666.720 596.000 668.120 ;
        RECT 4.000 659.960 596.000 666.720 ;
        RECT 4.400 658.560 596.000 659.960 ;
        RECT 4.000 651.800 596.000 658.560 ;
        RECT 4.400 650.400 596.000 651.800 ;
        RECT 4.000 643.640 596.000 650.400 ;
        RECT 4.400 642.240 596.000 643.640 ;
        RECT 4.000 636.160 596.000 642.240 ;
        RECT 4.400 634.760 596.000 636.160 ;
        RECT 4.000 628.000 596.000 634.760 ;
        RECT 4.400 626.600 596.000 628.000 ;
        RECT 4.000 619.840 596.000 626.600 ;
        RECT 4.400 618.440 596.000 619.840 ;
        RECT 4.000 611.680 596.000 618.440 ;
        RECT 4.400 610.280 596.000 611.680 ;
        RECT 4.000 604.200 596.000 610.280 ;
        RECT 4.400 602.800 596.000 604.200 ;
        RECT 4.000 600.800 596.000 602.800 ;
        RECT 4.000 599.400 595.600 600.800 ;
        RECT 4.000 596.040 596.000 599.400 ;
        RECT 4.400 594.640 596.000 596.040 ;
        RECT 4.000 587.880 596.000 594.640 ;
        RECT 4.400 586.480 596.000 587.880 ;
        RECT 4.000 579.720 596.000 586.480 ;
        RECT 4.400 578.320 596.000 579.720 ;
        RECT 4.000 571.560 596.000 578.320 ;
        RECT 4.400 570.160 596.000 571.560 ;
        RECT 4.000 564.080 596.000 570.160 ;
        RECT 4.400 562.680 596.000 564.080 ;
        RECT 4.000 555.920 596.000 562.680 ;
        RECT 4.400 554.520 596.000 555.920 ;
        RECT 4.000 547.760 596.000 554.520 ;
        RECT 4.400 546.360 596.000 547.760 ;
        RECT 4.000 539.600 596.000 546.360 ;
        RECT 4.400 538.200 596.000 539.600 ;
        RECT 4.000 532.120 596.000 538.200 ;
        RECT 4.400 530.720 596.000 532.120 ;
        RECT 4.000 523.960 596.000 530.720 ;
        RECT 4.400 522.560 596.000 523.960 ;
        RECT 4.000 515.800 596.000 522.560 ;
        RECT 4.400 514.400 596.000 515.800 ;
        RECT 4.000 507.640 596.000 514.400 ;
        RECT 4.400 506.240 596.000 507.640 ;
        RECT 4.000 500.160 596.000 506.240 ;
        RECT 4.400 498.760 596.000 500.160 ;
        RECT 4.000 492.000 596.000 498.760 ;
        RECT 4.400 490.600 596.000 492.000 ;
        RECT 4.000 483.840 596.000 490.600 ;
        RECT 4.400 482.440 596.000 483.840 ;
        RECT 4.000 475.680 596.000 482.440 ;
        RECT 4.400 474.280 596.000 475.680 ;
        RECT 4.000 468.200 596.000 474.280 ;
        RECT 4.400 467.520 596.000 468.200 ;
        RECT 4.400 466.800 595.600 467.520 ;
        RECT 4.000 466.120 595.600 466.800 ;
        RECT 4.000 460.040 596.000 466.120 ;
        RECT 4.400 458.640 596.000 460.040 ;
        RECT 4.000 451.880 596.000 458.640 ;
        RECT 4.400 450.480 596.000 451.880 ;
        RECT 4.000 443.720 596.000 450.480 ;
        RECT 4.400 442.320 596.000 443.720 ;
        RECT 4.000 436.240 596.000 442.320 ;
        RECT 4.400 434.840 596.000 436.240 ;
        RECT 4.000 428.080 596.000 434.840 ;
        RECT 4.400 426.680 596.000 428.080 ;
        RECT 4.000 419.920 596.000 426.680 ;
        RECT 4.400 418.520 596.000 419.920 ;
        RECT 4.000 411.760 596.000 418.520 ;
        RECT 4.400 410.360 596.000 411.760 ;
        RECT 4.000 404.280 596.000 410.360 ;
        RECT 4.400 402.880 596.000 404.280 ;
        RECT 4.000 396.120 596.000 402.880 ;
        RECT 4.400 394.720 596.000 396.120 ;
        RECT 4.000 387.960 596.000 394.720 ;
        RECT 4.400 386.560 596.000 387.960 ;
        RECT 4.000 379.800 596.000 386.560 ;
        RECT 4.400 378.400 596.000 379.800 ;
        RECT 4.000 371.640 596.000 378.400 ;
        RECT 4.400 370.240 596.000 371.640 ;
        RECT 4.000 364.160 596.000 370.240 ;
        RECT 4.400 362.760 596.000 364.160 ;
        RECT 4.000 356.000 596.000 362.760 ;
        RECT 4.400 354.600 596.000 356.000 ;
        RECT 4.000 347.840 596.000 354.600 ;
        RECT 4.400 346.440 596.000 347.840 ;
        RECT 4.000 339.680 596.000 346.440 ;
        RECT 4.400 338.280 596.000 339.680 ;
        RECT 4.000 334.240 596.000 338.280 ;
        RECT 4.000 332.840 595.600 334.240 ;
        RECT 4.000 332.200 596.000 332.840 ;
        RECT 4.400 330.800 596.000 332.200 ;
        RECT 4.000 324.040 596.000 330.800 ;
        RECT 4.400 322.640 596.000 324.040 ;
        RECT 4.000 315.880 596.000 322.640 ;
        RECT 4.400 314.480 596.000 315.880 ;
        RECT 4.000 307.720 596.000 314.480 ;
        RECT 4.400 306.320 596.000 307.720 ;
        RECT 4.000 300.240 596.000 306.320 ;
        RECT 4.400 298.840 596.000 300.240 ;
        RECT 4.000 292.080 596.000 298.840 ;
        RECT 4.400 290.680 596.000 292.080 ;
        RECT 4.000 283.920 596.000 290.680 ;
        RECT 4.400 282.520 596.000 283.920 ;
        RECT 4.000 275.760 596.000 282.520 ;
        RECT 4.400 274.360 596.000 275.760 ;
        RECT 4.000 268.280 596.000 274.360 ;
        RECT 4.400 266.880 596.000 268.280 ;
        RECT 4.000 260.120 596.000 266.880 ;
        RECT 4.400 258.720 596.000 260.120 ;
        RECT 4.000 251.960 596.000 258.720 ;
        RECT 4.400 250.560 596.000 251.960 ;
        RECT 4.000 243.800 596.000 250.560 ;
        RECT 4.400 242.400 596.000 243.800 ;
        RECT 4.000 236.320 596.000 242.400 ;
        RECT 4.400 234.920 596.000 236.320 ;
        RECT 4.000 228.160 596.000 234.920 ;
        RECT 4.400 226.760 596.000 228.160 ;
        RECT 4.000 220.000 596.000 226.760 ;
        RECT 4.400 218.600 596.000 220.000 ;
        RECT 4.000 211.840 596.000 218.600 ;
        RECT 4.400 210.440 596.000 211.840 ;
        RECT 4.000 204.360 596.000 210.440 ;
        RECT 4.400 202.960 596.000 204.360 ;
        RECT 4.000 200.960 596.000 202.960 ;
        RECT 4.000 199.560 595.600 200.960 ;
        RECT 4.000 196.200 596.000 199.560 ;
        RECT 4.400 194.800 596.000 196.200 ;
        RECT 4.000 188.040 596.000 194.800 ;
        RECT 4.400 186.640 596.000 188.040 ;
        RECT 4.000 179.880 596.000 186.640 ;
        RECT 4.400 178.480 596.000 179.880 ;
        RECT 4.000 171.720 596.000 178.480 ;
        RECT 4.400 170.320 596.000 171.720 ;
        RECT 4.000 164.240 596.000 170.320 ;
        RECT 4.400 162.840 596.000 164.240 ;
        RECT 4.000 156.080 596.000 162.840 ;
        RECT 4.400 154.680 596.000 156.080 ;
        RECT 4.000 147.920 596.000 154.680 ;
        RECT 4.400 146.520 596.000 147.920 ;
        RECT 4.000 139.760 596.000 146.520 ;
        RECT 4.400 138.360 596.000 139.760 ;
        RECT 4.000 132.280 596.000 138.360 ;
        RECT 4.400 130.880 596.000 132.280 ;
        RECT 4.000 124.120 596.000 130.880 ;
        RECT 4.400 122.720 596.000 124.120 ;
        RECT 4.000 115.960 596.000 122.720 ;
        RECT 4.400 114.560 596.000 115.960 ;
        RECT 4.000 107.800 596.000 114.560 ;
        RECT 4.400 106.400 596.000 107.800 ;
        RECT 4.000 100.320 596.000 106.400 ;
        RECT 4.400 98.920 596.000 100.320 ;
        RECT 4.000 92.160 596.000 98.920 ;
        RECT 4.400 90.760 596.000 92.160 ;
        RECT 4.000 84.000 596.000 90.760 ;
        RECT 4.400 82.600 596.000 84.000 ;
        RECT 4.000 75.840 596.000 82.600 ;
        RECT 4.400 74.440 596.000 75.840 ;
        RECT 4.000 68.360 596.000 74.440 ;
        RECT 4.400 67.680 596.000 68.360 ;
        RECT 4.400 66.960 595.600 67.680 ;
        RECT 4.000 66.280 595.600 66.960 ;
        RECT 4.000 60.200 596.000 66.280 ;
        RECT 4.400 58.800 596.000 60.200 ;
        RECT 4.000 52.040 596.000 58.800 ;
        RECT 4.400 50.640 596.000 52.040 ;
        RECT 4.000 43.880 596.000 50.640 ;
        RECT 4.400 42.480 596.000 43.880 ;
        RECT 4.000 36.400 596.000 42.480 ;
        RECT 4.400 35.000 596.000 36.400 ;
        RECT 4.000 28.240 596.000 35.000 ;
        RECT 4.400 26.840 596.000 28.240 ;
        RECT 4.000 20.080 596.000 26.840 ;
        RECT 4.400 18.680 596.000 20.080 ;
        RECT 4.000 11.920 596.000 18.680 ;
        RECT 4.400 10.520 596.000 11.920 ;
        RECT 4.000 4.440 596.000 10.520 ;
        RECT 4.400 3.575 596.000 4.440 ;
      LAYER met4 ;
        RECT 16.855 19.895 20.640 780.465 ;
        RECT 23.040 19.895 97.440 780.465 ;
        RECT 99.840 19.895 174.240 780.465 ;
        RECT 176.640 19.895 251.040 780.465 ;
        RECT 253.440 19.895 327.840 780.465 ;
        RECT 330.240 19.895 404.640 780.465 ;
        RECT 407.040 19.895 481.440 780.465 ;
        RECT 483.840 19.895 558.240 780.465 ;
        RECT 560.640 19.895 581.145 780.465 ;
  END
END Peripherals
END LIBRARY

