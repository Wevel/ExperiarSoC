magic
tech sky130A
magscale 1 2
timestamp 1683844190
<< obsli1 >>
rect 1104 2159 78844 82705
<< obsm1 >>
rect 566 76 79934 84108
<< metal2 >>
rect 570 84200 626 85000
rect 1306 84200 1362 85000
rect 2042 84200 2098 85000
rect 2778 84200 2834 85000
rect 3514 84200 3570 85000
rect 4250 84200 4306 85000
rect 4986 84200 5042 85000
rect 5722 84200 5778 85000
rect 6458 84200 6514 85000
rect 7194 84200 7250 85000
rect 7930 84200 7986 85000
rect 8666 84200 8722 85000
rect 9402 84200 9458 85000
rect 10138 84200 10194 85000
rect 10874 84200 10930 85000
rect 11610 84200 11666 85000
rect 12346 84200 12402 85000
rect 13082 84200 13138 85000
rect 13818 84200 13874 85000
rect 14554 84200 14610 85000
rect 15290 84200 15346 85000
rect 16026 84200 16082 85000
rect 16762 84200 16818 85000
rect 17498 84200 17554 85000
rect 18234 84200 18290 85000
rect 18970 84200 19026 85000
rect 19706 84200 19762 85000
rect 20442 84200 20498 85000
rect 21178 84200 21234 85000
rect 21914 84200 21970 85000
rect 22650 84200 22706 85000
rect 23386 84200 23442 85000
rect 24122 84200 24178 85000
rect 24858 84200 24914 85000
rect 25594 84200 25650 85000
rect 26330 84200 26386 85000
rect 27066 84200 27122 85000
rect 27802 84200 27858 85000
rect 28538 84200 28594 85000
rect 29274 84200 29330 85000
rect 30010 84200 30066 85000
rect 30746 84200 30802 85000
rect 31482 84200 31538 85000
rect 32218 84200 32274 85000
rect 32954 84200 33010 85000
rect 33690 84200 33746 85000
rect 34426 84200 34482 85000
rect 35162 84200 35218 85000
rect 35898 84200 35954 85000
rect 36634 84200 36690 85000
rect 37370 84200 37426 85000
rect 38106 84200 38162 85000
rect 38842 84200 38898 85000
rect 39578 84200 39634 85000
rect 40314 84200 40370 85000
rect 41050 84200 41106 85000
rect 41786 84200 41842 85000
rect 42522 84200 42578 85000
rect 43258 84200 43314 85000
rect 43994 84200 44050 85000
rect 44730 84200 44786 85000
rect 45466 84200 45522 85000
rect 46202 84200 46258 85000
rect 46938 84200 46994 85000
rect 47674 84200 47730 85000
rect 48410 84200 48466 85000
rect 49146 84200 49202 85000
rect 49882 84200 49938 85000
rect 50618 84200 50674 85000
rect 51354 84200 51410 85000
rect 52090 84200 52146 85000
rect 52826 84200 52882 85000
rect 53562 84200 53618 85000
rect 54298 84200 54354 85000
rect 55034 84200 55090 85000
rect 55770 84200 55826 85000
rect 56506 84200 56562 85000
rect 57242 84200 57298 85000
rect 57978 84200 58034 85000
rect 58714 84200 58770 85000
rect 59450 84200 59506 85000
rect 60186 84200 60242 85000
rect 60922 84200 60978 85000
rect 61658 84200 61714 85000
rect 62394 84200 62450 85000
rect 63130 84200 63186 85000
rect 63866 84200 63922 85000
rect 64602 84200 64658 85000
rect 65338 84200 65394 85000
rect 66074 84200 66130 85000
rect 66810 84200 66866 85000
rect 67546 84200 67602 85000
rect 68282 84200 68338 85000
rect 69018 84200 69074 85000
rect 69754 84200 69810 85000
rect 70490 84200 70546 85000
rect 71226 84200 71282 85000
rect 71962 84200 72018 85000
rect 72698 84200 72754 85000
rect 73434 84200 73490 85000
rect 74170 84200 74226 85000
rect 74906 84200 74962 85000
rect 75642 84200 75698 85000
rect 76378 84200 76434 85000
rect 77114 84200 77170 85000
rect 77850 84200 77906 85000
rect 78586 84200 78642 85000
rect 79322 84200 79378 85000
rect 1306 0 1362 800
rect 2042 0 2098 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14554 0 14610 800
rect 15290 0 15346 800
rect 16026 0 16082 800
rect 16762 0 16818 800
rect 17498 0 17554 800
rect 18234 0 18290 800
rect 18970 0 19026 800
rect 19706 0 19762 800
rect 20442 0 20498 800
rect 21178 0 21234 800
rect 21914 0 21970 800
rect 22650 0 22706 800
rect 23386 0 23442 800
rect 24122 0 24178 800
rect 24858 0 24914 800
rect 25594 0 25650 800
rect 26330 0 26386 800
rect 27066 0 27122 800
rect 27802 0 27858 800
rect 28538 0 28594 800
rect 29274 0 29330 800
rect 30010 0 30066 800
rect 30746 0 30802 800
rect 31482 0 31538 800
rect 32218 0 32274 800
rect 32954 0 33010 800
rect 33690 0 33746 800
rect 34426 0 34482 800
rect 35162 0 35218 800
rect 35898 0 35954 800
rect 36634 0 36690 800
rect 37370 0 37426 800
rect 38106 0 38162 800
rect 38842 0 38898 800
rect 39578 0 39634 800
rect 40314 0 40370 800
rect 41050 0 41106 800
rect 41786 0 41842 800
rect 42522 0 42578 800
rect 43258 0 43314 800
rect 43994 0 44050 800
rect 44730 0 44786 800
rect 45466 0 45522 800
rect 46202 0 46258 800
rect 46938 0 46994 800
rect 47674 0 47730 800
rect 48410 0 48466 800
rect 49146 0 49202 800
rect 49882 0 49938 800
rect 50618 0 50674 800
rect 51354 0 51410 800
rect 52090 0 52146 800
rect 52826 0 52882 800
rect 53562 0 53618 800
rect 54298 0 54354 800
rect 55034 0 55090 800
rect 55770 0 55826 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57978 0 58034 800
rect 58714 0 58770 800
rect 59450 0 59506 800
rect 60186 0 60242 800
rect 60922 0 60978 800
rect 61658 0 61714 800
rect 62394 0 62450 800
rect 63130 0 63186 800
rect 63866 0 63922 800
rect 64602 0 64658 800
rect 65338 0 65394 800
rect 66074 0 66130 800
rect 66810 0 66866 800
rect 67546 0 67602 800
rect 68282 0 68338 800
rect 69018 0 69074 800
rect 69754 0 69810 800
rect 70490 0 70546 800
rect 71226 0 71282 800
rect 71962 0 72018 800
rect 72698 0 72754 800
rect 73434 0 73490 800
rect 74170 0 74226 800
rect 74906 0 74962 800
rect 75642 0 75698 800
rect 76378 0 76434 800
rect 77114 0 77170 800
rect 77850 0 77906 800
rect 78586 0 78642 800
<< obsm2 >>
rect 682 84144 1250 84266
rect 1418 84144 1986 84266
rect 2154 84144 2722 84266
rect 2890 84144 3458 84266
rect 3626 84144 4194 84266
rect 4362 84144 4930 84266
rect 5098 84144 5666 84266
rect 5834 84144 6402 84266
rect 6570 84144 7138 84266
rect 7306 84144 7874 84266
rect 8042 84144 8610 84266
rect 8778 84144 9346 84266
rect 9514 84144 10082 84266
rect 10250 84144 10818 84266
rect 10986 84144 11554 84266
rect 11722 84144 12290 84266
rect 12458 84144 13026 84266
rect 13194 84144 13762 84266
rect 13930 84144 14498 84266
rect 14666 84144 15234 84266
rect 15402 84144 15970 84266
rect 16138 84144 16706 84266
rect 16874 84144 17442 84266
rect 17610 84144 18178 84266
rect 18346 84144 18914 84266
rect 19082 84144 19650 84266
rect 19818 84144 20386 84266
rect 20554 84144 21122 84266
rect 21290 84144 21858 84266
rect 22026 84144 22594 84266
rect 22762 84144 23330 84266
rect 23498 84144 24066 84266
rect 24234 84144 24802 84266
rect 24970 84144 25538 84266
rect 25706 84144 26274 84266
rect 26442 84144 27010 84266
rect 27178 84144 27746 84266
rect 27914 84144 28482 84266
rect 28650 84144 29218 84266
rect 29386 84144 29954 84266
rect 30122 84144 30690 84266
rect 30858 84144 31426 84266
rect 31594 84144 32162 84266
rect 32330 84144 32898 84266
rect 33066 84144 33634 84266
rect 33802 84144 34370 84266
rect 34538 84144 35106 84266
rect 35274 84144 35842 84266
rect 36010 84144 36578 84266
rect 36746 84144 37314 84266
rect 37482 84144 38050 84266
rect 38218 84144 38786 84266
rect 38954 84144 39522 84266
rect 39690 84144 40258 84266
rect 40426 84144 40994 84266
rect 41162 84144 41730 84266
rect 41898 84144 42466 84266
rect 42634 84144 43202 84266
rect 43370 84144 43938 84266
rect 44106 84144 44674 84266
rect 44842 84144 45410 84266
rect 45578 84144 46146 84266
rect 46314 84144 46882 84266
rect 47050 84144 47618 84266
rect 47786 84144 48354 84266
rect 48522 84144 49090 84266
rect 49258 84144 49826 84266
rect 49994 84144 50562 84266
rect 50730 84144 51298 84266
rect 51466 84144 52034 84266
rect 52202 84144 52770 84266
rect 52938 84144 53506 84266
rect 53674 84144 54242 84266
rect 54410 84144 54978 84266
rect 55146 84144 55714 84266
rect 55882 84144 56450 84266
rect 56618 84144 57186 84266
rect 57354 84144 57922 84266
rect 58090 84144 58658 84266
rect 58826 84144 59394 84266
rect 59562 84144 60130 84266
rect 60298 84144 60866 84266
rect 61034 84144 61602 84266
rect 61770 84144 62338 84266
rect 62506 84144 63074 84266
rect 63242 84144 63810 84266
rect 63978 84144 64546 84266
rect 64714 84144 65282 84266
rect 65450 84144 66018 84266
rect 66186 84144 66754 84266
rect 66922 84144 67490 84266
rect 67658 84144 68226 84266
rect 68394 84144 68962 84266
rect 69130 84144 69698 84266
rect 69866 84144 70434 84266
rect 70602 84144 71170 84266
rect 71338 84144 71906 84266
rect 72074 84144 72642 84266
rect 72810 84144 73378 84266
rect 73546 84144 74114 84266
rect 74282 84144 74850 84266
rect 75018 84144 75586 84266
rect 75754 84144 76322 84266
rect 76490 84144 77058 84266
rect 77226 84144 77794 84266
rect 77962 84144 78530 84266
rect 78698 84144 79266 84266
rect 79434 84144 79928 84266
rect 572 856 79928 84144
rect 572 70 1250 856
rect 1418 70 1986 856
rect 2154 70 2722 856
rect 2890 70 3458 856
rect 3626 70 4194 856
rect 4362 70 4930 856
rect 5098 70 5666 856
rect 5834 70 6402 856
rect 6570 70 7138 856
rect 7306 70 7874 856
rect 8042 70 8610 856
rect 8778 70 9346 856
rect 9514 70 10082 856
rect 10250 70 10818 856
rect 10986 70 11554 856
rect 11722 70 12290 856
rect 12458 70 13026 856
rect 13194 70 13762 856
rect 13930 70 14498 856
rect 14666 70 15234 856
rect 15402 70 15970 856
rect 16138 70 16706 856
rect 16874 70 17442 856
rect 17610 70 18178 856
rect 18346 70 18914 856
rect 19082 70 19650 856
rect 19818 70 20386 856
rect 20554 70 21122 856
rect 21290 70 21858 856
rect 22026 70 22594 856
rect 22762 70 23330 856
rect 23498 70 24066 856
rect 24234 70 24802 856
rect 24970 70 25538 856
rect 25706 70 26274 856
rect 26442 70 27010 856
rect 27178 70 27746 856
rect 27914 70 28482 856
rect 28650 70 29218 856
rect 29386 70 29954 856
rect 30122 70 30690 856
rect 30858 70 31426 856
rect 31594 70 32162 856
rect 32330 70 32898 856
rect 33066 70 33634 856
rect 33802 70 34370 856
rect 34538 70 35106 856
rect 35274 70 35842 856
rect 36010 70 36578 856
rect 36746 70 37314 856
rect 37482 70 38050 856
rect 38218 70 38786 856
rect 38954 70 39522 856
rect 39690 70 40258 856
rect 40426 70 40994 856
rect 41162 70 41730 856
rect 41898 70 42466 856
rect 42634 70 43202 856
rect 43370 70 43938 856
rect 44106 70 44674 856
rect 44842 70 45410 856
rect 45578 70 46146 856
rect 46314 70 46882 856
rect 47050 70 47618 856
rect 47786 70 48354 856
rect 48522 70 49090 856
rect 49258 70 49826 856
rect 49994 70 50562 856
rect 50730 70 51298 856
rect 51466 70 52034 856
rect 52202 70 52770 856
rect 52938 70 53506 856
rect 53674 70 54242 856
rect 54410 70 54978 856
rect 55146 70 55714 856
rect 55882 70 56450 856
rect 56618 70 57186 856
rect 57354 70 57922 856
rect 58090 70 58658 856
rect 58826 70 59394 856
rect 59562 70 60130 856
rect 60298 70 60866 856
rect 61034 70 61602 856
rect 61770 70 62338 856
rect 62506 70 63074 856
rect 63242 70 63810 856
rect 63978 70 64546 856
rect 64714 70 65282 856
rect 65450 70 66018 856
rect 66186 70 66754 856
rect 66922 70 67490 856
rect 67658 70 68226 856
rect 68394 70 68962 856
rect 69130 70 69698 856
rect 69866 70 70434 856
rect 70602 70 71170 856
rect 71338 70 71906 856
rect 72074 70 72642 856
rect 72810 70 73378 856
rect 73546 70 74114 856
rect 74282 70 74850 856
rect 75018 70 75586 856
rect 75754 70 76322 856
rect 76490 70 77058 856
rect 77226 70 77794 856
rect 77962 70 78530 856
rect 78698 70 79928 856
<< metal3 >>
rect 0 83104 800 83224
rect 0 81336 800 81456
rect 0 79568 800 79688
rect 0 77800 800 77920
rect 0 76032 800 76152
rect 0 74264 800 74384
rect 79200 73040 80000 73160
rect 79200 72768 80000 72888
rect 0 72496 800 72616
rect 79200 72496 80000 72616
rect 79200 72224 80000 72344
rect 79200 71952 80000 72072
rect 79200 71680 80000 71800
rect 79200 71408 80000 71528
rect 79200 71136 80000 71256
rect 0 70728 800 70848
rect 79200 70864 80000 70984
rect 79200 70592 80000 70712
rect 79200 70320 80000 70440
rect 79200 70048 80000 70168
rect 79200 69776 80000 69896
rect 79200 69504 80000 69624
rect 79200 69232 80000 69352
rect 0 68960 800 69080
rect 79200 68960 80000 69080
rect 79200 68688 80000 68808
rect 79200 68416 80000 68536
rect 79200 68144 80000 68264
rect 79200 67872 80000 67992
rect 79200 67600 80000 67720
rect 0 67192 800 67312
rect 79200 67328 80000 67448
rect 79200 67056 80000 67176
rect 79200 66784 80000 66904
rect 79200 66512 80000 66632
rect 79200 66240 80000 66360
rect 79200 65968 80000 66088
rect 79200 65696 80000 65816
rect 0 65424 800 65544
rect 79200 65424 80000 65544
rect 79200 65152 80000 65272
rect 79200 64880 80000 65000
rect 79200 64608 80000 64728
rect 79200 64336 80000 64456
rect 79200 64064 80000 64184
rect 0 63656 800 63776
rect 79200 63792 80000 63912
rect 79200 63520 80000 63640
rect 79200 63248 80000 63368
rect 79200 62976 80000 63096
rect 79200 62704 80000 62824
rect 79200 62432 80000 62552
rect 79200 62160 80000 62280
rect 0 61888 800 62008
rect 79200 61888 80000 62008
rect 79200 61616 80000 61736
rect 79200 61344 80000 61464
rect 79200 61072 80000 61192
rect 79200 60800 80000 60920
rect 79200 60528 80000 60648
rect 0 60120 800 60240
rect 79200 60256 80000 60376
rect 79200 59984 80000 60104
rect 79200 59712 80000 59832
rect 79200 59440 80000 59560
rect 79200 59168 80000 59288
rect 79200 58896 80000 59016
rect 79200 58624 80000 58744
rect 0 58352 800 58472
rect 79200 58352 80000 58472
rect 79200 58080 80000 58200
rect 79200 57808 80000 57928
rect 79200 57536 80000 57656
rect 79200 57264 80000 57384
rect 79200 56992 80000 57112
rect 0 56584 800 56704
rect 79200 56720 80000 56840
rect 79200 56448 80000 56568
rect 79200 56176 80000 56296
rect 79200 55904 80000 56024
rect 79200 55632 80000 55752
rect 79200 55360 80000 55480
rect 79200 55088 80000 55208
rect 0 54816 800 54936
rect 79200 54816 80000 54936
rect 79200 54544 80000 54664
rect 79200 54272 80000 54392
rect 79200 54000 80000 54120
rect 79200 53728 80000 53848
rect 79200 53456 80000 53576
rect 0 53048 800 53168
rect 79200 53184 80000 53304
rect 79200 52912 80000 53032
rect 79200 52640 80000 52760
rect 79200 52368 80000 52488
rect 79200 52096 80000 52216
rect 79200 51824 80000 51944
rect 79200 51552 80000 51672
rect 0 51280 800 51400
rect 79200 51280 80000 51400
rect 79200 51008 80000 51128
rect 79200 50736 80000 50856
rect 79200 50464 80000 50584
rect 79200 50192 80000 50312
rect 79200 49920 80000 50040
rect 0 49512 800 49632
rect 79200 49648 80000 49768
rect 79200 49376 80000 49496
rect 79200 49104 80000 49224
rect 79200 48832 80000 48952
rect 79200 48560 80000 48680
rect 79200 48288 80000 48408
rect 79200 48016 80000 48136
rect 0 47744 800 47864
rect 79200 47744 80000 47864
rect 79200 47472 80000 47592
rect 79200 47200 80000 47320
rect 79200 46928 80000 47048
rect 79200 46656 80000 46776
rect 79200 46384 80000 46504
rect 0 45976 800 46096
rect 79200 46112 80000 46232
rect 79200 45840 80000 45960
rect 79200 45568 80000 45688
rect 79200 45296 80000 45416
rect 79200 45024 80000 45144
rect 79200 44752 80000 44872
rect 79200 44480 80000 44600
rect 0 44208 800 44328
rect 79200 44208 80000 44328
rect 79200 43936 80000 44056
rect 79200 43664 80000 43784
rect 79200 43392 80000 43512
rect 79200 43120 80000 43240
rect 79200 42848 80000 42968
rect 0 42440 800 42560
rect 79200 42576 80000 42696
rect 79200 42304 80000 42424
rect 79200 42032 80000 42152
rect 79200 41760 80000 41880
rect 79200 41488 80000 41608
rect 79200 41216 80000 41336
rect 79200 40944 80000 41064
rect 0 40672 800 40792
rect 79200 40672 80000 40792
rect 79200 40400 80000 40520
rect 79200 40128 80000 40248
rect 79200 39856 80000 39976
rect 79200 39584 80000 39704
rect 79200 39312 80000 39432
rect 0 38904 800 39024
rect 79200 39040 80000 39160
rect 79200 38768 80000 38888
rect 79200 38496 80000 38616
rect 79200 38224 80000 38344
rect 79200 37952 80000 38072
rect 79200 37680 80000 37800
rect 79200 37408 80000 37528
rect 0 37136 800 37256
rect 79200 37136 80000 37256
rect 79200 36864 80000 36984
rect 79200 36592 80000 36712
rect 79200 36320 80000 36440
rect 79200 36048 80000 36168
rect 79200 35776 80000 35896
rect 0 35368 800 35488
rect 79200 35504 80000 35624
rect 79200 35232 80000 35352
rect 79200 34960 80000 35080
rect 79200 34688 80000 34808
rect 79200 34416 80000 34536
rect 79200 34144 80000 34264
rect 79200 33872 80000 33992
rect 0 33600 800 33720
rect 79200 33600 80000 33720
rect 79200 33328 80000 33448
rect 79200 33056 80000 33176
rect 79200 32784 80000 32904
rect 79200 32512 80000 32632
rect 79200 32240 80000 32360
rect 0 31832 800 31952
rect 79200 31968 80000 32088
rect 79200 31696 80000 31816
rect 79200 31424 80000 31544
rect 79200 31152 80000 31272
rect 79200 30880 80000 31000
rect 79200 30608 80000 30728
rect 79200 30336 80000 30456
rect 0 30064 800 30184
rect 79200 30064 80000 30184
rect 79200 29792 80000 29912
rect 79200 29520 80000 29640
rect 79200 29248 80000 29368
rect 79200 28976 80000 29096
rect 79200 28704 80000 28824
rect 0 28296 800 28416
rect 79200 28432 80000 28552
rect 79200 28160 80000 28280
rect 79200 27888 80000 28008
rect 79200 27616 80000 27736
rect 79200 27344 80000 27464
rect 79200 27072 80000 27192
rect 79200 26800 80000 26920
rect 0 26528 800 26648
rect 79200 26528 80000 26648
rect 79200 26256 80000 26376
rect 79200 25984 80000 26104
rect 79200 25712 80000 25832
rect 79200 25440 80000 25560
rect 79200 25168 80000 25288
rect 0 24760 800 24880
rect 79200 24896 80000 25016
rect 79200 24624 80000 24744
rect 79200 24352 80000 24472
rect 79200 24080 80000 24200
rect 79200 23808 80000 23928
rect 79200 23536 80000 23656
rect 79200 23264 80000 23384
rect 0 22992 800 23112
rect 79200 22992 80000 23112
rect 79200 22720 80000 22840
rect 79200 22448 80000 22568
rect 79200 22176 80000 22296
rect 79200 21904 80000 22024
rect 79200 21632 80000 21752
rect 0 21224 800 21344
rect 79200 21360 80000 21480
rect 79200 21088 80000 21208
rect 79200 20816 80000 20936
rect 79200 20544 80000 20664
rect 79200 20272 80000 20392
rect 79200 20000 80000 20120
rect 79200 19728 80000 19848
rect 0 19456 800 19576
rect 79200 19456 80000 19576
rect 79200 19184 80000 19304
rect 79200 18912 80000 19032
rect 79200 18640 80000 18760
rect 79200 18368 80000 18488
rect 79200 18096 80000 18216
rect 0 17688 800 17808
rect 79200 17824 80000 17944
rect 79200 17552 80000 17672
rect 79200 17280 80000 17400
rect 79200 17008 80000 17128
rect 79200 16736 80000 16856
rect 79200 16464 80000 16584
rect 79200 16192 80000 16312
rect 0 15920 800 16040
rect 79200 15920 80000 16040
rect 79200 15648 80000 15768
rect 79200 15376 80000 15496
rect 79200 15104 80000 15224
rect 79200 14832 80000 14952
rect 79200 14560 80000 14680
rect 0 14152 800 14272
rect 79200 14288 80000 14408
rect 79200 14016 80000 14136
rect 79200 13744 80000 13864
rect 79200 13472 80000 13592
rect 79200 13200 80000 13320
rect 79200 12928 80000 13048
rect 79200 12656 80000 12776
rect 0 12384 800 12504
rect 79200 12384 80000 12504
rect 79200 12112 80000 12232
rect 79200 11840 80000 11960
rect 0 10616 800 10736
rect 0 8848 800 8968
rect 0 7080 800 7200
rect 0 5312 800 5432
rect 0 3544 800 3664
rect 0 1776 800 1896
<< obsm3 >>
rect 880 83024 79200 83197
rect 800 81536 79200 83024
rect 880 81256 79200 81536
rect 800 79768 79200 81256
rect 880 79488 79200 79768
rect 800 78000 79200 79488
rect 880 77720 79200 78000
rect 800 76232 79200 77720
rect 880 75952 79200 76232
rect 800 74464 79200 75952
rect 880 74184 79200 74464
rect 800 73240 79200 74184
rect 800 72696 79120 73240
rect 880 72416 79120 72696
rect 800 70928 79120 72416
rect 880 70648 79120 70928
rect 800 69160 79120 70648
rect 880 68880 79120 69160
rect 800 67392 79120 68880
rect 880 67112 79120 67392
rect 800 65624 79120 67112
rect 880 65344 79120 65624
rect 800 63856 79120 65344
rect 880 63576 79120 63856
rect 800 62088 79120 63576
rect 880 61808 79120 62088
rect 800 60320 79120 61808
rect 880 60040 79120 60320
rect 800 58552 79120 60040
rect 880 58272 79120 58552
rect 800 56784 79120 58272
rect 880 56504 79120 56784
rect 800 55016 79120 56504
rect 880 54736 79120 55016
rect 800 53248 79120 54736
rect 880 52968 79120 53248
rect 800 51480 79120 52968
rect 880 51200 79120 51480
rect 800 49712 79120 51200
rect 880 49432 79120 49712
rect 800 47944 79120 49432
rect 880 47664 79120 47944
rect 800 46176 79120 47664
rect 880 45896 79120 46176
rect 800 44408 79120 45896
rect 880 44128 79120 44408
rect 800 42640 79120 44128
rect 880 42360 79120 42640
rect 800 40872 79120 42360
rect 880 40592 79120 40872
rect 800 39104 79120 40592
rect 880 38824 79120 39104
rect 800 37336 79120 38824
rect 880 37056 79120 37336
rect 800 35568 79120 37056
rect 880 35288 79120 35568
rect 800 33800 79120 35288
rect 880 33520 79120 33800
rect 800 32032 79120 33520
rect 880 31752 79120 32032
rect 800 30264 79120 31752
rect 880 29984 79120 30264
rect 800 28496 79120 29984
rect 880 28216 79120 28496
rect 800 26728 79120 28216
rect 880 26448 79120 26728
rect 800 24960 79120 26448
rect 880 24680 79120 24960
rect 800 23192 79120 24680
rect 880 22912 79120 23192
rect 800 21424 79120 22912
rect 880 21144 79120 21424
rect 800 19656 79120 21144
rect 880 19376 79120 19656
rect 800 17888 79120 19376
rect 880 17608 79120 17888
rect 800 16120 79120 17608
rect 880 15840 79120 16120
rect 800 14352 79120 15840
rect 880 14072 79120 14352
rect 800 12584 79120 14072
rect 880 12304 79120 12584
rect 800 11760 79120 12304
rect 800 10816 79200 11760
rect 880 10536 79200 10816
rect 800 9048 79200 10536
rect 880 8768 79200 9048
rect 800 7280 79200 8768
rect 880 7000 79200 7280
rect 800 5512 79200 7000
rect 880 5232 79200 5512
rect 800 3744 79200 5232
rect 880 3464 79200 3744
rect 800 1976 79200 3464
rect 880 1803 79200 1976
<< metal4 >>
rect 4208 2128 4528 82736
rect 19568 2128 19888 82736
rect 34928 2128 35248 82736
rect 50288 2128 50608 82736
rect 65648 2128 65968 82736
<< obsm4 >>
rect 1715 2347 4128 81565
rect 4608 2347 19488 81565
rect 19968 2347 34848 81565
rect 35328 2347 50208 81565
rect 50688 2347 65568 81565
rect 66048 2347 77037 81565
<< labels >>
rlabel metal2 s 77114 84200 77170 85000 6 caravel_irq[0]
port 1 nsew signal output
rlabel metal2 s 77850 84200 77906 85000 6 caravel_irq[1]
port 2 nsew signal output
rlabel metal2 s 78586 84200 78642 85000 6 caravel_irq[2]
port 3 nsew signal output
rlabel metal2 s 79322 84200 79378 85000 6 caravel_irq[3]
port 4 nsew signal output
rlabel metal2 s 75642 84200 75698 85000 6 caravel_uart_rx
port 5 nsew signal input
rlabel metal2 s 76378 84200 76434 85000 6 caravel_uart_tx
port 6 nsew signal output
rlabel metal2 s 570 84200 626 85000 6 caravel_wb_ack_i
port 7 nsew signal input
rlabel metal2 s 4986 84200 5042 85000 6 caravel_wb_adr_o[0]
port 8 nsew signal output
rlabel metal2 s 30010 84200 30066 85000 6 caravel_wb_adr_o[10]
port 9 nsew signal output
rlabel metal2 s 32218 84200 32274 85000 6 caravel_wb_adr_o[11]
port 10 nsew signal output
rlabel metal2 s 34426 84200 34482 85000 6 caravel_wb_adr_o[12]
port 11 nsew signal output
rlabel metal2 s 36634 84200 36690 85000 6 caravel_wb_adr_o[13]
port 12 nsew signal output
rlabel metal2 s 38842 84200 38898 85000 6 caravel_wb_adr_o[14]
port 13 nsew signal output
rlabel metal2 s 41050 84200 41106 85000 6 caravel_wb_adr_o[15]
port 14 nsew signal output
rlabel metal2 s 43258 84200 43314 85000 6 caravel_wb_adr_o[16]
port 15 nsew signal output
rlabel metal2 s 45466 84200 45522 85000 6 caravel_wb_adr_o[17]
port 16 nsew signal output
rlabel metal2 s 47674 84200 47730 85000 6 caravel_wb_adr_o[18]
port 17 nsew signal output
rlabel metal2 s 49882 84200 49938 85000 6 caravel_wb_adr_o[19]
port 18 nsew signal output
rlabel metal2 s 7930 84200 7986 85000 6 caravel_wb_adr_o[1]
port 19 nsew signal output
rlabel metal2 s 52090 84200 52146 85000 6 caravel_wb_adr_o[20]
port 20 nsew signal output
rlabel metal2 s 54298 84200 54354 85000 6 caravel_wb_adr_o[21]
port 21 nsew signal output
rlabel metal2 s 56506 84200 56562 85000 6 caravel_wb_adr_o[22]
port 22 nsew signal output
rlabel metal2 s 58714 84200 58770 85000 6 caravel_wb_adr_o[23]
port 23 nsew signal output
rlabel metal2 s 60922 84200 60978 85000 6 caravel_wb_adr_o[24]
port 24 nsew signal output
rlabel metal2 s 63130 84200 63186 85000 6 caravel_wb_adr_o[25]
port 25 nsew signal output
rlabel metal2 s 65338 84200 65394 85000 6 caravel_wb_adr_o[26]
port 26 nsew signal output
rlabel metal2 s 67546 84200 67602 85000 6 caravel_wb_adr_o[27]
port 27 nsew signal output
rlabel metal2 s 10874 84200 10930 85000 6 caravel_wb_adr_o[2]
port 28 nsew signal output
rlabel metal2 s 13818 84200 13874 85000 6 caravel_wb_adr_o[3]
port 29 nsew signal output
rlabel metal2 s 16762 84200 16818 85000 6 caravel_wb_adr_o[4]
port 30 nsew signal output
rlabel metal2 s 18970 84200 19026 85000 6 caravel_wb_adr_o[5]
port 31 nsew signal output
rlabel metal2 s 21178 84200 21234 85000 6 caravel_wb_adr_o[6]
port 32 nsew signal output
rlabel metal2 s 23386 84200 23442 85000 6 caravel_wb_adr_o[7]
port 33 nsew signal output
rlabel metal2 s 25594 84200 25650 85000 6 caravel_wb_adr_o[8]
port 34 nsew signal output
rlabel metal2 s 27802 84200 27858 85000 6 caravel_wb_adr_o[9]
port 35 nsew signal output
rlabel metal2 s 1306 84200 1362 85000 6 caravel_wb_cyc_o
port 36 nsew signal output
rlabel metal2 s 5722 84200 5778 85000 6 caravel_wb_data_i[0]
port 37 nsew signal input
rlabel metal2 s 30746 84200 30802 85000 6 caravel_wb_data_i[10]
port 38 nsew signal input
rlabel metal2 s 32954 84200 33010 85000 6 caravel_wb_data_i[11]
port 39 nsew signal input
rlabel metal2 s 35162 84200 35218 85000 6 caravel_wb_data_i[12]
port 40 nsew signal input
rlabel metal2 s 37370 84200 37426 85000 6 caravel_wb_data_i[13]
port 41 nsew signal input
rlabel metal2 s 39578 84200 39634 85000 6 caravel_wb_data_i[14]
port 42 nsew signal input
rlabel metal2 s 41786 84200 41842 85000 6 caravel_wb_data_i[15]
port 43 nsew signal input
rlabel metal2 s 43994 84200 44050 85000 6 caravel_wb_data_i[16]
port 44 nsew signal input
rlabel metal2 s 46202 84200 46258 85000 6 caravel_wb_data_i[17]
port 45 nsew signal input
rlabel metal2 s 48410 84200 48466 85000 6 caravel_wb_data_i[18]
port 46 nsew signal input
rlabel metal2 s 50618 84200 50674 85000 6 caravel_wb_data_i[19]
port 47 nsew signal input
rlabel metal2 s 8666 84200 8722 85000 6 caravel_wb_data_i[1]
port 48 nsew signal input
rlabel metal2 s 52826 84200 52882 85000 6 caravel_wb_data_i[20]
port 49 nsew signal input
rlabel metal2 s 55034 84200 55090 85000 6 caravel_wb_data_i[21]
port 50 nsew signal input
rlabel metal2 s 57242 84200 57298 85000 6 caravel_wb_data_i[22]
port 51 nsew signal input
rlabel metal2 s 59450 84200 59506 85000 6 caravel_wb_data_i[23]
port 52 nsew signal input
rlabel metal2 s 61658 84200 61714 85000 6 caravel_wb_data_i[24]
port 53 nsew signal input
rlabel metal2 s 63866 84200 63922 85000 6 caravel_wb_data_i[25]
port 54 nsew signal input
rlabel metal2 s 66074 84200 66130 85000 6 caravel_wb_data_i[26]
port 55 nsew signal input
rlabel metal2 s 68282 84200 68338 85000 6 caravel_wb_data_i[27]
port 56 nsew signal input
rlabel metal2 s 69754 84200 69810 85000 6 caravel_wb_data_i[28]
port 57 nsew signal input
rlabel metal2 s 71226 84200 71282 85000 6 caravel_wb_data_i[29]
port 58 nsew signal input
rlabel metal2 s 11610 84200 11666 85000 6 caravel_wb_data_i[2]
port 59 nsew signal input
rlabel metal2 s 72698 84200 72754 85000 6 caravel_wb_data_i[30]
port 60 nsew signal input
rlabel metal2 s 74170 84200 74226 85000 6 caravel_wb_data_i[31]
port 61 nsew signal input
rlabel metal2 s 14554 84200 14610 85000 6 caravel_wb_data_i[3]
port 62 nsew signal input
rlabel metal2 s 17498 84200 17554 85000 6 caravel_wb_data_i[4]
port 63 nsew signal input
rlabel metal2 s 19706 84200 19762 85000 6 caravel_wb_data_i[5]
port 64 nsew signal input
rlabel metal2 s 21914 84200 21970 85000 6 caravel_wb_data_i[6]
port 65 nsew signal input
rlabel metal2 s 24122 84200 24178 85000 6 caravel_wb_data_i[7]
port 66 nsew signal input
rlabel metal2 s 26330 84200 26386 85000 6 caravel_wb_data_i[8]
port 67 nsew signal input
rlabel metal2 s 28538 84200 28594 85000 6 caravel_wb_data_i[9]
port 68 nsew signal input
rlabel metal2 s 6458 84200 6514 85000 6 caravel_wb_data_o[0]
port 69 nsew signal output
rlabel metal2 s 31482 84200 31538 85000 6 caravel_wb_data_o[10]
port 70 nsew signal output
rlabel metal2 s 33690 84200 33746 85000 6 caravel_wb_data_o[11]
port 71 nsew signal output
rlabel metal2 s 35898 84200 35954 85000 6 caravel_wb_data_o[12]
port 72 nsew signal output
rlabel metal2 s 38106 84200 38162 85000 6 caravel_wb_data_o[13]
port 73 nsew signal output
rlabel metal2 s 40314 84200 40370 85000 6 caravel_wb_data_o[14]
port 74 nsew signal output
rlabel metal2 s 42522 84200 42578 85000 6 caravel_wb_data_o[15]
port 75 nsew signal output
rlabel metal2 s 44730 84200 44786 85000 6 caravel_wb_data_o[16]
port 76 nsew signal output
rlabel metal2 s 46938 84200 46994 85000 6 caravel_wb_data_o[17]
port 77 nsew signal output
rlabel metal2 s 49146 84200 49202 85000 6 caravel_wb_data_o[18]
port 78 nsew signal output
rlabel metal2 s 51354 84200 51410 85000 6 caravel_wb_data_o[19]
port 79 nsew signal output
rlabel metal2 s 9402 84200 9458 85000 6 caravel_wb_data_o[1]
port 80 nsew signal output
rlabel metal2 s 53562 84200 53618 85000 6 caravel_wb_data_o[20]
port 81 nsew signal output
rlabel metal2 s 55770 84200 55826 85000 6 caravel_wb_data_o[21]
port 82 nsew signal output
rlabel metal2 s 57978 84200 58034 85000 6 caravel_wb_data_o[22]
port 83 nsew signal output
rlabel metal2 s 60186 84200 60242 85000 6 caravel_wb_data_o[23]
port 84 nsew signal output
rlabel metal2 s 62394 84200 62450 85000 6 caravel_wb_data_o[24]
port 85 nsew signal output
rlabel metal2 s 64602 84200 64658 85000 6 caravel_wb_data_o[25]
port 86 nsew signal output
rlabel metal2 s 66810 84200 66866 85000 6 caravel_wb_data_o[26]
port 87 nsew signal output
rlabel metal2 s 69018 84200 69074 85000 6 caravel_wb_data_o[27]
port 88 nsew signal output
rlabel metal2 s 70490 84200 70546 85000 6 caravel_wb_data_o[28]
port 89 nsew signal output
rlabel metal2 s 71962 84200 72018 85000 6 caravel_wb_data_o[29]
port 90 nsew signal output
rlabel metal2 s 12346 84200 12402 85000 6 caravel_wb_data_o[2]
port 91 nsew signal output
rlabel metal2 s 73434 84200 73490 85000 6 caravel_wb_data_o[30]
port 92 nsew signal output
rlabel metal2 s 74906 84200 74962 85000 6 caravel_wb_data_o[31]
port 93 nsew signal output
rlabel metal2 s 15290 84200 15346 85000 6 caravel_wb_data_o[3]
port 94 nsew signal output
rlabel metal2 s 18234 84200 18290 85000 6 caravel_wb_data_o[4]
port 95 nsew signal output
rlabel metal2 s 20442 84200 20498 85000 6 caravel_wb_data_o[5]
port 96 nsew signal output
rlabel metal2 s 22650 84200 22706 85000 6 caravel_wb_data_o[6]
port 97 nsew signal output
rlabel metal2 s 24858 84200 24914 85000 6 caravel_wb_data_o[7]
port 98 nsew signal output
rlabel metal2 s 27066 84200 27122 85000 6 caravel_wb_data_o[8]
port 99 nsew signal output
rlabel metal2 s 29274 84200 29330 85000 6 caravel_wb_data_o[9]
port 100 nsew signal output
rlabel metal2 s 2042 84200 2098 85000 6 caravel_wb_error_i
port 101 nsew signal input
rlabel metal2 s 7194 84200 7250 85000 6 caravel_wb_sel_o[0]
port 102 nsew signal output
rlabel metal2 s 10138 84200 10194 85000 6 caravel_wb_sel_o[1]
port 103 nsew signal output
rlabel metal2 s 13082 84200 13138 85000 6 caravel_wb_sel_o[2]
port 104 nsew signal output
rlabel metal2 s 16026 84200 16082 85000 6 caravel_wb_sel_o[3]
port 105 nsew signal output
rlabel metal2 s 2778 84200 2834 85000 6 caravel_wb_stall_i
port 106 nsew signal input
rlabel metal2 s 3514 84200 3570 85000 6 caravel_wb_stb_o
port 107 nsew signal output
rlabel metal2 s 4250 84200 4306 85000 6 caravel_wb_we_o
port 108 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 core0Index[0]
port 109 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 core0Index[1]
port 110 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 core0Index[2]
port 111 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 core0Index[3]
port 112 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 core0Index[4]
port 113 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 core0Index[5]
port 114 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 core0Index[6]
port 115 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 core0Index[7]
port 116 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 core1Index[0]
port 117 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 core1Index[1]
port 118 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 core1Index[2]
port 119 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 core1Index[3]
port 120 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 core1Index[4]
port 121 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 core1Index[5]
port 122 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 core1Index[6]
port 123 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 core1Index[7]
port 124 nsew signal output
rlabel metal3 s 79200 11840 80000 11960 6 la_data_out[0]
port 125 nsew signal output
rlabel metal3 s 79200 39040 80000 39160 6 la_data_out[100]
port 126 nsew signal output
rlabel metal3 s 79200 39312 80000 39432 6 la_data_out[101]
port 127 nsew signal output
rlabel metal3 s 79200 39584 80000 39704 6 la_data_out[102]
port 128 nsew signal output
rlabel metal3 s 79200 39856 80000 39976 6 la_data_out[103]
port 129 nsew signal output
rlabel metal3 s 79200 40128 80000 40248 6 la_data_out[104]
port 130 nsew signal output
rlabel metal3 s 79200 40400 80000 40520 6 la_data_out[105]
port 131 nsew signal output
rlabel metal3 s 79200 40672 80000 40792 6 la_data_out[106]
port 132 nsew signal output
rlabel metal3 s 79200 40944 80000 41064 6 la_data_out[107]
port 133 nsew signal output
rlabel metal3 s 79200 41216 80000 41336 6 la_data_out[108]
port 134 nsew signal output
rlabel metal3 s 79200 41488 80000 41608 6 la_data_out[109]
port 135 nsew signal output
rlabel metal3 s 79200 14560 80000 14680 6 la_data_out[10]
port 136 nsew signal output
rlabel metal3 s 79200 41760 80000 41880 6 la_data_out[110]
port 137 nsew signal output
rlabel metal3 s 79200 42032 80000 42152 6 la_data_out[111]
port 138 nsew signal output
rlabel metal3 s 79200 42304 80000 42424 6 la_data_out[112]
port 139 nsew signal output
rlabel metal3 s 79200 42576 80000 42696 6 la_data_out[113]
port 140 nsew signal output
rlabel metal3 s 79200 42848 80000 42968 6 la_data_out[114]
port 141 nsew signal output
rlabel metal3 s 79200 43120 80000 43240 6 la_data_out[115]
port 142 nsew signal output
rlabel metal3 s 79200 43392 80000 43512 6 la_data_out[116]
port 143 nsew signal output
rlabel metal3 s 79200 43664 80000 43784 6 la_data_out[117]
port 144 nsew signal output
rlabel metal3 s 79200 43936 80000 44056 6 la_data_out[118]
port 145 nsew signal output
rlabel metal3 s 79200 44208 80000 44328 6 la_data_out[119]
port 146 nsew signal output
rlabel metal3 s 79200 14832 80000 14952 6 la_data_out[11]
port 147 nsew signal output
rlabel metal3 s 79200 44480 80000 44600 6 la_data_out[120]
port 148 nsew signal output
rlabel metal3 s 79200 44752 80000 44872 6 la_data_out[121]
port 149 nsew signal output
rlabel metal3 s 79200 45024 80000 45144 6 la_data_out[122]
port 150 nsew signal output
rlabel metal3 s 79200 45296 80000 45416 6 la_data_out[123]
port 151 nsew signal output
rlabel metal3 s 79200 45568 80000 45688 6 la_data_out[124]
port 152 nsew signal output
rlabel metal3 s 79200 45840 80000 45960 6 la_data_out[125]
port 153 nsew signal output
rlabel metal3 s 79200 46112 80000 46232 6 la_data_out[126]
port 154 nsew signal output
rlabel metal3 s 79200 46384 80000 46504 6 la_data_out[127]
port 155 nsew signal output
rlabel metal3 s 79200 15104 80000 15224 6 la_data_out[12]
port 156 nsew signal output
rlabel metal3 s 79200 15376 80000 15496 6 la_data_out[13]
port 157 nsew signal output
rlabel metal3 s 79200 15648 80000 15768 6 la_data_out[14]
port 158 nsew signal output
rlabel metal3 s 79200 15920 80000 16040 6 la_data_out[15]
port 159 nsew signal output
rlabel metal3 s 79200 16192 80000 16312 6 la_data_out[16]
port 160 nsew signal output
rlabel metal3 s 79200 16464 80000 16584 6 la_data_out[17]
port 161 nsew signal output
rlabel metal3 s 79200 16736 80000 16856 6 la_data_out[18]
port 162 nsew signal output
rlabel metal3 s 79200 17008 80000 17128 6 la_data_out[19]
port 163 nsew signal output
rlabel metal3 s 79200 12112 80000 12232 6 la_data_out[1]
port 164 nsew signal output
rlabel metal3 s 79200 17280 80000 17400 6 la_data_out[20]
port 165 nsew signal output
rlabel metal3 s 79200 17552 80000 17672 6 la_data_out[21]
port 166 nsew signal output
rlabel metal3 s 79200 17824 80000 17944 6 la_data_out[22]
port 167 nsew signal output
rlabel metal3 s 79200 18096 80000 18216 6 la_data_out[23]
port 168 nsew signal output
rlabel metal3 s 79200 18368 80000 18488 6 la_data_out[24]
port 169 nsew signal output
rlabel metal3 s 79200 18640 80000 18760 6 la_data_out[25]
port 170 nsew signal output
rlabel metal3 s 79200 18912 80000 19032 6 la_data_out[26]
port 171 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 la_data_out[27]
port 172 nsew signal output
rlabel metal3 s 79200 19456 80000 19576 6 la_data_out[28]
port 173 nsew signal output
rlabel metal3 s 79200 19728 80000 19848 6 la_data_out[29]
port 174 nsew signal output
rlabel metal3 s 79200 12384 80000 12504 6 la_data_out[2]
port 175 nsew signal output
rlabel metal3 s 79200 20000 80000 20120 6 la_data_out[30]
port 176 nsew signal output
rlabel metal3 s 79200 20272 80000 20392 6 la_data_out[31]
port 177 nsew signal output
rlabel metal3 s 79200 20544 80000 20664 6 la_data_out[32]
port 178 nsew signal output
rlabel metal3 s 79200 20816 80000 20936 6 la_data_out[33]
port 179 nsew signal output
rlabel metal3 s 79200 21088 80000 21208 6 la_data_out[34]
port 180 nsew signal output
rlabel metal3 s 79200 21360 80000 21480 6 la_data_out[35]
port 181 nsew signal output
rlabel metal3 s 79200 21632 80000 21752 6 la_data_out[36]
port 182 nsew signal output
rlabel metal3 s 79200 21904 80000 22024 6 la_data_out[37]
port 183 nsew signal output
rlabel metal3 s 79200 22176 80000 22296 6 la_data_out[38]
port 184 nsew signal output
rlabel metal3 s 79200 22448 80000 22568 6 la_data_out[39]
port 185 nsew signal output
rlabel metal3 s 79200 12656 80000 12776 6 la_data_out[3]
port 186 nsew signal output
rlabel metal3 s 79200 22720 80000 22840 6 la_data_out[40]
port 187 nsew signal output
rlabel metal3 s 79200 22992 80000 23112 6 la_data_out[41]
port 188 nsew signal output
rlabel metal3 s 79200 23264 80000 23384 6 la_data_out[42]
port 189 nsew signal output
rlabel metal3 s 79200 23536 80000 23656 6 la_data_out[43]
port 190 nsew signal output
rlabel metal3 s 79200 23808 80000 23928 6 la_data_out[44]
port 191 nsew signal output
rlabel metal3 s 79200 24080 80000 24200 6 la_data_out[45]
port 192 nsew signal output
rlabel metal3 s 79200 24352 80000 24472 6 la_data_out[46]
port 193 nsew signal output
rlabel metal3 s 79200 24624 80000 24744 6 la_data_out[47]
port 194 nsew signal output
rlabel metal3 s 79200 24896 80000 25016 6 la_data_out[48]
port 195 nsew signal output
rlabel metal3 s 79200 25168 80000 25288 6 la_data_out[49]
port 196 nsew signal output
rlabel metal3 s 79200 12928 80000 13048 6 la_data_out[4]
port 197 nsew signal output
rlabel metal3 s 79200 25440 80000 25560 6 la_data_out[50]
port 198 nsew signal output
rlabel metal3 s 79200 25712 80000 25832 6 la_data_out[51]
port 199 nsew signal output
rlabel metal3 s 79200 25984 80000 26104 6 la_data_out[52]
port 200 nsew signal output
rlabel metal3 s 79200 26256 80000 26376 6 la_data_out[53]
port 201 nsew signal output
rlabel metal3 s 79200 26528 80000 26648 6 la_data_out[54]
port 202 nsew signal output
rlabel metal3 s 79200 26800 80000 26920 6 la_data_out[55]
port 203 nsew signal output
rlabel metal3 s 79200 27072 80000 27192 6 la_data_out[56]
port 204 nsew signal output
rlabel metal3 s 79200 27344 80000 27464 6 la_data_out[57]
port 205 nsew signal output
rlabel metal3 s 79200 27616 80000 27736 6 la_data_out[58]
port 206 nsew signal output
rlabel metal3 s 79200 27888 80000 28008 6 la_data_out[59]
port 207 nsew signal output
rlabel metal3 s 79200 13200 80000 13320 6 la_data_out[5]
port 208 nsew signal output
rlabel metal3 s 79200 28160 80000 28280 6 la_data_out[60]
port 209 nsew signal output
rlabel metal3 s 79200 28432 80000 28552 6 la_data_out[61]
port 210 nsew signal output
rlabel metal3 s 79200 28704 80000 28824 6 la_data_out[62]
port 211 nsew signal output
rlabel metal3 s 79200 28976 80000 29096 6 la_data_out[63]
port 212 nsew signal output
rlabel metal3 s 79200 29248 80000 29368 6 la_data_out[64]
port 213 nsew signal output
rlabel metal3 s 79200 29520 80000 29640 6 la_data_out[65]
port 214 nsew signal output
rlabel metal3 s 79200 29792 80000 29912 6 la_data_out[66]
port 215 nsew signal output
rlabel metal3 s 79200 30064 80000 30184 6 la_data_out[67]
port 216 nsew signal output
rlabel metal3 s 79200 30336 80000 30456 6 la_data_out[68]
port 217 nsew signal output
rlabel metal3 s 79200 30608 80000 30728 6 la_data_out[69]
port 218 nsew signal output
rlabel metal3 s 79200 13472 80000 13592 6 la_data_out[6]
port 219 nsew signal output
rlabel metal3 s 79200 30880 80000 31000 6 la_data_out[70]
port 220 nsew signal output
rlabel metal3 s 79200 31152 80000 31272 6 la_data_out[71]
port 221 nsew signal output
rlabel metal3 s 79200 31424 80000 31544 6 la_data_out[72]
port 222 nsew signal output
rlabel metal3 s 79200 31696 80000 31816 6 la_data_out[73]
port 223 nsew signal output
rlabel metal3 s 79200 31968 80000 32088 6 la_data_out[74]
port 224 nsew signal output
rlabel metal3 s 79200 32240 80000 32360 6 la_data_out[75]
port 225 nsew signal output
rlabel metal3 s 79200 32512 80000 32632 6 la_data_out[76]
port 226 nsew signal output
rlabel metal3 s 79200 32784 80000 32904 6 la_data_out[77]
port 227 nsew signal output
rlabel metal3 s 79200 33056 80000 33176 6 la_data_out[78]
port 228 nsew signal output
rlabel metal3 s 79200 33328 80000 33448 6 la_data_out[79]
port 229 nsew signal output
rlabel metal3 s 79200 13744 80000 13864 6 la_data_out[7]
port 230 nsew signal output
rlabel metal3 s 79200 33600 80000 33720 6 la_data_out[80]
port 231 nsew signal output
rlabel metal3 s 79200 33872 80000 33992 6 la_data_out[81]
port 232 nsew signal output
rlabel metal3 s 79200 34144 80000 34264 6 la_data_out[82]
port 233 nsew signal output
rlabel metal3 s 79200 34416 80000 34536 6 la_data_out[83]
port 234 nsew signal output
rlabel metal3 s 79200 34688 80000 34808 6 la_data_out[84]
port 235 nsew signal output
rlabel metal3 s 79200 34960 80000 35080 6 la_data_out[85]
port 236 nsew signal output
rlabel metal3 s 79200 35232 80000 35352 6 la_data_out[86]
port 237 nsew signal output
rlabel metal3 s 79200 35504 80000 35624 6 la_data_out[87]
port 238 nsew signal output
rlabel metal3 s 79200 35776 80000 35896 6 la_data_out[88]
port 239 nsew signal output
rlabel metal3 s 79200 36048 80000 36168 6 la_data_out[89]
port 240 nsew signal output
rlabel metal3 s 79200 14016 80000 14136 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 79200 36320 80000 36440 6 la_data_out[90]
port 242 nsew signal output
rlabel metal3 s 79200 36592 80000 36712 6 la_data_out[91]
port 243 nsew signal output
rlabel metal3 s 79200 36864 80000 36984 6 la_data_out[92]
port 244 nsew signal output
rlabel metal3 s 79200 37136 80000 37256 6 la_data_out[93]
port 245 nsew signal output
rlabel metal3 s 79200 37408 80000 37528 6 la_data_out[94]
port 246 nsew signal output
rlabel metal3 s 79200 37680 80000 37800 6 la_data_out[95]
port 247 nsew signal output
rlabel metal3 s 79200 37952 80000 38072 6 la_data_out[96]
port 248 nsew signal output
rlabel metal3 s 79200 38224 80000 38344 6 la_data_out[97]
port 249 nsew signal output
rlabel metal3 s 79200 38496 80000 38616 6 la_data_out[98]
port 250 nsew signal output
rlabel metal3 s 79200 38768 80000 38888 6 la_data_out[99]
port 251 nsew signal output
rlabel metal3 s 79200 14288 80000 14408 6 la_data_out[9]
port 252 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 manufacturerID[0]
port 253 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 manufacturerID[10]
port 254 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 manufacturerID[1]
port 255 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 manufacturerID[2]
port 256 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 manufacturerID[3]
port 257 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 manufacturerID[4]
port 258 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 manufacturerID[5]
port 259 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 manufacturerID[6]
port 260 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 manufacturerID[7]
port 261 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 manufacturerID[8]
port 262 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 manufacturerID[9]
port 263 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 partID[0]
port 264 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 partID[10]
port 265 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 partID[11]
port 266 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 partID[12]
port 267 nsew signal output
rlabel metal3 s 0 72496 800 72616 6 partID[13]
port 268 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 partID[14]
port 269 nsew signal output
rlabel metal3 s 0 76032 800 76152 6 partID[15]
port 270 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 partID[1]
port 271 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 partID[2]
port 272 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 partID[3]
port 273 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 partID[4]
port 274 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 partID[5]
port 275 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 partID[6]
port 276 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 partID[7]
port 277 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 partID[8]
port 278 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 partID[9]
port 279 nsew signal output
rlabel metal3 s 79200 46656 80000 46776 6 probe_out[0]
port 280 nsew signal input
rlabel metal3 s 79200 49376 80000 49496 6 probe_out[10]
port 281 nsew signal input
rlabel metal3 s 79200 49648 80000 49768 6 probe_out[11]
port 282 nsew signal input
rlabel metal3 s 79200 49920 80000 50040 6 probe_out[12]
port 283 nsew signal input
rlabel metal3 s 79200 50192 80000 50312 6 probe_out[13]
port 284 nsew signal input
rlabel metal3 s 79200 50464 80000 50584 6 probe_out[14]
port 285 nsew signal input
rlabel metal3 s 79200 50736 80000 50856 6 probe_out[15]
port 286 nsew signal input
rlabel metal3 s 79200 51008 80000 51128 6 probe_out[16]
port 287 nsew signal input
rlabel metal3 s 79200 51280 80000 51400 6 probe_out[17]
port 288 nsew signal input
rlabel metal3 s 79200 51552 80000 51672 6 probe_out[18]
port 289 nsew signal input
rlabel metal3 s 79200 51824 80000 51944 6 probe_out[19]
port 290 nsew signal input
rlabel metal3 s 79200 46928 80000 47048 6 probe_out[1]
port 291 nsew signal input
rlabel metal3 s 79200 52096 80000 52216 6 probe_out[20]
port 292 nsew signal input
rlabel metal3 s 79200 52368 80000 52488 6 probe_out[21]
port 293 nsew signal input
rlabel metal3 s 79200 52640 80000 52760 6 probe_out[22]
port 294 nsew signal input
rlabel metal3 s 79200 52912 80000 53032 6 probe_out[23]
port 295 nsew signal input
rlabel metal3 s 79200 53184 80000 53304 6 probe_out[24]
port 296 nsew signal input
rlabel metal3 s 79200 53456 80000 53576 6 probe_out[25]
port 297 nsew signal input
rlabel metal3 s 79200 53728 80000 53848 6 probe_out[26]
port 298 nsew signal input
rlabel metal3 s 79200 54000 80000 54120 6 probe_out[27]
port 299 nsew signal input
rlabel metal3 s 79200 54272 80000 54392 6 probe_out[28]
port 300 nsew signal input
rlabel metal3 s 79200 54544 80000 54664 6 probe_out[29]
port 301 nsew signal input
rlabel metal3 s 79200 47200 80000 47320 6 probe_out[2]
port 302 nsew signal input
rlabel metal3 s 79200 54816 80000 54936 6 probe_out[30]
port 303 nsew signal input
rlabel metal3 s 79200 55088 80000 55208 6 probe_out[31]
port 304 nsew signal input
rlabel metal3 s 79200 55360 80000 55480 6 probe_out[32]
port 305 nsew signal input
rlabel metal3 s 79200 55632 80000 55752 6 probe_out[33]
port 306 nsew signal input
rlabel metal3 s 79200 55904 80000 56024 6 probe_out[34]
port 307 nsew signal input
rlabel metal3 s 79200 56176 80000 56296 6 probe_out[35]
port 308 nsew signal input
rlabel metal3 s 79200 56448 80000 56568 6 probe_out[36]
port 309 nsew signal input
rlabel metal3 s 79200 56720 80000 56840 6 probe_out[37]
port 310 nsew signal input
rlabel metal3 s 79200 56992 80000 57112 6 probe_out[38]
port 311 nsew signal input
rlabel metal3 s 79200 57264 80000 57384 6 probe_out[39]
port 312 nsew signal input
rlabel metal3 s 79200 47472 80000 47592 6 probe_out[3]
port 313 nsew signal input
rlabel metal3 s 79200 57536 80000 57656 6 probe_out[40]
port 314 nsew signal input
rlabel metal3 s 79200 57808 80000 57928 6 probe_out[41]
port 315 nsew signal input
rlabel metal3 s 79200 58080 80000 58200 6 probe_out[42]
port 316 nsew signal input
rlabel metal3 s 79200 58352 80000 58472 6 probe_out[43]
port 317 nsew signal input
rlabel metal3 s 79200 58624 80000 58744 6 probe_out[44]
port 318 nsew signal input
rlabel metal3 s 79200 58896 80000 59016 6 probe_out[45]
port 319 nsew signal input
rlabel metal3 s 79200 59168 80000 59288 6 probe_out[46]
port 320 nsew signal input
rlabel metal3 s 79200 59440 80000 59560 6 probe_out[47]
port 321 nsew signal input
rlabel metal3 s 79200 59712 80000 59832 6 probe_out[48]
port 322 nsew signal input
rlabel metal3 s 79200 59984 80000 60104 6 probe_out[49]
port 323 nsew signal input
rlabel metal3 s 79200 47744 80000 47864 6 probe_out[4]
port 324 nsew signal input
rlabel metal3 s 79200 60256 80000 60376 6 probe_out[50]
port 325 nsew signal input
rlabel metal3 s 79200 60528 80000 60648 6 probe_out[51]
port 326 nsew signal input
rlabel metal3 s 79200 60800 80000 60920 6 probe_out[52]
port 327 nsew signal input
rlabel metal3 s 79200 61072 80000 61192 6 probe_out[53]
port 328 nsew signal input
rlabel metal3 s 79200 61344 80000 61464 6 probe_out[54]
port 329 nsew signal input
rlabel metal3 s 79200 61616 80000 61736 6 probe_out[55]
port 330 nsew signal input
rlabel metal3 s 79200 61888 80000 62008 6 probe_out[56]
port 331 nsew signal input
rlabel metal3 s 79200 62160 80000 62280 6 probe_out[57]
port 332 nsew signal input
rlabel metal3 s 79200 62432 80000 62552 6 probe_out[58]
port 333 nsew signal input
rlabel metal3 s 79200 62704 80000 62824 6 probe_out[59]
port 334 nsew signal input
rlabel metal3 s 79200 48016 80000 48136 6 probe_out[5]
port 335 nsew signal input
rlabel metal3 s 79200 62976 80000 63096 6 probe_out[60]
port 336 nsew signal input
rlabel metal3 s 79200 63248 80000 63368 6 probe_out[61]
port 337 nsew signal input
rlabel metal3 s 79200 63520 80000 63640 6 probe_out[62]
port 338 nsew signal input
rlabel metal3 s 79200 63792 80000 63912 6 probe_out[63]
port 339 nsew signal input
rlabel metal3 s 79200 64064 80000 64184 6 probe_out[64]
port 340 nsew signal input
rlabel metal3 s 79200 64336 80000 64456 6 probe_out[65]
port 341 nsew signal input
rlabel metal3 s 79200 64608 80000 64728 6 probe_out[66]
port 342 nsew signal input
rlabel metal3 s 79200 64880 80000 65000 6 probe_out[67]
port 343 nsew signal input
rlabel metal3 s 79200 65152 80000 65272 6 probe_out[68]
port 344 nsew signal input
rlabel metal3 s 79200 65424 80000 65544 6 probe_out[69]
port 345 nsew signal input
rlabel metal3 s 79200 48288 80000 48408 6 probe_out[6]
port 346 nsew signal input
rlabel metal3 s 79200 65696 80000 65816 6 probe_out[70]
port 347 nsew signal input
rlabel metal3 s 79200 65968 80000 66088 6 probe_out[71]
port 348 nsew signal input
rlabel metal3 s 79200 66240 80000 66360 6 probe_out[72]
port 349 nsew signal input
rlabel metal3 s 79200 66512 80000 66632 6 probe_out[73]
port 350 nsew signal input
rlabel metal3 s 79200 66784 80000 66904 6 probe_out[74]
port 351 nsew signal input
rlabel metal3 s 79200 67056 80000 67176 6 probe_out[75]
port 352 nsew signal input
rlabel metal3 s 79200 67328 80000 67448 6 probe_out[76]
port 353 nsew signal input
rlabel metal3 s 79200 67600 80000 67720 6 probe_out[77]
port 354 nsew signal input
rlabel metal3 s 79200 67872 80000 67992 6 probe_out[78]
port 355 nsew signal input
rlabel metal3 s 79200 68144 80000 68264 6 probe_out[79]
port 356 nsew signal input
rlabel metal3 s 79200 48560 80000 48680 6 probe_out[7]
port 357 nsew signal input
rlabel metal3 s 79200 68416 80000 68536 6 probe_out[80]
port 358 nsew signal input
rlabel metal3 s 79200 68688 80000 68808 6 probe_out[81]
port 359 nsew signal input
rlabel metal3 s 79200 68960 80000 69080 6 probe_out[82]
port 360 nsew signal input
rlabel metal3 s 79200 69232 80000 69352 6 probe_out[83]
port 361 nsew signal input
rlabel metal3 s 79200 69504 80000 69624 6 probe_out[84]
port 362 nsew signal input
rlabel metal3 s 79200 69776 80000 69896 6 probe_out[85]
port 363 nsew signal input
rlabel metal3 s 79200 70048 80000 70168 6 probe_out[86]
port 364 nsew signal input
rlabel metal3 s 79200 70320 80000 70440 6 probe_out[87]
port 365 nsew signal input
rlabel metal3 s 79200 70592 80000 70712 6 probe_out[88]
port 366 nsew signal input
rlabel metal3 s 79200 70864 80000 70984 6 probe_out[89]
port 367 nsew signal input
rlabel metal3 s 79200 48832 80000 48952 6 probe_out[8]
port 368 nsew signal input
rlabel metal3 s 79200 71136 80000 71256 6 probe_out[90]
port 369 nsew signal input
rlabel metal3 s 79200 71408 80000 71528 6 probe_out[91]
port 370 nsew signal input
rlabel metal3 s 79200 71680 80000 71800 6 probe_out[92]
port 371 nsew signal input
rlabel metal3 s 79200 71952 80000 72072 6 probe_out[93]
port 372 nsew signal input
rlabel metal3 s 79200 72224 80000 72344 6 probe_out[94]
port 373 nsew signal input
rlabel metal3 s 79200 72496 80000 72616 6 probe_out[95]
port 374 nsew signal input
rlabel metal3 s 79200 72768 80000 72888 6 probe_out[96]
port 375 nsew signal input
rlabel metal3 s 79200 73040 80000 73160 6 probe_out[97]
port 376 nsew signal input
rlabel metal3 s 79200 49104 80000 49224 6 probe_out[9]
port 377 nsew signal input
rlabel metal4 s 4208 2128 4528 82736 6 vccd1
port 378 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 82736 6 vccd1
port 378 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 82736 6 vccd1
port 378 nsew power bidirectional
rlabel metal3 s 0 77800 800 77920 6 versionID[0]
port 379 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 versionID[1]
port 380 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 versionID[2]
port 381 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 versionID[3]
port 382 nsew signal output
rlabel metal4 s 19568 2128 19888 82736 6 vssd1
port 383 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 82736 6 vssd1
port 383 nsew ground bidirectional
rlabel metal2 s 1306 0 1362 800 6 wb_clk_i
port 384 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wb_rst_i
port 385 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 386 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[0]
port 387 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[10]
port 388 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[11]
port 389 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[12]
port 390 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[13]
port 391 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[14]
port 392 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_adr_i[15]
port 393 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_adr_i[16]
port 394 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_adr_i[17]
port 395 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wbs_adr_i[18]
port 396 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_adr_i[19]
port 397 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[1]
port 398 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[20]
port 399 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_adr_i[21]
port 400 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_adr_i[22]
port 401 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_adr_i[23]
port 402 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_adr_i[24]
port 403 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 wbs_adr_i[25]
port 404 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 wbs_adr_i[26]
port 405 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_adr_i[27]
port 406 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 wbs_adr_i[28]
port 407 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_adr_i[29]
port 408 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[2]
port 409 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 wbs_adr_i[30]
port 410 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 wbs_adr_i[31]
port 411 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[3]
port 412 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[4]
port 413 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[5]
port 414 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[6]
port 415 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[7]
port 416 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[8]
port 417 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[9]
port 418 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_cyc_i
port 419 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_data_i[0]
port 420 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_data_i[10]
port 421 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_data_i[11]
port 422 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_data_i[12]
port 423 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_data_i[13]
port 424 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_data_i[14]
port 425 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_data_i[15]
port 426 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_data_i[16]
port 427 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_data_i[17]
port 428 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_data_i[18]
port 429 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 wbs_data_i[19]
port 430 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_data_i[1]
port 431 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wbs_data_i[20]
port 432 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 wbs_data_i[21]
port 433 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_data_i[22]
port 434 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_data_i[23]
port 435 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 wbs_data_i[24]
port 436 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_data_i[25]
port 437 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_data_i[26]
port 438 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 wbs_data_i[27]
port 439 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 wbs_data_i[28]
port 440 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 wbs_data_i[29]
port 441 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_data_i[2]
port 442 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 wbs_data_i[30]
port 443 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 wbs_data_i[31]
port 444 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_data_i[3]
port 445 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_data_i[4]
port 446 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_data_i[5]
port 447 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_data_i[6]
port 448 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_data_i[7]
port 449 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_data_i[8]
port 450 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_data_i[9]
port 451 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_data_o[0]
port 452 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_data_o[10]
port 453 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_data_o[11]
port 454 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_data_o[12]
port 455 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_data_o[13]
port 456 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_data_o[14]
port 457 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_data_o[15]
port 458 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_data_o[16]
port 459 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_data_o[17]
port 460 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_data_o[18]
port 461 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_data_o[19]
port 462 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_data_o[1]
port 463 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_data_o[20]
port 464 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 wbs_data_o[21]
port 465 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_data_o[22]
port 466 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_data_o[23]
port 467 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 wbs_data_o[24]
port 468 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 wbs_data_o[25]
port 469 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 wbs_data_o[26]
port 470 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 wbs_data_o[27]
port 471 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 wbs_data_o[28]
port 472 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 wbs_data_o[29]
port 473 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_data_o[2]
port 474 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 wbs_data_o[30]
port 475 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 wbs_data_o[31]
port 476 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 wbs_data_o[3]
port 477 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_data_o[4]
port 478 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_data_o[5]
port 479 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_data_o[6]
port 480 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_data_o[7]
port 481 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_data_o[8]
port 482 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_data_o[9]
port 483 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_sel_i[0]
port 484 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[1]
port 485 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_sel_i[2]
port 486 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_sel_i[3]
port 487 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_stb_i
port 488 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_we_i
port 489 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 85000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14070718
string GDS_FILE /mnt/f/WSL/ASIC/ExperiarSoC/openlane/CaravelHost/runs/23_05_11_23_18/results/signoff/CaravelHost.magic.gds
string GDS_START 981186
<< end >>

