magic
tech sky130A
magscale 1 2
timestamp 1652998313
<< obsli1 >>
rect 1104 2159 68816 97393
<< obsm1 >>
rect 14 416 69998 97424
<< metal2 >>
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2318 0 2374 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6550 0 6606 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9310 0 9366 800
rect 10046 0 10102 800
rect 10782 0 10838 800
rect 11426 0 11482 800
rect 12162 0 12218 800
rect 12806 0 12862 800
rect 13542 0 13598 800
rect 14278 0 14334 800
rect 14922 0 14978 800
rect 15658 0 15714 800
rect 16394 0 16450 800
rect 17038 0 17094 800
rect 17774 0 17830 800
rect 18418 0 18474 800
rect 19154 0 19210 800
rect 19890 0 19946 800
rect 20534 0 20590 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22650 0 22706 800
rect 23386 0 23442 800
rect 24030 0 24086 800
rect 24766 0 24822 800
rect 25410 0 25466 800
rect 26146 0 26202 800
rect 26882 0 26938 800
rect 27526 0 27582 800
rect 28262 0 28318 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30378 0 30434 800
rect 31022 0 31078 800
rect 31758 0 31814 800
rect 32494 0 32550 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34518 0 34574 800
rect 35254 0 35310 800
rect 35990 0 36046 800
rect 36634 0 36690 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38750 0 38806 800
rect 39486 0 39542 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41510 0 41566 800
rect 42246 0 42302 800
rect 42982 0 43038 800
rect 43626 0 43682 800
rect 44362 0 44418 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46478 0 46534 800
rect 47122 0 47178 800
rect 47858 0 47914 800
rect 48594 0 48650 800
rect 49238 0 49294 800
rect 49974 0 50030 800
rect 50618 0 50674 800
rect 51354 0 51410 800
rect 52090 0 52146 800
rect 52734 0 52790 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54850 0 54906 800
rect 55586 0 55642 800
rect 56230 0 56286 800
rect 56966 0 57022 800
rect 57702 0 57758 800
rect 58346 0 58402 800
rect 59082 0 59138 800
rect 59726 0 59782 800
rect 60462 0 60518 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62578 0 62634 800
rect 63222 0 63278 800
rect 63958 0 64014 800
rect 64694 0 64750 800
rect 65338 0 65394 800
rect 66074 0 66130 800
rect 66718 0 66774 800
rect 67454 0 67510 800
rect 68190 0 68246 800
rect 68834 0 68890 800
rect 69570 0 69626 800
<< obsm2 >>
rect 20 856 69994 99521
rect 20 167 238 856
rect 406 167 882 856
rect 1050 167 1618 856
rect 1786 167 2262 856
rect 2430 167 2998 856
rect 3166 167 3734 856
rect 3902 167 4378 856
rect 4546 167 5114 856
rect 5282 167 5758 856
rect 5926 167 6494 856
rect 6662 167 7230 856
rect 7398 167 7874 856
rect 8042 167 8610 856
rect 8778 167 9254 856
rect 9422 167 9990 856
rect 10158 167 10726 856
rect 10894 167 11370 856
rect 11538 167 12106 856
rect 12274 167 12750 856
rect 12918 167 13486 856
rect 13654 167 14222 856
rect 14390 167 14866 856
rect 15034 167 15602 856
rect 15770 167 16338 856
rect 16506 167 16982 856
rect 17150 167 17718 856
rect 17886 167 18362 856
rect 18530 167 19098 856
rect 19266 167 19834 856
rect 20002 167 20478 856
rect 20646 167 21214 856
rect 21382 167 21858 856
rect 22026 167 22594 856
rect 22762 167 23330 856
rect 23498 167 23974 856
rect 24142 167 24710 856
rect 24878 167 25354 856
rect 25522 167 26090 856
rect 26258 167 26826 856
rect 26994 167 27470 856
rect 27638 167 28206 856
rect 28374 167 28942 856
rect 29110 167 29586 856
rect 29754 167 30322 856
rect 30490 167 30966 856
rect 31134 167 31702 856
rect 31870 167 32438 856
rect 32606 167 33082 856
rect 33250 167 33818 856
rect 33986 167 34462 856
rect 34630 167 35198 856
rect 35366 167 35934 856
rect 36102 167 36578 856
rect 36746 167 37314 856
rect 37482 167 37958 856
rect 38126 167 38694 856
rect 38862 167 39430 856
rect 39598 167 40074 856
rect 40242 167 40810 856
rect 40978 167 41454 856
rect 41622 167 42190 856
rect 42358 167 42926 856
rect 43094 167 43570 856
rect 43738 167 44306 856
rect 44474 167 45042 856
rect 45210 167 45686 856
rect 45854 167 46422 856
rect 46590 167 47066 856
rect 47234 167 47802 856
rect 47970 167 48538 856
rect 48706 167 49182 856
rect 49350 167 49918 856
rect 50086 167 50562 856
rect 50730 167 51298 856
rect 51466 167 52034 856
rect 52202 167 52678 856
rect 52846 167 53414 856
rect 53582 167 54058 856
rect 54226 167 54794 856
rect 54962 167 55530 856
rect 55698 167 56174 856
rect 56342 167 56910 856
rect 57078 167 57646 856
rect 57814 167 58290 856
rect 58458 167 59026 856
rect 59194 167 59670 856
rect 59838 167 60406 856
rect 60574 167 61142 856
rect 61310 167 61786 856
rect 61954 167 62522 856
rect 62690 167 63166 856
rect 63334 167 63902 856
rect 64070 167 64638 856
rect 64806 167 65282 856
rect 65450 167 66018 856
rect 66186 167 66662 856
rect 66830 167 67398 856
rect 67566 167 68134 856
rect 68302 167 68778 856
rect 68946 167 69514 856
rect 69682 167 69994 856
<< metal3 >>
rect 69200 99696 70000 99816
rect 69200 99424 70000 99544
rect 69200 99152 70000 99272
rect 69200 98880 70000 99000
rect 69200 98472 70000 98592
rect 69200 98200 70000 98320
rect 69200 97928 70000 98048
rect 69200 97656 70000 97776
rect 69200 97248 70000 97368
rect 69200 96976 70000 97096
rect 69200 96704 70000 96824
rect 69200 96432 70000 96552
rect 69200 96024 70000 96144
rect 69200 95752 70000 95872
rect 69200 95480 70000 95600
rect 69200 95208 70000 95328
rect 69200 94936 70000 95056
rect 69200 94528 70000 94648
rect 69200 94256 70000 94376
rect 69200 93984 70000 94104
rect 69200 93712 70000 93832
rect 69200 93304 70000 93424
rect 69200 93032 70000 93152
rect 69200 92760 70000 92880
rect 69200 92488 70000 92608
rect 69200 92080 70000 92200
rect 69200 91808 70000 91928
rect 69200 91536 70000 91656
rect 69200 91264 70000 91384
rect 69200 90856 70000 90976
rect 69200 90584 70000 90704
rect 69200 90312 70000 90432
rect 69200 90040 70000 90160
rect 69200 89768 70000 89888
rect 69200 89360 70000 89480
rect 69200 89088 70000 89208
rect 69200 88816 70000 88936
rect 69200 88544 70000 88664
rect 69200 88136 70000 88256
rect 69200 87864 70000 87984
rect 69200 87592 70000 87712
rect 69200 87320 70000 87440
rect 69200 86912 70000 87032
rect 69200 86640 70000 86760
rect 69200 86368 70000 86488
rect 69200 86096 70000 86216
rect 69200 85824 70000 85944
rect 69200 85416 70000 85536
rect 69200 85144 70000 85264
rect 69200 84872 70000 84992
rect 69200 84600 70000 84720
rect 69200 84192 70000 84312
rect 69200 83920 70000 84040
rect 69200 83648 70000 83768
rect 69200 83376 70000 83496
rect 69200 82968 70000 83088
rect 69200 82696 70000 82816
rect 69200 82424 70000 82544
rect 69200 82152 70000 82272
rect 69200 81744 70000 81864
rect 69200 81472 70000 81592
rect 69200 81200 70000 81320
rect 69200 80928 70000 81048
rect 69200 80656 70000 80776
rect 69200 80248 70000 80368
rect 69200 79976 70000 80096
rect 69200 79704 70000 79824
rect 69200 79432 70000 79552
rect 69200 79024 70000 79144
rect 69200 78752 70000 78872
rect 69200 78480 70000 78600
rect 69200 78208 70000 78328
rect 69200 77800 70000 77920
rect 69200 77528 70000 77648
rect 69200 77256 70000 77376
rect 69200 76984 70000 77104
rect 69200 76576 70000 76696
rect 69200 76304 70000 76424
rect 69200 76032 70000 76152
rect 69200 75760 70000 75880
rect 69200 75488 70000 75608
rect 69200 75080 70000 75200
rect 69200 74808 70000 74928
rect 69200 74536 70000 74656
rect 69200 74264 70000 74384
rect 69200 73856 70000 73976
rect 69200 73584 70000 73704
rect 69200 73312 70000 73432
rect 69200 73040 70000 73160
rect 69200 72632 70000 72752
rect 69200 72360 70000 72480
rect 69200 72088 70000 72208
rect 69200 71816 70000 71936
rect 69200 71544 70000 71664
rect 69200 71136 70000 71256
rect 69200 70864 70000 70984
rect 69200 70592 70000 70712
rect 69200 70320 70000 70440
rect 69200 69912 70000 70032
rect 69200 69640 70000 69760
rect 69200 69368 70000 69488
rect 69200 69096 70000 69216
rect 69200 68688 70000 68808
rect 69200 68416 70000 68536
rect 69200 68144 70000 68264
rect 69200 67872 70000 67992
rect 69200 67464 70000 67584
rect 69200 67192 70000 67312
rect 69200 66920 70000 67040
rect 69200 66648 70000 66768
rect 69200 66376 70000 66496
rect 69200 65968 70000 66088
rect 69200 65696 70000 65816
rect 69200 65424 70000 65544
rect 69200 65152 70000 65272
rect 69200 64744 70000 64864
rect 69200 64472 70000 64592
rect 69200 64200 70000 64320
rect 69200 63928 70000 64048
rect 69200 63520 70000 63640
rect 69200 63248 70000 63368
rect 69200 62976 70000 63096
rect 69200 62704 70000 62824
rect 69200 62296 70000 62416
rect 69200 62024 70000 62144
rect 69200 61752 70000 61872
rect 69200 61480 70000 61600
rect 69200 61208 70000 61328
rect 69200 60800 70000 60920
rect 69200 60528 70000 60648
rect 69200 60256 70000 60376
rect 69200 59984 70000 60104
rect 69200 59576 70000 59696
rect 69200 59304 70000 59424
rect 69200 59032 70000 59152
rect 69200 58760 70000 58880
rect 69200 58352 70000 58472
rect 69200 58080 70000 58200
rect 69200 57808 70000 57928
rect 69200 57536 70000 57656
rect 69200 57264 70000 57384
rect 69200 56856 70000 56976
rect 69200 56584 70000 56704
rect 69200 56312 70000 56432
rect 69200 56040 70000 56160
rect 69200 55632 70000 55752
rect 69200 55360 70000 55480
rect 69200 55088 70000 55208
rect 69200 54816 70000 54936
rect 69200 54408 70000 54528
rect 69200 54136 70000 54256
rect 69200 53864 70000 53984
rect 69200 53592 70000 53712
rect 69200 53184 70000 53304
rect 69200 52912 70000 53032
rect 69200 52640 70000 52760
rect 69200 52368 70000 52488
rect 69200 52096 70000 52216
rect 69200 51688 70000 51808
rect 69200 51416 70000 51536
rect 69200 51144 70000 51264
rect 69200 50872 70000 50992
rect 69200 50464 70000 50584
rect 69200 50192 70000 50312
rect 69200 49920 70000 50040
rect 69200 49648 70000 49768
rect 69200 49240 70000 49360
rect 69200 48968 70000 49088
rect 69200 48696 70000 48816
rect 69200 48424 70000 48544
rect 69200 48016 70000 48136
rect 69200 47744 70000 47864
rect 69200 47472 70000 47592
rect 69200 47200 70000 47320
rect 69200 46928 70000 47048
rect 69200 46520 70000 46640
rect 69200 46248 70000 46368
rect 69200 45976 70000 46096
rect 69200 45704 70000 45824
rect 69200 45296 70000 45416
rect 69200 45024 70000 45144
rect 69200 44752 70000 44872
rect 69200 44480 70000 44600
rect 69200 44072 70000 44192
rect 69200 43800 70000 43920
rect 69200 43528 70000 43648
rect 69200 43256 70000 43376
rect 69200 42984 70000 43104
rect 69200 42576 70000 42696
rect 69200 42304 70000 42424
rect 69200 42032 70000 42152
rect 69200 41760 70000 41880
rect 69200 41352 70000 41472
rect 69200 41080 70000 41200
rect 69200 40808 70000 40928
rect 69200 40536 70000 40656
rect 69200 40128 70000 40248
rect 69200 39856 70000 39976
rect 69200 39584 70000 39704
rect 69200 39312 70000 39432
rect 69200 38904 70000 39024
rect 69200 38632 70000 38752
rect 69200 38360 70000 38480
rect 69200 38088 70000 38208
rect 69200 37816 70000 37936
rect 69200 37408 70000 37528
rect 69200 37136 70000 37256
rect 69200 36864 70000 36984
rect 69200 36592 70000 36712
rect 69200 36184 70000 36304
rect 69200 35912 70000 36032
rect 69200 35640 70000 35760
rect 69200 35368 70000 35488
rect 69200 34960 70000 35080
rect 69200 34688 70000 34808
rect 69200 34416 70000 34536
rect 69200 34144 70000 34264
rect 69200 33736 70000 33856
rect 69200 33464 70000 33584
rect 69200 33192 70000 33312
rect 69200 32920 70000 33040
rect 69200 32648 70000 32768
rect 69200 32240 70000 32360
rect 69200 31968 70000 32088
rect 69200 31696 70000 31816
rect 69200 31424 70000 31544
rect 69200 31016 70000 31136
rect 69200 30744 70000 30864
rect 69200 30472 70000 30592
rect 69200 30200 70000 30320
rect 69200 29792 70000 29912
rect 69200 29520 70000 29640
rect 69200 29248 70000 29368
rect 69200 28976 70000 29096
rect 69200 28704 70000 28824
rect 69200 28296 70000 28416
rect 69200 28024 70000 28144
rect 69200 27752 70000 27872
rect 69200 27480 70000 27600
rect 69200 27072 70000 27192
rect 69200 26800 70000 26920
rect 69200 26528 70000 26648
rect 69200 26256 70000 26376
rect 69200 25848 70000 25968
rect 69200 25576 70000 25696
rect 69200 25304 70000 25424
rect 69200 25032 70000 25152
rect 69200 24624 70000 24744
rect 69200 24352 70000 24472
rect 69200 24080 70000 24200
rect 69200 23808 70000 23928
rect 69200 23536 70000 23656
rect 69200 23128 70000 23248
rect 69200 22856 70000 22976
rect 69200 22584 70000 22704
rect 69200 22312 70000 22432
rect 69200 21904 70000 22024
rect 69200 21632 70000 21752
rect 69200 21360 70000 21480
rect 69200 21088 70000 21208
rect 69200 20680 70000 20800
rect 69200 20408 70000 20528
rect 69200 20136 70000 20256
rect 69200 19864 70000 19984
rect 69200 19456 70000 19576
rect 69200 19184 70000 19304
rect 69200 18912 70000 19032
rect 69200 18640 70000 18760
rect 69200 18368 70000 18488
rect 69200 17960 70000 18080
rect 69200 17688 70000 17808
rect 69200 17416 70000 17536
rect 69200 17144 70000 17264
rect 69200 16736 70000 16856
rect 69200 16464 70000 16584
rect 69200 16192 70000 16312
rect 69200 15920 70000 16040
rect 69200 15512 70000 15632
rect 69200 15240 70000 15360
rect 69200 14968 70000 15088
rect 69200 14696 70000 14816
rect 69200 14424 70000 14544
rect 69200 14016 70000 14136
rect 69200 13744 70000 13864
rect 69200 13472 70000 13592
rect 69200 13200 70000 13320
rect 69200 12792 70000 12912
rect 69200 12520 70000 12640
rect 69200 12248 70000 12368
rect 69200 11976 70000 12096
rect 69200 11568 70000 11688
rect 69200 11296 70000 11416
rect 69200 11024 70000 11144
rect 69200 10752 70000 10872
rect 69200 10344 70000 10464
rect 69200 10072 70000 10192
rect 69200 9800 70000 9920
rect 69200 9528 70000 9648
rect 69200 9256 70000 9376
rect 69200 8848 70000 8968
rect 69200 8576 70000 8696
rect 69200 8304 70000 8424
rect 69200 8032 70000 8152
rect 69200 7624 70000 7744
rect 69200 7352 70000 7472
rect 69200 7080 70000 7200
rect 69200 6808 70000 6928
rect 69200 6400 70000 6520
rect 69200 6128 70000 6248
rect 69200 5856 70000 5976
rect 69200 5584 70000 5704
rect 69200 5176 70000 5296
rect 69200 4904 70000 5024
rect 69200 4632 70000 4752
rect 69200 4360 70000 4480
rect 69200 4088 70000 4208
rect 69200 3680 70000 3800
rect 69200 3408 70000 3528
rect 69200 3136 70000 3256
rect 69200 2864 70000 2984
rect 69200 2456 70000 2576
rect 69200 2184 70000 2304
rect 69200 1912 70000 2032
rect 69200 1640 70000 1760
rect 69200 1232 70000 1352
rect 69200 960 70000 1080
rect 69200 688 70000 808
rect 69200 416 70000 536
rect 69200 144 70000 264
<< obsm3 >>
rect 4210 98800 69120 99517
rect 4210 98672 69999 98800
rect 4210 97576 69120 98672
rect 4210 97448 69999 97576
rect 4210 96352 69120 97448
rect 4210 96224 69999 96352
rect 4210 94856 69120 96224
rect 4210 94728 69999 94856
rect 4210 93632 69120 94728
rect 4210 93504 69999 93632
rect 4210 92408 69120 93504
rect 4210 92280 69999 92408
rect 4210 91184 69120 92280
rect 4210 91056 69999 91184
rect 4210 89688 69120 91056
rect 4210 89560 69999 89688
rect 4210 88464 69120 89560
rect 4210 88336 69999 88464
rect 4210 87240 69120 88336
rect 4210 87112 69999 87240
rect 4210 85744 69120 87112
rect 4210 85616 69999 85744
rect 4210 84520 69120 85616
rect 4210 84392 69999 84520
rect 4210 83296 69120 84392
rect 4210 83168 69999 83296
rect 4210 82072 69120 83168
rect 4210 81944 69999 82072
rect 4210 80576 69120 81944
rect 4210 80448 69999 80576
rect 4210 79352 69120 80448
rect 4210 79224 69999 79352
rect 4210 78128 69120 79224
rect 4210 78000 69999 78128
rect 4210 76904 69120 78000
rect 4210 76776 69999 76904
rect 4210 75408 69120 76776
rect 4210 75280 69999 75408
rect 4210 74184 69120 75280
rect 4210 74056 69999 74184
rect 4210 72960 69120 74056
rect 4210 72832 69999 72960
rect 4210 71464 69120 72832
rect 4210 71336 69999 71464
rect 4210 70240 69120 71336
rect 4210 70112 69999 70240
rect 4210 69016 69120 70112
rect 4210 68888 69999 69016
rect 4210 67792 69120 68888
rect 4210 67664 69999 67792
rect 4210 66296 69120 67664
rect 4210 66168 69999 66296
rect 4210 65072 69120 66168
rect 4210 64944 69999 65072
rect 4210 63848 69120 64944
rect 4210 63720 69999 63848
rect 4210 62624 69120 63720
rect 4210 62496 69999 62624
rect 4210 61128 69120 62496
rect 4210 61000 69999 61128
rect 4210 59904 69120 61000
rect 4210 59776 69999 59904
rect 4210 58680 69120 59776
rect 4210 58552 69999 58680
rect 4210 57184 69120 58552
rect 4210 57056 69999 57184
rect 4210 55960 69120 57056
rect 4210 55832 69999 55960
rect 4210 54736 69120 55832
rect 4210 54608 69999 54736
rect 4210 53512 69120 54608
rect 4210 53384 69999 53512
rect 4210 52016 69120 53384
rect 4210 51888 69999 52016
rect 4210 50792 69120 51888
rect 4210 50664 69999 50792
rect 4210 49568 69120 50664
rect 4210 49440 69999 49568
rect 4210 48344 69120 49440
rect 4210 48216 69999 48344
rect 4210 46848 69120 48216
rect 4210 46720 69999 46848
rect 4210 45624 69120 46720
rect 4210 45496 69999 45624
rect 4210 44400 69120 45496
rect 4210 44272 69999 44400
rect 4210 42904 69120 44272
rect 4210 42776 69999 42904
rect 4210 41680 69120 42776
rect 4210 41552 69999 41680
rect 4210 40456 69120 41552
rect 4210 40328 69999 40456
rect 4210 39232 69120 40328
rect 4210 39104 69999 39232
rect 4210 37736 69120 39104
rect 4210 37608 69999 37736
rect 4210 36512 69120 37608
rect 4210 36384 69999 36512
rect 4210 35288 69120 36384
rect 4210 35160 69999 35288
rect 4210 34064 69120 35160
rect 4210 33936 69999 34064
rect 4210 32568 69120 33936
rect 4210 32440 69999 32568
rect 4210 31344 69120 32440
rect 4210 31216 69999 31344
rect 4210 30120 69120 31216
rect 4210 29992 69999 30120
rect 4210 28624 69120 29992
rect 4210 28496 69999 28624
rect 4210 27400 69120 28496
rect 4210 27272 69999 27400
rect 4210 26176 69120 27272
rect 4210 26048 69999 26176
rect 4210 24952 69120 26048
rect 4210 24824 69999 24952
rect 4210 23456 69120 24824
rect 4210 23328 69999 23456
rect 4210 22232 69120 23328
rect 4210 22104 69999 22232
rect 4210 21008 69120 22104
rect 4210 20880 69999 21008
rect 4210 19784 69120 20880
rect 4210 19656 69999 19784
rect 4210 18288 69120 19656
rect 4210 18160 69999 18288
rect 4210 17064 69120 18160
rect 4210 16936 69999 17064
rect 4210 15840 69120 16936
rect 4210 15712 69999 15840
rect 4210 14344 69120 15712
rect 4210 14216 69999 14344
rect 4210 13120 69120 14216
rect 4210 12992 69999 13120
rect 4210 11896 69120 12992
rect 4210 11768 69999 11896
rect 4210 10672 69120 11768
rect 4210 10544 69999 10672
rect 4210 9176 69120 10544
rect 4210 9048 69999 9176
rect 4210 7952 69120 9048
rect 4210 7824 69999 7952
rect 4210 6728 69120 7824
rect 4210 6600 69999 6728
rect 4210 5504 69120 6600
rect 4210 5376 69999 5504
rect 4210 4008 69120 5376
rect 4210 3880 69999 4008
rect 4210 2784 69120 3880
rect 4210 2656 69999 2784
rect 4210 1560 69120 2656
rect 4210 1432 69999 1560
rect 4210 171 69120 1432
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
<< obsm4 >>
rect 38331 3571 50208 94213
rect 50688 3571 65568 94213
rect 66048 3571 69677 94213
<< labels >>
rlabel metal3 s 69200 3408 70000 3528 6 sram_addr0[0]
port 1 nsew signal output
rlabel metal3 s 69200 5856 70000 5976 6 sram_addr0[1]
port 2 nsew signal output
rlabel metal3 s 69200 8304 70000 8424 6 sram_addr0[2]
port 3 nsew signal output
rlabel metal3 s 69200 10752 70000 10872 6 sram_addr0[3]
port 4 nsew signal output
rlabel metal3 s 69200 13200 70000 13320 6 sram_addr0[4]
port 5 nsew signal output
rlabel metal3 s 69200 14696 70000 14816 6 sram_addr0[5]
port 6 nsew signal output
rlabel metal3 s 69200 16192 70000 16312 6 sram_addr0[6]
port 7 nsew signal output
rlabel metal3 s 69200 17688 70000 17808 6 sram_addr0[7]
port 8 nsew signal output
rlabel metal3 s 69200 19184 70000 19304 6 sram_addr0[8]
port 9 nsew signal output
rlabel metal3 s 69200 3680 70000 3800 6 sram_addr1[0]
port 10 nsew signal output
rlabel metal3 s 69200 6128 70000 6248 6 sram_addr1[1]
port 11 nsew signal output
rlabel metal3 s 69200 8576 70000 8696 6 sram_addr1[2]
port 12 nsew signal output
rlabel metal3 s 69200 11024 70000 11144 6 sram_addr1[3]
port 13 nsew signal output
rlabel metal3 s 69200 13472 70000 13592 6 sram_addr1[4]
port 14 nsew signal output
rlabel metal3 s 69200 14968 70000 15088 6 sram_addr1[5]
port 15 nsew signal output
rlabel metal3 s 69200 16464 70000 16584 6 sram_addr1[6]
port 16 nsew signal output
rlabel metal3 s 69200 17960 70000 18080 6 sram_addr1[7]
port 17 nsew signal output
rlabel metal3 s 69200 19456 70000 19576 6 sram_addr1[8]
port 18 nsew signal output
rlabel metal3 s 69200 2456 70000 2576 6 sram_clk0
port 19 nsew signal output
rlabel metal3 s 69200 2864 70000 2984 6 sram_clk1
port 20 nsew signal output
rlabel metal3 s 69200 4088 70000 4208 6 sram_csb0[0]
port 21 nsew signal output
rlabel metal3 s 69200 6400 70000 6520 6 sram_csb0[1]
port 22 nsew signal output
rlabel metal3 s 69200 8848 70000 8968 6 sram_csb0[2]
port 23 nsew signal output
rlabel metal3 s 69200 11296 70000 11416 6 sram_csb0[3]
port 24 nsew signal output
rlabel metal3 s 69200 4360 70000 4480 6 sram_csb1[0]
port 25 nsew signal output
rlabel metal3 s 69200 6808 70000 6928 6 sram_csb1[1]
port 26 nsew signal output
rlabel metal3 s 69200 9256 70000 9376 6 sram_csb1[2]
port 27 nsew signal output
rlabel metal3 s 69200 11568 70000 11688 6 sram_csb1[3]
port 28 nsew signal output
rlabel metal3 s 69200 4632 70000 4752 6 sram_din0[0]
port 29 nsew signal output
rlabel metal3 s 69200 21632 70000 21752 6 sram_din0[10]
port 30 nsew signal output
rlabel metal3 s 69200 22584 70000 22704 6 sram_din0[11]
port 31 nsew signal output
rlabel metal3 s 69200 23536 70000 23656 6 sram_din0[12]
port 32 nsew signal output
rlabel metal3 s 69200 24352 70000 24472 6 sram_din0[13]
port 33 nsew signal output
rlabel metal3 s 69200 25304 70000 25424 6 sram_din0[14]
port 34 nsew signal output
rlabel metal3 s 69200 26256 70000 26376 6 sram_din0[15]
port 35 nsew signal output
rlabel metal3 s 69200 27072 70000 27192 6 sram_din0[16]
port 36 nsew signal output
rlabel metal3 s 69200 28024 70000 28144 6 sram_din0[17]
port 37 nsew signal output
rlabel metal3 s 69200 28976 70000 29096 6 sram_din0[18]
port 38 nsew signal output
rlabel metal3 s 69200 29792 70000 29912 6 sram_din0[19]
port 39 nsew signal output
rlabel metal3 s 69200 7080 70000 7200 6 sram_din0[1]
port 40 nsew signal output
rlabel metal3 s 69200 30744 70000 30864 6 sram_din0[20]
port 41 nsew signal output
rlabel metal3 s 69200 31696 70000 31816 6 sram_din0[21]
port 42 nsew signal output
rlabel metal3 s 69200 32648 70000 32768 6 sram_din0[22]
port 43 nsew signal output
rlabel metal3 s 69200 33464 70000 33584 6 sram_din0[23]
port 44 nsew signal output
rlabel metal3 s 69200 34416 70000 34536 6 sram_din0[24]
port 45 nsew signal output
rlabel metal3 s 69200 35368 70000 35488 6 sram_din0[25]
port 46 nsew signal output
rlabel metal3 s 69200 36184 70000 36304 6 sram_din0[26]
port 47 nsew signal output
rlabel metal3 s 69200 37136 70000 37256 6 sram_din0[27]
port 48 nsew signal output
rlabel metal3 s 69200 38088 70000 38208 6 sram_din0[28]
port 49 nsew signal output
rlabel metal3 s 69200 38904 70000 39024 6 sram_din0[29]
port 50 nsew signal output
rlabel metal3 s 69200 9528 70000 9648 6 sram_din0[2]
port 51 nsew signal output
rlabel metal3 s 69200 39856 70000 39976 6 sram_din0[30]
port 52 nsew signal output
rlabel metal3 s 69200 40808 70000 40928 6 sram_din0[31]
port 53 nsew signal output
rlabel metal3 s 69200 11976 70000 12096 6 sram_din0[3]
port 54 nsew signal output
rlabel metal3 s 69200 13744 70000 13864 6 sram_din0[4]
port 55 nsew signal output
rlabel metal3 s 69200 15240 70000 15360 6 sram_din0[5]
port 56 nsew signal output
rlabel metal3 s 69200 16736 70000 16856 6 sram_din0[6]
port 57 nsew signal output
rlabel metal3 s 69200 18368 70000 18488 6 sram_din0[7]
port 58 nsew signal output
rlabel metal3 s 69200 19864 70000 19984 6 sram_din0[8]
port 59 nsew signal output
rlabel metal3 s 69200 20680 70000 20800 6 sram_din0[9]
port 60 nsew signal output
rlabel metal3 s 69200 4904 70000 5024 6 sram_dout0[0]
port 61 nsew signal input
rlabel metal3 s 69200 82968 70000 83088 6 sram_dout0[100]
port 62 nsew signal input
rlabel metal3 s 69200 83648 70000 83768 6 sram_dout0[101]
port 63 nsew signal input
rlabel metal3 s 69200 84192 70000 84312 6 sram_dout0[102]
port 64 nsew signal input
rlabel metal3 s 69200 84872 70000 84992 6 sram_dout0[103]
port 65 nsew signal input
rlabel metal3 s 69200 85416 70000 85536 6 sram_dout0[104]
port 66 nsew signal input
rlabel metal3 s 69200 86096 70000 86216 6 sram_dout0[105]
port 67 nsew signal input
rlabel metal3 s 69200 86640 70000 86760 6 sram_dout0[106]
port 68 nsew signal input
rlabel metal3 s 69200 87320 70000 87440 6 sram_dout0[107]
port 69 nsew signal input
rlabel metal3 s 69200 87864 70000 87984 6 sram_dout0[108]
port 70 nsew signal input
rlabel metal3 s 69200 88544 70000 88664 6 sram_dout0[109]
port 71 nsew signal input
rlabel metal3 s 69200 21904 70000 22024 6 sram_dout0[10]
port 72 nsew signal input
rlabel metal3 s 69200 89088 70000 89208 6 sram_dout0[110]
port 73 nsew signal input
rlabel metal3 s 69200 89768 70000 89888 6 sram_dout0[111]
port 74 nsew signal input
rlabel metal3 s 69200 90312 70000 90432 6 sram_dout0[112]
port 75 nsew signal input
rlabel metal3 s 69200 90856 70000 90976 6 sram_dout0[113]
port 76 nsew signal input
rlabel metal3 s 69200 91536 70000 91656 6 sram_dout0[114]
port 77 nsew signal input
rlabel metal3 s 69200 92080 70000 92200 6 sram_dout0[115]
port 78 nsew signal input
rlabel metal3 s 69200 92760 70000 92880 6 sram_dout0[116]
port 79 nsew signal input
rlabel metal3 s 69200 93304 70000 93424 6 sram_dout0[117]
port 80 nsew signal input
rlabel metal3 s 69200 93984 70000 94104 6 sram_dout0[118]
port 81 nsew signal input
rlabel metal3 s 69200 94528 70000 94648 6 sram_dout0[119]
port 82 nsew signal input
rlabel metal3 s 69200 22856 70000 22976 6 sram_dout0[11]
port 83 nsew signal input
rlabel metal3 s 69200 95208 70000 95328 6 sram_dout0[120]
port 84 nsew signal input
rlabel metal3 s 69200 95752 70000 95872 6 sram_dout0[121]
port 85 nsew signal input
rlabel metal3 s 69200 96432 70000 96552 6 sram_dout0[122]
port 86 nsew signal input
rlabel metal3 s 69200 96976 70000 97096 6 sram_dout0[123]
port 87 nsew signal input
rlabel metal3 s 69200 97656 70000 97776 6 sram_dout0[124]
port 88 nsew signal input
rlabel metal3 s 69200 98200 70000 98320 6 sram_dout0[125]
port 89 nsew signal input
rlabel metal3 s 69200 98880 70000 99000 6 sram_dout0[126]
port 90 nsew signal input
rlabel metal3 s 69200 99424 70000 99544 6 sram_dout0[127]
port 91 nsew signal input
rlabel metal3 s 69200 23808 70000 23928 6 sram_dout0[12]
port 92 nsew signal input
rlabel metal3 s 69200 24624 70000 24744 6 sram_dout0[13]
port 93 nsew signal input
rlabel metal3 s 69200 25576 70000 25696 6 sram_dout0[14]
port 94 nsew signal input
rlabel metal3 s 69200 26528 70000 26648 6 sram_dout0[15]
port 95 nsew signal input
rlabel metal3 s 69200 27480 70000 27600 6 sram_dout0[16]
port 96 nsew signal input
rlabel metal3 s 69200 28296 70000 28416 6 sram_dout0[17]
port 97 nsew signal input
rlabel metal3 s 69200 29248 70000 29368 6 sram_dout0[18]
port 98 nsew signal input
rlabel metal3 s 69200 30200 70000 30320 6 sram_dout0[19]
port 99 nsew signal input
rlabel metal3 s 69200 7352 70000 7472 6 sram_dout0[1]
port 100 nsew signal input
rlabel metal3 s 69200 31016 70000 31136 6 sram_dout0[20]
port 101 nsew signal input
rlabel metal3 s 69200 31968 70000 32088 6 sram_dout0[21]
port 102 nsew signal input
rlabel metal3 s 69200 32920 70000 33040 6 sram_dout0[22]
port 103 nsew signal input
rlabel metal3 s 69200 33736 70000 33856 6 sram_dout0[23]
port 104 nsew signal input
rlabel metal3 s 69200 34688 70000 34808 6 sram_dout0[24]
port 105 nsew signal input
rlabel metal3 s 69200 35640 70000 35760 6 sram_dout0[25]
port 106 nsew signal input
rlabel metal3 s 69200 36592 70000 36712 6 sram_dout0[26]
port 107 nsew signal input
rlabel metal3 s 69200 37408 70000 37528 6 sram_dout0[27]
port 108 nsew signal input
rlabel metal3 s 69200 38360 70000 38480 6 sram_dout0[28]
port 109 nsew signal input
rlabel metal3 s 69200 39312 70000 39432 6 sram_dout0[29]
port 110 nsew signal input
rlabel metal3 s 69200 9800 70000 9920 6 sram_dout0[2]
port 111 nsew signal input
rlabel metal3 s 69200 40128 70000 40248 6 sram_dout0[30]
port 112 nsew signal input
rlabel metal3 s 69200 41080 70000 41200 6 sram_dout0[31]
port 113 nsew signal input
rlabel metal3 s 69200 41760 70000 41880 6 sram_dout0[32]
port 114 nsew signal input
rlabel metal3 s 69200 42304 70000 42424 6 sram_dout0[33]
port 115 nsew signal input
rlabel metal3 s 69200 42984 70000 43104 6 sram_dout0[34]
port 116 nsew signal input
rlabel metal3 s 69200 43528 70000 43648 6 sram_dout0[35]
port 117 nsew signal input
rlabel metal3 s 69200 44072 70000 44192 6 sram_dout0[36]
port 118 nsew signal input
rlabel metal3 s 69200 44752 70000 44872 6 sram_dout0[37]
port 119 nsew signal input
rlabel metal3 s 69200 45296 70000 45416 6 sram_dout0[38]
port 120 nsew signal input
rlabel metal3 s 69200 45976 70000 46096 6 sram_dout0[39]
port 121 nsew signal input
rlabel metal3 s 69200 12248 70000 12368 6 sram_dout0[3]
port 122 nsew signal input
rlabel metal3 s 69200 46520 70000 46640 6 sram_dout0[40]
port 123 nsew signal input
rlabel metal3 s 69200 47200 70000 47320 6 sram_dout0[41]
port 124 nsew signal input
rlabel metal3 s 69200 47744 70000 47864 6 sram_dout0[42]
port 125 nsew signal input
rlabel metal3 s 69200 48424 70000 48544 6 sram_dout0[43]
port 126 nsew signal input
rlabel metal3 s 69200 48968 70000 49088 6 sram_dout0[44]
port 127 nsew signal input
rlabel metal3 s 69200 49648 70000 49768 6 sram_dout0[45]
port 128 nsew signal input
rlabel metal3 s 69200 50192 70000 50312 6 sram_dout0[46]
port 129 nsew signal input
rlabel metal3 s 69200 50872 70000 50992 6 sram_dout0[47]
port 130 nsew signal input
rlabel metal3 s 69200 51416 70000 51536 6 sram_dout0[48]
port 131 nsew signal input
rlabel metal3 s 69200 52096 70000 52216 6 sram_dout0[49]
port 132 nsew signal input
rlabel metal3 s 69200 14016 70000 14136 6 sram_dout0[4]
port 133 nsew signal input
rlabel metal3 s 69200 52640 70000 52760 6 sram_dout0[50]
port 134 nsew signal input
rlabel metal3 s 69200 53184 70000 53304 6 sram_dout0[51]
port 135 nsew signal input
rlabel metal3 s 69200 53864 70000 53984 6 sram_dout0[52]
port 136 nsew signal input
rlabel metal3 s 69200 54408 70000 54528 6 sram_dout0[53]
port 137 nsew signal input
rlabel metal3 s 69200 55088 70000 55208 6 sram_dout0[54]
port 138 nsew signal input
rlabel metal3 s 69200 55632 70000 55752 6 sram_dout0[55]
port 139 nsew signal input
rlabel metal3 s 69200 56312 70000 56432 6 sram_dout0[56]
port 140 nsew signal input
rlabel metal3 s 69200 56856 70000 56976 6 sram_dout0[57]
port 141 nsew signal input
rlabel metal3 s 69200 57536 70000 57656 6 sram_dout0[58]
port 142 nsew signal input
rlabel metal3 s 69200 58080 70000 58200 6 sram_dout0[59]
port 143 nsew signal input
rlabel metal3 s 69200 15512 70000 15632 6 sram_dout0[5]
port 144 nsew signal input
rlabel metal3 s 69200 58760 70000 58880 6 sram_dout0[60]
port 145 nsew signal input
rlabel metal3 s 69200 59304 70000 59424 6 sram_dout0[61]
port 146 nsew signal input
rlabel metal3 s 69200 59984 70000 60104 6 sram_dout0[62]
port 147 nsew signal input
rlabel metal3 s 69200 60528 70000 60648 6 sram_dout0[63]
port 148 nsew signal input
rlabel metal3 s 69200 61208 70000 61328 6 sram_dout0[64]
port 149 nsew signal input
rlabel metal3 s 69200 61752 70000 61872 6 sram_dout0[65]
port 150 nsew signal input
rlabel metal3 s 69200 62296 70000 62416 6 sram_dout0[66]
port 151 nsew signal input
rlabel metal3 s 69200 62976 70000 63096 6 sram_dout0[67]
port 152 nsew signal input
rlabel metal3 s 69200 63520 70000 63640 6 sram_dout0[68]
port 153 nsew signal input
rlabel metal3 s 69200 64200 70000 64320 6 sram_dout0[69]
port 154 nsew signal input
rlabel metal3 s 69200 17144 70000 17264 6 sram_dout0[6]
port 155 nsew signal input
rlabel metal3 s 69200 64744 70000 64864 6 sram_dout0[70]
port 156 nsew signal input
rlabel metal3 s 69200 65424 70000 65544 6 sram_dout0[71]
port 157 nsew signal input
rlabel metal3 s 69200 65968 70000 66088 6 sram_dout0[72]
port 158 nsew signal input
rlabel metal3 s 69200 66648 70000 66768 6 sram_dout0[73]
port 159 nsew signal input
rlabel metal3 s 69200 67192 70000 67312 6 sram_dout0[74]
port 160 nsew signal input
rlabel metal3 s 69200 67872 70000 67992 6 sram_dout0[75]
port 161 nsew signal input
rlabel metal3 s 69200 68416 70000 68536 6 sram_dout0[76]
port 162 nsew signal input
rlabel metal3 s 69200 69096 70000 69216 6 sram_dout0[77]
port 163 nsew signal input
rlabel metal3 s 69200 69640 70000 69760 6 sram_dout0[78]
port 164 nsew signal input
rlabel metal3 s 69200 70320 70000 70440 6 sram_dout0[79]
port 165 nsew signal input
rlabel metal3 s 69200 18640 70000 18760 6 sram_dout0[7]
port 166 nsew signal input
rlabel metal3 s 69200 70864 70000 70984 6 sram_dout0[80]
port 167 nsew signal input
rlabel metal3 s 69200 71544 70000 71664 6 sram_dout0[81]
port 168 nsew signal input
rlabel metal3 s 69200 72088 70000 72208 6 sram_dout0[82]
port 169 nsew signal input
rlabel metal3 s 69200 72632 70000 72752 6 sram_dout0[83]
port 170 nsew signal input
rlabel metal3 s 69200 73312 70000 73432 6 sram_dout0[84]
port 171 nsew signal input
rlabel metal3 s 69200 73856 70000 73976 6 sram_dout0[85]
port 172 nsew signal input
rlabel metal3 s 69200 74536 70000 74656 6 sram_dout0[86]
port 173 nsew signal input
rlabel metal3 s 69200 75080 70000 75200 6 sram_dout0[87]
port 174 nsew signal input
rlabel metal3 s 69200 75760 70000 75880 6 sram_dout0[88]
port 175 nsew signal input
rlabel metal3 s 69200 76304 70000 76424 6 sram_dout0[89]
port 176 nsew signal input
rlabel metal3 s 69200 20136 70000 20256 6 sram_dout0[8]
port 177 nsew signal input
rlabel metal3 s 69200 76984 70000 77104 6 sram_dout0[90]
port 178 nsew signal input
rlabel metal3 s 69200 77528 70000 77648 6 sram_dout0[91]
port 179 nsew signal input
rlabel metal3 s 69200 78208 70000 78328 6 sram_dout0[92]
port 180 nsew signal input
rlabel metal3 s 69200 78752 70000 78872 6 sram_dout0[93]
port 181 nsew signal input
rlabel metal3 s 69200 79432 70000 79552 6 sram_dout0[94]
port 182 nsew signal input
rlabel metal3 s 69200 79976 70000 80096 6 sram_dout0[95]
port 183 nsew signal input
rlabel metal3 s 69200 80656 70000 80776 6 sram_dout0[96]
port 184 nsew signal input
rlabel metal3 s 69200 81200 70000 81320 6 sram_dout0[97]
port 185 nsew signal input
rlabel metal3 s 69200 81744 70000 81864 6 sram_dout0[98]
port 186 nsew signal input
rlabel metal3 s 69200 82424 70000 82544 6 sram_dout0[99]
port 187 nsew signal input
rlabel metal3 s 69200 21088 70000 21208 6 sram_dout0[9]
port 188 nsew signal input
rlabel metal3 s 69200 5176 70000 5296 6 sram_dout1[0]
port 189 nsew signal input
rlabel metal3 s 69200 83376 70000 83496 6 sram_dout1[100]
port 190 nsew signal input
rlabel metal3 s 69200 83920 70000 84040 6 sram_dout1[101]
port 191 nsew signal input
rlabel metal3 s 69200 84600 70000 84720 6 sram_dout1[102]
port 192 nsew signal input
rlabel metal3 s 69200 85144 70000 85264 6 sram_dout1[103]
port 193 nsew signal input
rlabel metal3 s 69200 85824 70000 85944 6 sram_dout1[104]
port 194 nsew signal input
rlabel metal3 s 69200 86368 70000 86488 6 sram_dout1[105]
port 195 nsew signal input
rlabel metal3 s 69200 86912 70000 87032 6 sram_dout1[106]
port 196 nsew signal input
rlabel metal3 s 69200 87592 70000 87712 6 sram_dout1[107]
port 197 nsew signal input
rlabel metal3 s 69200 88136 70000 88256 6 sram_dout1[108]
port 198 nsew signal input
rlabel metal3 s 69200 88816 70000 88936 6 sram_dout1[109]
port 199 nsew signal input
rlabel metal3 s 69200 22312 70000 22432 6 sram_dout1[10]
port 200 nsew signal input
rlabel metal3 s 69200 89360 70000 89480 6 sram_dout1[110]
port 201 nsew signal input
rlabel metal3 s 69200 90040 70000 90160 6 sram_dout1[111]
port 202 nsew signal input
rlabel metal3 s 69200 90584 70000 90704 6 sram_dout1[112]
port 203 nsew signal input
rlabel metal3 s 69200 91264 70000 91384 6 sram_dout1[113]
port 204 nsew signal input
rlabel metal3 s 69200 91808 70000 91928 6 sram_dout1[114]
port 205 nsew signal input
rlabel metal3 s 69200 92488 70000 92608 6 sram_dout1[115]
port 206 nsew signal input
rlabel metal3 s 69200 93032 70000 93152 6 sram_dout1[116]
port 207 nsew signal input
rlabel metal3 s 69200 93712 70000 93832 6 sram_dout1[117]
port 208 nsew signal input
rlabel metal3 s 69200 94256 70000 94376 6 sram_dout1[118]
port 209 nsew signal input
rlabel metal3 s 69200 94936 70000 95056 6 sram_dout1[119]
port 210 nsew signal input
rlabel metal3 s 69200 23128 70000 23248 6 sram_dout1[11]
port 211 nsew signal input
rlabel metal3 s 69200 95480 70000 95600 6 sram_dout1[120]
port 212 nsew signal input
rlabel metal3 s 69200 96024 70000 96144 6 sram_dout1[121]
port 213 nsew signal input
rlabel metal3 s 69200 96704 70000 96824 6 sram_dout1[122]
port 214 nsew signal input
rlabel metal3 s 69200 97248 70000 97368 6 sram_dout1[123]
port 215 nsew signal input
rlabel metal3 s 69200 97928 70000 98048 6 sram_dout1[124]
port 216 nsew signal input
rlabel metal3 s 69200 98472 70000 98592 6 sram_dout1[125]
port 217 nsew signal input
rlabel metal3 s 69200 99152 70000 99272 6 sram_dout1[126]
port 218 nsew signal input
rlabel metal3 s 69200 99696 70000 99816 6 sram_dout1[127]
port 219 nsew signal input
rlabel metal3 s 69200 24080 70000 24200 6 sram_dout1[12]
port 220 nsew signal input
rlabel metal3 s 69200 25032 70000 25152 6 sram_dout1[13]
port 221 nsew signal input
rlabel metal3 s 69200 25848 70000 25968 6 sram_dout1[14]
port 222 nsew signal input
rlabel metal3 s 69200 26800 70000 26920 6 sram_dout1[15]
port 223 nsew signal input
rlabel metal3 s 69200 27752 70000 27872 6 sram_dout1[16]
port 224 nsew signal input
rlabel metal3 s 69200 28704 70000 28824 6 sram_dout1[17]
port 225 nsew signal input
rlabel metal3 s 69200 29520 70000 29640 6 sram_dout1[18]
port 226 nsew signal input
rlabel metal3 s 69200 30472 70000 30592 6 sram_dout1[19]
port 227 nsew signal input
rlabel metal3 s 69200 7624 70000 7744 6 sram_dout1[1]
port 228 nsew signal input
rlabel metal3 s 69200 31424 70000 31544 6 sram_dout1[20]
port 229 nsew signal input
rlabel metal3 s 69200 32240 70000 32360 6 sram_dout1[21]
port 230 nsew signal input
rlabel metal3 s 69200 33192 70000 33312 6 sram_dout1[22]
port 231 nsew signal input
rlabel metal3 s 69200 34144 70000 34264 6 sram_dout1[23]
port 232 nsew signal input
rlabel metal3 s 69200 34960 70000 35080 6 sram_dout1[24]
port 233 nsew signal input
rlabel metal3 s 69200 35912 70000 36032 6 sram_dout1[25]
port 234 nsew signal input
rlabel metal3 s 69200 36864 70000 36984 6 sram_dout1[26]
port 235 nsew signal input
rlabel metal3 s 69200 37816 70000 37936 6 sram_dout1[27]
port 236 nsew signal input
rlabel metal3 s 69200 38632 70000 38752 6 sram_dout1[28]
port 237 nsew signal input
rlabel metal3 s 69200 39584 70000 39704 6 sram_dout1[29]
port 238 nsew signal input
rlabel metal3 s 69200 10072 70000 10192 6 sram_dout1[2]
port 239 nsew signal input
rlabel metal3 s 69200 40536 70000 40656 6 sram_dout1[30]
port 240 nsew signal input
rlabel metal3 s 69200 41352 70000 41472 6 sram_dout1[31]
port 241 nsew signal input
rlabel metal3 s 69200 42032 70000 42152 6 sram_dout1[32]
port 242 nsew signal input
rlabel metal3 s 69200 42576 70000 42696 6 sram_dout1[33]
port 243 nsew signal input
rlabel metal3 s 69200 43256 70000 43376 6 sram_dout1[34]
port 244 nsew signal input
rlabel metal3 s 69200 43800 70000 43920 6 sram_dout1[35]
port 245 nsew signal input
rlabel metal3 s 69200 44480 70000 44600 6 sram_dout1[36]
port 246 nsew signal input
rlabel metal3 s 69200 45024 70000 45144 6 sram_dout1[37]
port 247 nsew signal input
rlabel metal3 s 69200 45704 70000 45824 6 sram_dout1[38]
port 248 nsew signal input
rlabel metal3 s 69200 46248 70000 46368 6 sram_dout1[39]
port 249 nsew signal input
rlabel metal3 s 69200 12520 70000 12640 6 sram_dout1[3]
port 250 nsew signal input
rlabel metal3 s 69200 46928 70000 47048 6 sram_dout1[40]
port 251 nsew signal input
rlabel metal3 s 69200 47472 70000 47592 6 sram_dout1[41]
port 252 nsew signal input
rlabel metal3 s 69200 48016 70000 48136 6 sram_dout1[42]
port 253 nsew signal input
rlabel metal3 s 69200 48696 70000 48816 6 sram_dout1[43]
port 254 nsew signal input
rlabel metal3 s 69200 49240 70000 49360 6 sram_dout1[44]
port 255 nsew signal input
rlabel metal3 s 69200 49920 70000 50040 6 sram_dout1[45]
port 256 nsew signal input
rlabel metal3 s 69200 50464 70000 50584 6 sram_dout1[46]
port 257 nsew signal input
rlabel metal3 s 69200 51144 70000 51264 6 sram_dout1[47]
port 258 nsew signal input
rlabel metal3 s 69200 51688 70000 51808 6 sram_dout1[48]
port 259 nsew signal input
rlabel metal3 s 69200 52368 70000 52488 6 sram_dout1[49]
port 260 nsew signal input
rlabel metal3 s 69200 14424 70000 14544 6 sram_dout1[4]
port 261 nsew signal input
rlabel metal3 s 69200 52912 70000 53032 6 sram_dout1[50]
port 262 nsew signal input
rlabel metal3 s 69200 53592 70000 53712 6 sram_dout1[51]
port 263 nsew signal input
rlabel metal3 s 69200 54136 70000 54256 6 sram_dout1[52]
port 264 nsew signal input
rlabel metal3 s 69200 54816 70000 54936 6 sram_dout1[53]
port 265 nsew signal input
rlabel metal3 s 69200 55360 70000 55480 6 sram_dout1[54]
port 266 nsew signal input
rlabel metal3 s 69200 56040 70000 56160 6 sram_dout1[55]
port 267 nsew signal input
rlabel metal3 s 69200 56584 70000 56704 6 sram_dout1[56]
port 268 nsew signal input
rlabel metal3 s 69200 57264 70000 57384 6 sram_dout1[57]
port 269 nsew signal input
rlabel metal3 s 69200 57808 70000 57928 6 sram_dout1[58]
port 270 nsew signal input
rlabel metal3 s 69200 58352 70000 58472 6 sram_dout1[59]
port 271 nsew signal input
rlabel metal3 s 69200 15920 70000 16040 6 sram_dout1[5]
port 272 nsew signal input
rlabel metal3 s 69200 59032 70000 59152 6 sram_dout1[60]
port 273 nsew signal input
rlabel metal3 s 69200 59576 70000 59696 6 sram_dout1[61]
port 274 nsew signal input
rlabel metal3 s 69200 60256 70000 60376 6 sram_dout1[62]
port 275 nsew signal input
rlabel metal3 s 69200 60800 70000 60920 6 sram_dout1[63]
port 276 nsew signal input
rlabel metal3 s 69200 61480 70000 61600 6 sram_dout1[64]
port 277 nsew signal input
rlabel metal3 s 69200 62024 70000 62144 6 sram_dout1[65]
port 278 nsew signal input
rlabel metal3 s 69200 62704 70000 62824 6 sram_dout1[66]
port 279 nsew signal input
rlabel metal3 s 69200 63248 70000 63368 6 sram_dout1[67]
port 280 nsew signal input
rlabel metal3 s 69200 63928 70000 64048 6 sram_dout1[68]
port 281 nsew signal input
rlabel metal3 s 69200 64472 70000 64592 6 sram_dout1[69]
port 282 nsew signal input
rlabel metal3 s 69200 17416 70000 17536 6 sram_dout1[6]
port 283 nsew signal input
rlabel metal3 s 69200 65152 70000 65272 6 sram_dout1[70]
port 284 nsew signal input
rlabel metal3 s 69200 65696 70000 65816 6 sram_dout1[71]
port 285 nsew signal input
rlabel metal3 s 69200 66376 70000 66496 6 sram_dout1[72]
port 286 nsew signal input
rlabel metal3 s 69200 66920 70000 67040 6 sram_dout1[73]
port 287 nsew signal input
rlabel metal3 s 69200 67464 70000 67584 6 sram_dout1[74]
port 288 nsew signal input
rlabel metal3 s 69200 68144 70000 68264 6 sram_dout1[75]
port 289 nsew signal input
rlabel metal3 s 69200 68688 70000 68808 6 sram_dout1[76]
port 290 nsew signal input
rlabel metal3 s 69200 69368 70000 69488 6 sram_dout1[77]
port 291 nsew signal input
rlabel metal3 s 69200 69912 70000 70032 6 sram_dout1[78]
port 292 nsew signal input
rlabel metal3 s 69200 70592 70000 70712 6 sram_dout1[79]
port 293 nsew signal input
rlabel metal3 s 69200 18912 70000 19032 6 sram_dout1[7]
port 294 nsew signal input
rlabel metal3 s 69200 71136 70000 71256 6 sram_dout1[80]
port 295 nsew signal input
rlabel metal3 s 69200 71816 70000 71936 6 sram_dout1[81]
port 296 nsew signal input
rlabel metal3 s 69200 72360 70000 72480 6 sram_dout1[82]
port 297 nsew signal input
rlabel metal3 s 69200 73040 70000 73160 6 sram_dout1[83]
port 298 nsew signal input
rlabel metal3 s 69200 73584 70000 73704 6 sram_dout1[84]
port 299 nsew signal input
rlabel metal3 s 69200 74264 70000 74384 6 sram_dout1[85]
port 300 nsew signal input
rlabel metal3 s 69200 74808 70000 74928 6 sram_dout1[86]
port 301 nsew signal input
rlabel metal3 s 69200 75488 70000 75608 6 sram_dout1[87]
port 302 nsew signal input
rlabel metal3 s 69200 76032 70000 76152 6 sram_dout1[88]
port 303 nsew signal input
rlabel metal3 s 69200 76576 70000 76696 6 sram_dout1[89]
port 304 nsew signal input
rlabel metal3 s 69200 20408 70000 20528 6 sram_dout1[8]
port 305 nsew signal input
rlabel metal3 s 69200 77256 70000 77376 6 sram_dout1[90]
port 306 nsew signal input
rlabel metal3 s 69200 77800 70000 77920 6 sram_dout1[91]
port 307 nsew signal input
rlabel metal3 s 69200 78480 70000 78600 6 sram_dout1[92]
port 308 nsew signal input
rlabel metal3 s 69200 79024 70000 79144 6 sram_dout1[93]
port 309 nsew signal input
rlabel metal3 s 69200 79704 70000 79824 6 sram_dout1[94]
port 310 nsew signal input
rlabel metal3 s 69200 80248 70000 80368 6 sram_dout1[95]
port 311 nsew signal input
rlabel metal3 s 69200 80928 70000 81048 6 sram_dout1[96]
port 312 nsew signal input
rlabel metal3 s 69200 81472 70000 81592 6 sram_dout1[97]
port 313 nsew signal input
rlabel metal3 s 69200 82152 70000 82272 6 sram_dout1[98]
port 314 nsew signal input
rlabel metal3 s 69200 82696 70000 82816 6 sram_dout1[99]
port 315 nsew signal input
rlabel metal3 s 69200 21360 70000 21480 6 sram_dout1[9]
port 316 nsew signal input
rlabel metal3 s 69200 3136 70000 3256 6 sram_web0
port 317 nsew signal output
rlabel metal3 s 69200 5584 70000 5704 6 sram_wmask0[0]
port 318 nsew signal output
rlabel metal3 s 69200 8032 70000 8152 6 sram_wmask0[1]
port 319 nsew signal output
rlabel metal3 s 69200 10344 70000 10464 6 sram_wmask0[2]
port 320 nsew signal output
rlabel metal3 s 69200 12792 70000 12912 6 sram_wmask0[3]
port 321 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal3 s 69200 688 70000 808 6 vga_b[0]
port 323 nsew signal output
rlabel metal3 s 69200 1640 70000 1760 6 vga_b[1]
port 324 nsew signal output
rlabel metal3 s 69200 960 70000 1080 6 vga_g[0]
port 325 nsew signal output
rlabel metal3 s 69200 1912 70000 2032 6 vga_g[1]
port 326 nsew signal output
rlabel metal3 s 69200 144 70000 264 6 vga_hsync
port 327 nsew signal output
rlabel metal3 s 69200 1232 70000 1352 6 vga_r[0]
port 328 nsew signal output
rlabel metal3 s 69200 2184 70000 2304 6 vga_r[1]
port 329 nsew signal output
rlabel metal3 s 69200 416 70000 536 6 vga_vsync
port 330 nsew signal output
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal2 s 294 0 350 800 6 wb_ack_o
port 332 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wb_adr_i[0]
port 333 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wb_adr_i[10]
port 334 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wb_adr_i[11]
port 335 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wb_adr_i[12]
port 336 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wb_adr_i[13]
port 337 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wb_adr_i[14]
port 338 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wb_adr_i[15]
port 339 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wb_adr_i[16]
port 340 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wb_adr_i[17]
port 341 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wb_adr_i[18]
port 342 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wb_adr_i[19]
port 343 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wb_adr_i[1]
port 344 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wb_adr_i[20]
port 345 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wb_adr_i[21]
port 346 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wb_adr_i[22]
port 347 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wb_adr_i[23]
port 348 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wb_adr_i[2]
port 349 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wb_adr_i[3]
port 350 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb_adr_i[4]
port 351 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wb_adr_i[5]
port 352 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wb_adr_i[6]
port 353 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wb_adr_i[7]
port 354 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wb_adr_i[8]
port 355 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wb_adr_i[9]
port 356 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_clk_i
port 357 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_cyc_i
port 358 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wb_data_i[0]
port 359 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wb_data_i[10]
port 360 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wb_data_i[11]
port 361 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wb_data_i[12]
port 362 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wb_data_i[13]
port 363 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wb_data_i[14]
port 364 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wb_data_i[15]
port 365 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wb_data_i[16]
port 366 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wb_data_i[17]
port 367 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wb_data_i[18]
port 368 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wb_data_i[19]
port 369 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wb_data_i[1]
port 370 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 wb_data_i[20]
port 371 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wb_data_i[21]
port 372 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 wb_data_i[22]
port 373 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wb_data_i[23]
port 374 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wb_data_i[24]
port 375 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wb_data_i[25]
port 376 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wb_data_i[26]
port 377 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wb_data_i[27]
port 378 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wb_data_i[28]
port 379 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 wb_data_i[29]
port 380 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wb_data_i[2]
port 381 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wb_data_i[30]
port 382 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 wb_data_i[31]
port 383 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wb_data_i[3]
port 384 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wb_data_i[4]
port 385 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wb_data_i[5]
port 386 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wb_data_i[6]
port 387 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wb_data_i[7]
port 388 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wb_data_i[8]
port 389 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wb_data_i[9]
port 390 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_data_o[0]
port 391 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 wb_data_o[10]
port 392 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wb_data_o[11]
port 393 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wb_data_o[12]
port 394 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wb_data_o[13]
port 395 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 wb_data_o[14]
port 396 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wb_data_o[15]
port 397 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wb_data_o[16]
port 398 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 wb_data_o[17]
port 399 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 wb_data_o[18]
port 400 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 wb_data_o[19]
port 401 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wb_data_o[1]
port 402 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wb_data_o[20]
port 403 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 wb_data_o[21]
port 404 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wb_data_o[22]
port 405 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wb_data_o[23]
port 406 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wb_data_o[24]
port 407 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wb_data_o[25]
port 408 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 wb_data_o[26]
port 409 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 wb_data_o[27]
port 410 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 wb_data_o[28]
port 411 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 wb_data_o[29]
port 412 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wb_data_o[2]
port 413 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 wb_data_o[30]
port 414 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 wb_data_o[31]
port 415 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wb_data_o[3]
port 416 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wb_data_o[4]
port 417 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wb_data_o[5]
port 418 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wb_data_o[6]
port 419 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 wb_data_o[7]
port 420 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wb_data_o[8]
port 421 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wb_data_o[9]
port 422 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 wb_error_o
port 423 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 wb_rst_i
port 424 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wb_sel_i[0]
port 425 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wb_sel_i[1]
port 426 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wb_sel_i[2]
port 427 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wb_sel_i[3]
port 428 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wb_stall_o
port 429 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wb_stb_i
port 430 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wb_we_i
port 431 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6970546
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Video/runs/Video/results/signoff/Video.magic.gds
string GDS_START 674100
<< end >>

