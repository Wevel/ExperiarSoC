VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 500.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 496.000 35.790 500.000 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 496.000 39.930 500.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 496.000 44.530 500.000 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 496.000 48.670 500.000 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 496.000 52.810 500.000 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 496.000 56.950 500.000 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 496.000 61.090 500.000 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 496.000 65.690 500.000 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 496.000 69.830 500.000 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 496.000 493.030 500.000 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 496.000 497.170 500.000 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 496.000 501.310 500.000 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 496.000 505.450 500.000 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 496.000 510.050 500.000 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 496.000 514.190 500.000 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 496.000 518.330 500.000 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 496.000 522.470 500.000 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 496.000 526.610 500.000 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 496.000 2.210 500.000 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 496.000 480.150 500.000 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 5.480 800.000 6.080 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 20.440 800.000 21.040 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 104.080 800.000 104.680 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 111.560 800.000 112.160 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 119.040 800.000 119.640 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 126.520 800.000 127.120 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 134.000 800.000 134.600 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 141.480 800.000 142.080 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 148.960 800.000 149.560 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 156.440 800.000 157.040 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 163.920 800.000 164.520 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 171.400 800.000 172.000 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 29.960 800.000 30.560 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 178.200 800.000 178.800 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 185.680 800.000 186.280 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 193.160 800.000 193.760 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 200.640 800.000 201.240 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 208.120 800.000 208.720 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 215.600 800.000 216.200 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 223.080 800.000 223.680 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 230.560 800.000 231.160 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 40.160 800.000 40.760 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 49.680 800.000 50.280 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 59.880 800.000 60.480 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 67.360 800.000 67.960 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 74.840 800.000 75.440 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 82.320 800.000 82.920 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 89.120 800.000 89.720 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 96.600 800.000 97.200 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 7.520 800.000 8.120 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 22.480 800.000 23.080 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 106.800 800.000 107.400 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 114.280 800.000 114.880 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 121.760 800.000 122.360 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 129.240 800.000 129.840 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 136.720 800.000 137.320 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 144.200 800.000 144.800 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 151.000 800.000 151.600 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 158.480 800.000 159.080 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 165.960 800.000 166.560 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 173.440 800.000 174.040 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 32.680 800.000 33.280 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 180.920 800.000 181.520 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 188.400 800.000 189.000 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 195.880 800.000 196.480 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 203.360 800.000 203.960 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 218.320 800.000 218.920 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 225.800 800.000 226.400 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 233.280 800.000 233.880 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 238.040 800.000 238.640 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 242.800 800.000 243.400 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 42.200 800.000 42.800 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 247.560 800.000 248.160 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 253.000 800.000 253.600 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 52.400 800.000 53.000 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 61.920 800.000 62.520 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 69.400 800.000 70.000 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 76.880 800.000 77.480 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 84.360 800.000 84.960 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 91.840 800.000 92.440 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 99.320 800.000 99.920 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 25.200 800.000 25.800 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 109.520 800.000 110.120 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 117.000 800.000 117.600 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 123.800 800.000 124.400 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 131.280 800.000 131.880 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 138.760 800.000 139.360 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 146.240 800.000 146.840 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 153.720 800.000 154.320 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 161.200 800.000 161.800 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 168.680 800.000 169.280 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.160 800.000 176.760 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 34.720 800.000 35.320 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 183.640 800.000 184.240 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 191.120 800.000 191.720 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 198.600 800.000 199.200 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 206.080 800.000 206.680 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 212.880 800.000 213.480 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 220.360 800.000 220.960 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 227.840 800.000 228.440 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 235.320 800.000 235.920 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 240.080 800.000 240.680 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 245.520 800.000 246.120 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 44.920 800.000 45.520 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 250.280 800.000 250.880 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 255.040 800.000 255.640 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 55.120 800.000 55.720 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 64.640 800.000 65.240 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 72.120 800.000 72.720 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 79.600 800.000 80.200 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 87.080 800.000 87.680 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 94.560 800.000 95.160 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 102.040 800.000 102.640 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 10.240 800.000 10.840 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 27.920 800.000 28.520 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 37.440 800.000 38.040 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 47.640 800.000 48.240 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 57.160 800.000 57.760 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 12.960 800.000 13.560 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 15.000 800.000 15.600 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 17.720 800.000 18.320 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 496.000 6.350 500.000 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 496.000 10.490 500.000 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 496.000 484.290 500.000 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 496.000 488.890 500.000 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 496.000 73.970 500.000 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 496.000 116.290 500.000 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 496.000 120.430 500.000 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 496.000 124.570 500.000 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 496.000 129.170 500.000 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 496.000 133.310 500.000 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 496.000 137.450 500.000 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 496.000 141.590 500.000 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 496.000 145.730 500.000 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 496.000 150.330 500.000 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 496.000 154.470 500.000 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 496.000 78.110 500.000 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 496.000 158.610 500.000 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 496.000 162.750 500.000 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 496.000 166.890 500.000 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 496.000 171.490 500.000 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 496.000 175.630 500.000 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 496.000 179.770 500.000 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 496.000 183.910 500.000 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 496.000 188.050 500.000 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 496.000 192.650 500.000 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 496.000 82.250 500.000 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 496.000 200.930 500.000 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 496.000 205.070 500.000 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 496.000 86.850 500.000 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 496.000 90.990 500.000 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 496.000 95.130 500.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 496.000 99.270 500.000 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 496.000 103.410 500.000 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 496.000 108.010 500.000 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 496.000 112.150 500.000 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 496.000 209.210 500.000 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 496.000 251.530 500.000 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 496.000 256.130 500.000 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 496.000 260.270 500.000 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 496.000 264.410 500.000 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 496.000 268.550 500.000 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 496.000 272.690 500.000 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 496.000 277.290 500.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 496.000 281.430 500.000 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 496.000 285.570 500.000 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 496.000 289.710 500.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 496.000 213.810 500.000 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 496.000 293.850 500.000 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 496.000 298.450 500.000 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 496.000 302.590 500.000 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 496.000 306.730 500.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 496.000 310.870 500.000 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 496.000 315.010 500.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 496.000 319.610 500.000 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 496.000 323.750 500.000 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 496.000 327.890 500.000 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 496.000 332.030 500.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 496.000 217.950 500.000 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 496.000 336.170 500.000 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 496.000 340.770 500.000 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 496.000 344.910 500.000 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 496.000 349.050 500.000 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 496.000 353.190 500.000 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 496.000 357.330 500.000 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 496.000 361.930 500.000 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 496.000 366.070 500.000 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 496.000 370.210 500.000 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 496.000 374.350 500.000 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 496.000 222.090 500.000 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 496.000 378.490 500.000 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 496.000 383.090 500.000 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 496.000 387.230 500.000 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 496.000 391.370 500.000 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 496.000 395.510 500.000 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 496.000 399.650 500.000 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 496.000 404.250 500.000 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 496.000 408.390 500.000 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 496.000 412.530 500.000 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 496.000 416.670 500.000 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 496.000 226.230 500.000 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 496.000 420.810 500.000 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 496.000 425.410 500.000 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 496.000 429.550 500.000 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 496.000 433.690 500.000 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 496.000 437.830 500.000 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 496.000 441.970 500.000 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 496.000 446.570 500.000 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 496.000 450.710 500.000 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 496.000 454.850 500.000 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 496.000 458.990 500.000 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 496.000 230.370 500.000 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 496.000 463.130 500.000 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 496.000 467.730 500.000 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 496.000 471.870 500.000 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 496.000 476.010 500.000 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 496.000 234.970 500.000 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 496.000 239.110 500.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 496.000 243.250 500.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 496.000 247.390 500.000 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 496.000 531.210 500.000 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 496.000 573.530 500.000 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 496.000 577.670 500.000 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 496.000 581.810 500.000 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 496.000 585.950 500.000 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 496.000 590.090 500.000 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 496.000 594.690 500.000 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 496.000 598.830 500.000 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 496.000 602.970 500.000 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 496.000 607.110 500.000 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 496.000 611.250 500.000 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 496.000 535.350 500.000 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 496.000 615.850 500.000 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 496.000 619.990 500.000 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 496.000 624.130 500.000 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 496.000 628.270 500.000 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 496.000 632.410 500.000 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 496.000 637.010 500.000 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 496.000 641.150 500.000 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 496.000 645.290 500.000 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 496.000 649.430 500.000 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 496.000 653.570 500.000 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 496.000 539.490 500.000 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 496.000 658.170 500.000 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 496.000 662.310 500.000 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 496.000 666.450 500.000 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 496.000 670.590 500.000 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 496.000 674.730 500.000 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 496.000 679.330 500.000 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 496.000 683.470 500.000 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 496.000 687.610 500.000 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 496.000 691.750 500.000 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 496.000 695.890 500.000 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 496.000 543.630 500.000 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 496.000 700.490 500.000 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 496.000 704.630 500.000 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 496.000 708.770 500.000 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 496.000 712.910 500.000 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 496.000 717.050 500.000 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 496.000 721.650 500.000 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 496.000 725.790 500.000 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 496.000 729.930 500.000 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 496.000 734.070 500.000 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 496.000 738.210 500.000 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 496.000 547.770 500.000 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 496.000 742.810 500.000 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 496.000 746.950 500.000 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 496.000 751.090 500.000 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 496.000 755.230 500.000 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 496.000 759.370 500.000 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 496.000 763.970 500.000 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 496.000 768.110 500.000 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 496.000 772.250 500.000 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 496.000 776.390 500.000 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 496.000 780.530 500.000 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 496.000 552.370 500.000 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 496.000 785.130 500.000 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 496.000 789.270 500.000 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 496.000 793.410 500.000 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 496.000 797.550 500.000 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 496.000 556.510 500.000 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 496.000 560.650 500.000 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 496.000 564.790 500.000 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 496.000 568.930 500.000 ;
    END
  END dout1[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 257.760 800.000 258.360 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 272.720 800.000 273.320 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 356.360 800.000 356.960 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 363.840 800.000 364.440 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 371.320 800.000 371.920 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 378.800 800.000 379.400 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 386.280 800.000 386.880 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 393.760 800.000 394.360 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 401.240 800.000 401.840 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 408.720 800.000 409.320 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 416.200 800.000 416.800 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 423.680 800.000 424.280 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 282.240 800.000 282.840 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 431.160 800.000 431.760 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 438.640 800.000 439.240 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 445.440 800.000 446.040 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 452.920 800.000 453.520 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 292.440 800.000 293.040 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 301.960 800.000 302.560 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 312.160 800.000 312.760 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 319.640 800.000 320.240 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 327.120 800.000 327.720 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 334.600 800.000 335.200 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 342.080 800.000 342.680 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 349.560 800.000 350.160 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 260.480 800.000 261.080 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 274.760 800.000 275.360 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 359.080 800.000 359.680 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 366.560 800.000 367.160 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 374.040 800.000 374.640 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 381.520 800.000 382.120 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 389.000 800.000 389.600 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 396.480 800.000 397.080 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 403.960 800.000 404.560 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 411.440 800.000 412.040 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 418.240 800.000 418.840 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.720 800.000 426.320 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 284.960 800.000 285.560 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 433.200 800.000 433.800 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 440.680 800.000 441.280 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 448.160 800.000 448.760 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 455.640 800.000 456.240 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 460.400 800.000 461.000 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 465.840 800.000 466.440 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 470.600 800.000 471.200 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 475.360 800.000 475.960 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 480.120 800.000 480.720 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 485.560 800.000 486.160 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 294.480 800.000 295.080 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 490.320 800.000 490.920 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 495.080 800.000 495.680 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 304.680 800.000 305.280 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 314.880 800.000 315.480 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 322.360 800.000 322.960 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 329.160 800.000 329.760 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 336.640 800.000 337.240 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 344.120 800.000 344.720 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 351.600 800.000 352.200 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 277.480 800.000 278.080 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 361.800 800.000 362.400 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 369.280 800.000 369.880 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 376.760 800.000 377.360 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 383.560 800.000 384.160 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 391.040 800.000 391.640 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 398.520 800.000 399.120 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 406.000 800.000 406.600 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 413.480 800.000 414.080 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 420.960 800.000 421.560 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 428.440 800.000 429.040 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 287.680 800.000 288.280 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 435.920 800.000 436.520 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 443.400 800.000 444.000 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 450.880 800.000 451.480 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 458.360 800.000 458.960 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 463.120 800.000 463.720 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 467.880 800.000 468.480 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 472.640 800.000 473.240 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 478.080 800.000 478.680 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 482.840 800.000 483.440 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 487.600 800.000 488.200 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 297.200 800.000 297.800 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.040 800.000 493.640 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 497.800 800.000 498.400 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 307.400 800.000 308.000 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.920 800.000 317.520 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 324.400 800.000 325.000 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 331.880 800.000 332.480 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 339.360 800.000 339.960 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 346.840 800.000 347.440 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 354.320 800.000 354.920 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 262.520 800.000 263.120 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 280.200 800.000 280.800 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 289.720 800.000 290.320 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.920 800.000 300.520 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 309.440 800.000 310.040 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 265.240 800.000 265.840 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 267.280 800.000 267.880 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 270.000 800.000 270.600 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 0.000 605.270 4.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 0.000 625.510 4.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END partID[9]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END probe_errorCode[1]
  PIN probe_errorCode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END probe_errorCode[2]
  PIN probe_errorCode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END probe_errorCode[3]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 487.120 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 0.720 800.000 1.320 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 2.760 800.000 3.360 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 496.000 14.630 500.000 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 496.000 18.770 500.000 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 496.000 23.370 500.000 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 496.000 27.510 500.000 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 496.000 31.650 500.000 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 486.965 ;
      LAYER met1 ;
        RECT 1.910 6.500 794.420 490.240 ;
      LAYER met2 ;
        RECT 2.490 495.720 5.790 498.285 ;
        RECT 6.630 495.720 9.930 498.285 ;
        RECT 10.770 495.720 14.070 498.285 ;
        RECT 14.910 495.720 18.210 498.285 ;
        RECT 19.050 495.720 22.810 498.285 ;
        RECT 23.650 495.720 26.950 498.285 ;
        RECT 27.790 495.720 31.090 498.285 ;
        RECT 31.930 495.720 35.230 498.285 ;
        RECT 36.070 495.720 39.370 498.285 ;
        RECT 40.210 495.720 43.970 498.285 ;
        RECT 44.810 495.720 48.110 498.285 ;
        RECT 48.950 495.720 52.250 498.285 ;
        RECT 53.090 495.720 56.390 498.285 ;
        RECT 57.230 495.720 60.530 498.285 ;
        RECT 61.370 495.720 65.130 498.285 ;
        RECT 65.970 495.720 69.270 498.285 ;
        RECT 70.110 495.720 73.410 498.285 ;
        RECT 74.250 495.720 77.550 498.285 ;
        RECT 78.390 495.720 81.690 498.285 ;
        RECT 82.530 495.720 86.290 498.285 ;
        RECT 87.130 495.720 90.430 498.285 ;
        RECT 91.270 495.720 94.570 498.285 ;
        RECT 95.410 495.720 98.710 498.285 ;
        RECT 99.550 495.720 102.850 498.285 ;
        RECT 103.690 495.720 107.450 498.285 ;
        RECT 108.290 495.720 111.590 498.285 ;
        RECT 112.430 495.720 115.730 498.285 ;
        RECT 116.570 495.720 119.870 498.285 ;
        RECT 120.710 495.720 124.010 498.285 ;
        RECT 124.850 495.720 128.610 498.285 ;
        RECT 129.450 495.720 132.750 498.285 ;
        RECT 133.590 495.720 136.890 498.285 ;
        RECT 137.730 495.720 141.030 498.285 ;
        RECT 141.870 495.720 145.170 498.285 ;
        RECT 146.010 495.720 149.770 498.285 ;
        RECT 150.610 495.720 153.910 498.285 ;
        RECT 154.750 495.720 158.050 498.285 ;
        RECT 158.890 495.720 162.190 498.285 ;
        RECT 163.030 495.720 166.330 498.285 ;
        RECT 167.170 495.720 170.930 498.285 ;
        RECT 171.770 495.720 175.070 498.285 ;
        RECT 175.910 495.720 179.210 498.285 ;
        RECT 180.050 495.720 183.350 498.285 ;
        RECT 184.190 495.720 187.490 498.285 ;
        RECT 188.330 495.720 192.090 498.285 ;
        RECT 192.930 495.720 196.230 498.285 ;
        RECT 197.070 495.720 200.370 498.285 ;
        RECT 201.210 495.720 204.510 498.285 ;
        RECT 205.350 495.720 208.650 498.285 ;
        RECT 209.490 495.720 213.250 498.285 ;
        RECT 214.090 495.720 217.390 498.285 ;
        RECT 218.230 495.720 221.530 498.285 ;
        RECT 222.370 495.720 225.670 498.285 ;
        RECT 226.510 495.720 229.810 498.285 ;
        RECT 230.650 495.720 234.410 498.285 ;
        RECT 235.250 495.720 238.550 498.285 ;
        RECT 239.390 495.720 242.690 498.285 ;
        RECT 243.530 495.720 246.830 498.285 ;
        RECT 247.670 495.720 250.970 498.285 ;
        RECT 251.810 495.720 255.570 498.285 ;
        RECT 256.410 495.720 259.710 498.285 ;
        RECT 260.550 495.720 263.850 498.285 ;
        RECT 264.690 495.720 267.990 498.285 ;
        RECT 268.830 495.720 272.130 498.285 ;
        RECT 272.970 495.720 276.730 498.285 ;
        RECT 277.570 495.720 280.870 498.285 ;
        RECT 281.710 495.720 285.010 498.285 ;
        RECT 285.850 495.720 289.150 498.285 ;
        RECT 289.990 495.720 293.290 498.285 ;
        RECT 294.130 495.720 297.890 498.285 ;
        RECT 298.730 495.720 302.030 498.285 ;
        RECT 302.870 495.720 306.170 498.285 ;
        RECT 307.010 495.720 310.310 498.285 ;
        RECT 311.150 495.720 314.450 498.285 ;
        RECT 315.290 495.720 319.050 498.285 ;
        RECT 319.890 495.720 323.190 498.285 ;
        RECT 324.030 495.720 327.330 498.285 ;
        RECT 328.170 495.720 331.470 498.285 ;
        RECT 332.310 495.720 335.610 498.285 ;
        RECT 336.450 495.720 340.210 498.285 ;
        RECT 341.050 495.720 344.350 498.285 ;
        RECT 345.190 495.720 348.490 498.285 ;
        RECT 349.330 495.720 352.630 498.285 ;
        RECT 353.470 495.720 356.770 498.285 ;
        RECT 357.610 495.720 361.370 498.285 ;
        RECT 362.210 495.720 365.510 498.285 ;
        RECT 366.350 495.720 369.650 498.285 ;
        RECT 370.490 495.720 373.790 498.285 ;
        RECT 374.630 495.720 377.930 498.285 ;
        RECT 378.770 495.720 382.530 498.285 ;
        RECT 383.370 495.720 386.670 498.285 ;
        RECT 387.510 495.720 390.810 498.285 ;
        RECT 391.650 495.720 394.950 498.285 ;
        RECT 395.790 495.720 399.090 498.285 ;
        RECT 399.930 495.720 403.690 498.285 ;
        RECT 404.530 495.720 407.830 498.285 ;
        RECT 408.670 495.720 411.970 498.285 ;
        RECT 412.810 495.720 416.110 498.285 ;
        RECT 416.950 495.720 420.250 498.285 ;
        RECT 421.090 495.720 424.850 498.285 ;
        RECT 425.690 495.720 428.990 498.285 ;
        RECT 429.830 495.720 433.130 498.285 ;
        RECT 433.970 495.720 437.270 498.285 ;
        RECT 438.110 495.720 441.410 498.285 ;
        RECT 442.250 495.720 446.010 498.285 ;
        RECT 446.850 495.720 450.150 498.285 ;
        RECT 450.990 495.720 454.290 498.285 ;
        RECT 455.130 495.720 458.430 498.285 ;
        RECT 459.270 495.720 462.570 498.285 ;
        RECT 463.410 495.720 467.170 498.285 ;
        RECT 468.010 495.720 471.310 498.285 ;
        RECT 472.150 495.720 475.450 498.285 ;
        RECT 476.290 495.720 479.590 498.285 ;
        RECT 480.430 495.720 483.730 498.285 ;
        RECT 484.570 495.720 488.330 498.285 ;
        RECT 489.170 495.720 492.470 498.285 ;
        RECT 493.310 495.720 496.610 498.285 ;
        RECT 497.450 495.720 500.750 498.285 ;
        RECT 501.590 495.720 504.890 498.285 ;
        RECT 505.730 495.720 509.490 498.285 ;
        RECT 510.330 495.720 513.630 498.285 ;
        RECT 514.470 495.720 517.770 498.285 ;
        RECT 518.610 495.720 521.910 498.285 ;
        RECT 522.750 495.720 526.050 498.285 ;
        RECT 526.890 495.720 530.650 498.285 ;
        RECT 531.490 495.720 534.790 498.285 ;
        RECT 535.630 495.720 538.930 498.285 ;
        RECT 539.770 495.720 543.070 498.285 ;
        RECT 543.910 495.720 547.210 498.285 ;
        RECT 548.050 495.720 551.810 498.285 ;
        RECT 552.650 495.720 555.950 498.285 ;
        RECT 556.790 495.720 560.090 498.285 ;
        RECT 560.930 495.720 564.230 498.285 ;
        RECT 565.070 495.720 568.370 498.285 ;
        RECT 569.210 495.720 572.970 498.285 ;
        RECT 573.810 495.720 577.110 498.285 ;
        RECT 577.950 495.720 581.250 498.285 ;
        RECT 582.090 495.720 585.390 498.285 ;
        RECT 586.230 495.720 589.530 498.285 ;
        RECT 590.370 495.720 594.130 498.285 ;
        RECT 594.970 495.720 598.270 498.285 ;
        RECT 599.110 495.720 602.410 498.285 ;
        RECT 603.250 495.720 606.550 498.285 ;
        RECT 607.390 495.720 610.690 498.285 ;
        RECT 611.530 495.720 615.290 498.285 ;
        RECT 616.130 495.720 619.430 498.285 ;
        RECT 620.270 495.720 623.570 498.285 ;
        RECT 624.410 495.720 627.710 498.285 ;
        RECT 628.550 495.720 631.850 498.285 ;
        RECT 632.690 495.720 636.450 498.285 ;
        RECT 637.290 495.720 640.590 498.285 ;
        RECT 641.430 495.720 644.730 498.285 ;
        RECT 645.570 495.720 648.870 498.285 ;
        RECT 649.710 495.720 653.010 498.285 ;
        RECT 653.850 495.720 657.610 498.285 ;
        RECT 658.450 495.720 661.750 498.285 ;
        RECT 662.590 495.720 665.890 498.285 ;
        RECT 666.730 495.720 670.030 498.285 ;
        RECT 670.870 495.720 674.170 498.285 ;
        RECT 675.010 495.720 678.770 498.285 ;
        RECT 679.610 495.720 682.910 498.285 ;
        RECT 683.750 495.720 687.050 498.285 ;
        RECT 687.890 495.720 691.190 498.285 ;
        RECT 692.030 495.720 695.330 498.285 ;
        RECT 696.170 495.720 699.930 498.285 ;
        RECT 700.770 495.720 704.070 498.285 ;
        RECT 704.910 495.720 708.210 498.285 ;
        RECT 709.050 495.720 712.350 498.285 ;
        RECT 713.190 495.720 716.490 498.285 ;
        RECT 717.330 495.720 721.090 498.285 ;
        RECT 721.930 495.720 725.230 498.285 ;
        RECT 726.070 495.720 729.370 498.285 ;
        RECT 730.210 495.720 733.510 498.285 ;
        RECT 734.350 495.720 737.650 498.285 ;
        RECT 738.490 495.720 742.250 498.285 ;
        RECT 743.090 495.720 746.390 498.285 ;
        RECT 747.230 495.720 750.530 498.285 ;
        RECT 751.370 495.720 754.670 498.285 ;
        RECT 755.510 495.720 758.810 498.285 ;
        RECT 759.650 495.720 763.410 498.285 ;
        RECT 764.250 495.720 767.550 498.285 ;
        RECT 768.390 495.720 771.690 498.285 ;
        RECT 772.530 495.720 775.830 498.285 ;
        RECT 776.670 495.720 779.970 498.285 ;
        RECT 780.810 495.720 784.570 498.285 ;
        RECT 785.410 495.720 788.710 498.285 ;
        RECT 789.550 495.720 792.490 498.285 ;
        RECT 1.940 4.280 792.490 495.720 ;
        RECT 1.940 0.835 9.930 4.280 ;
        RECT 10.770 0.835 30.170 4.280 ;
        RECT 31.010 0.835 50.870 4.280 ;
        RECT 51.710 0.835 71.110 4.280 ;
        RECT 71.950 0.835 91.810 4.280 ;
        RECT 92.650 0.835 112.050 4.280 ;
        RECT 112.890 0.835 132.750 4.280 ;
        RECT 133.590 0.835 153.450 4.280 ;
        RECT 154.290 0.835 173.690 4.280 ;
        RECT 174.530 0.835 194.390 4.280 ;
        RECT 195.230 0.835 214.630 4.280 ;
        RECT 215.470 0.835 235.330 4.280 ;
        RECT 236.170 0.835 256.030 4.280 ;
        RECT 256.870 0.835 276.270 4.280 ;
        RECT 277.110 0.835 296.970 4.280 ;
        RECT 297.810 0.835 317.210 4.280 ;
        RECT 318.050 0.835 337.910 4.280 ;
        RECT 338.750 0.835 358.610 4.280 ;
        RECT 359.450 0.835 378.850 4.280 ;
        RECT 379.690 0.835 399.550 4.280 ;
        RECT 400.390 0.835 419.790 4.280 ;
        RECT 420.630 0.835 440.490 4.280 ;
        RECT 441.330 0.835 460.730 4.280 ;
        RECT 461.570 0.835 481.430 4.280 ;
        RECT 482.270 0.835 502.130 4.280 ;
        RECT 502.970 0.835 522.370 4.280 ;
        RECT 523.210 0.835 543.070 4.280 ;
        RECT 543.910 0.835 563.310 4.280 ;
        RECT 564.150 0.835 584.010 4.280 ;
        RECT 584.850 0.835 604.710 4.280 ;
        RECT 605.550 0.835 624.950 4.280 ;
        RECT 625.790 0.835 645.650 4.280 ;
        RECT 646.490 0.835 665.890 4.280 ;
        RECT 666.730 0.835 686.590 4.280 ;
        RECT 687.430 0.835 707.290 4.280 ;
        RECT 708.130 0.835 727.530 4.280 ;
        RECT 728.370 0.835 748.230 4.280 ;
        RECT 749.070 0.835 768.470 4.280 ;
        RECT 769.310 0.835 789.170 4.280 ;
        RECT 790.010 0.835 792.490 4.280 ;
      LAYER met3 ;
        RECT 4.000 497.400 795.600 498.265 ;
        RECT 4.000 496.080 796.000 497.400 ;
        RECT 4.400 494.680 795.600 496.080 ;
        RECT 4.000 494.040 796.000 494.680 ;
        RECT 4.000 492.640 795.600 494.040 ;
        RECT 4.000 491.320 796.000 492.640 ;
        RECT 4.000 489.920 795.600 491.320 ;
        RECT 4.000 488.600 796.000 489.920 ;
        RECT 4.000 487.920 795.600 488.600 ;
        RECT 4.400 487.200 795.600 487.920 ;
        RECT 4.400 486.560 796.000 487.200 ;
        RECT 4.400 486.520 795.600 486.560 ;
        RECT 4.000 485.160 795.600 486.520 ;
        RECT 4.000 483.840 796.000 485.160 ;
        RECT 4.000 482.440 795.600 483.840 ;
        RECT 4.000 481.120 796.000 482.440 ;
        RECT 4.000 479.720 795.600 481.120 ;
        RECT 4.000 479.080 796.000 479.720 ;
        RECT 4.400 477.680 795.600 479.080 ;
        RECT 4.000 476.360 796.000 477.680 ;
        RECT 4.000 474.960 795.600 476.360 ;
        RECT 4.000 473.640 796.000 474.960 ;
        RECT 4.000 472.240 795.600 473.640 ;
        RECT 4.000 471.600 796.000 472.240 ;
        RECT 4.000 470.920 795.600 471.600 ;
        RECT 4.400 470.200 795.600 470.920 ;
        RECT 4.400 469.520 796.000 470.200 ;
        RECT 4.000 468.880 796.000 469.520 ;
        RECT 4.000 467.480 795.600 468.880 ;
        RECT 4.000 466.840 796.000 467.480 ;
        RECT 4.000 465.440 795.600 466.840 ;
        RECT 4.000 464.120 796.000 465.440 ;
        RECT 4.000 462.720 795.600 464.120 ;
        RECT 4.000 462.080 796.000 462.720 ;
        RECT 4.400 461.400 796.000 462.080 ;
        RECT 4.400 460.680 795.600 461.400 ;
        RECT 4.000 460.000 795.600 460.680 ;
        RECT 4.000 459.360 796.000 460.000 ;
        RECT 4.000 457.960 795.600 459.360 ;
        RECT 4.000 456.640 796.000 457.960 ;
        RECT 4.000 455.240 795.600 456.640 ;
        RECT 4.000 453.920 796.000 455.240 ;
        RECT 4.400 452.520 795.600 453.920 ;
        RECT 4.000 451.880 796.000 452.520 ;
        RECT 4.000 450.480 795.600 451.880 ;
        RECT 4.000 449.160 796.000 450.480 ;
        RECT 4.000 447.760 795.600 449.160 ;
        RECT 4.000 446.440 796.000 447.760 ;
        RECT 4.000 445.080 795.600 446.440 ;
        RECT 4.400 445.040 795.600 445.080 ;
        RECT 4.400 444.400 796.000 445.040 ;
        RECT 4.400 443.680 795.600 444.400 ;
        RECT 4.000 443.000 795.600 443.680 ;
        RECT 4.000 441.680 796.000 443.000 ;
        RECT 4.000 440.280 795.600 441.680 ;
        RECT 4.000 439.640 796.000 440.280 ;
        RECT 4.000 438.240 795.600 439.640 ;
        RECT 4.000 436.920 796.000 438.240 ;
        RECT 4.400 435.520 795.600 436.920 ;
        RECT 4.000 434.200 796.000 435.520 ;
        RECT 4.000 432.800 795.600 434.200 ;
        RECT 4.000 432.160 796.000 432.800 ;
        RECT 4.000 430.760 795.600 432.160 ;
        RECT 4.000 429.440 796.000 430.760 ;
        RECT 4.000 428.080 795.600 429.440 ;
        RECT 4.400 428.040 795.600 428.080 ;
        RECT 4.400 426.720 796.000 428.040 ;
        RECT 4.400 426.680 795.600 426.720 ;
        RECT 4.000 425.320 795.600 426.680 ;
        RECT 4.000 424.680 796.000 425.320 ;
        RECT 4.000 423.280 795.600 424.680 ;
        RECT 4.000 421.960 796.000 423.280 ;
        RECT 4.000 420.560 795.600 421.960 ;
        RECT 4.000 419.920 796.000 420.560 ;
        RECT 4.400 419.240 796.000 419.920 ;
        RECT 4.400 418.520 795.600 419.240 ;
        RECT 4.000 417.840 795.600 418.520 ;
        RECT 4.000 417.200 796.000 417.840 ;
        RECT 4.000 415.800 795.600 417.200 ;
        RECT 4.000 414.480 796.000 415.800 ;
        RECT 4.000 413.080 795.600 414.480 ;
        RECT 4.000 412.440 796.000 413.080 ;
        RECT 4.000 411.080 795.600 412.440 ;
        RECT 4.400 411.040 795.600 411.080 ;
        RECT 4.400 409.720 796.000 411.040 ;
        RECT 4.400 409.680 795.600 409.720 ;
        RECT 4.000 408.320 795.600 409.680 ;
        RECT 4.000 407.000 796.000 408.320 ;
        RECT 4.000 405.600 795.600 407.000 ;
        RECT 4.000 404.960 796.000 405.600 ;
        RECT 4.000 403.560 795.600 404.960 ;
        RECT 4.000 402.920 796.000 403.560 ;
        RECT 4.400 402.240 796.000 402.920 ;
        RECT 4.400 401.520 795.600 402.240 ;
        RECT 4.000 400.840 795.600 401.520 ;
        RECT 4.000 399.520 796.000 400.840 ;
        RECT 4.000 398.120 795.600 399.520 ;
        RECT 4.000 397.480 796.000 398.120 ;
        RECT 4.000 396.080 795.600 397.480 ;
        RECT 4.000 394.760 796.000 396.080 ;
        RECT 4.400 393.360 795.600 394.760 ;
        RECT 4.000 392.040 796.000 393.360 ;
        RECT 4.000 390.640 795.600 392.040 ;
        RECT 4.000 390.000 796.000 390.640 ;
        RECT 4.000 388.600 795.600 390.000 ;
        RECT 4.000 387.280 796.000 388.600 ;
        RECT 4.000 385.920 795.600 387.280 ;
        RECT 4.400 385.880 795.600 385.920 ;
        RECT 4.400 384.560 796.000 385.880 ;
        RECT 4.400 384.520 795.600 384.560 ;
        RECT 4.000 383.160 795.600 384.520 ;
        RECT 4.000 382.520 796.000 383.160 ;
        RECT 4.000 381.120 795.600 382.520 ;
        RECT 4.000 379.800 796.000 381.120 ;
        RECT 4.000 378.400 795.600 379.800 ;
        RECT 4.000 377.760 796.000 378.400 ;
        RECT 4.400 376.360 795.600 377.760 ;
        RECT 4.000 375.040 796.000 376.360 ;
        RECT 4.000 373.640 795.600 375.040 ;
        RECT 4.000 372.320 796.000 373.640 ;
        RECT 4.000 370.920 795.600 372.320 ;
        RECT 4.000 370.280 796.000 370.920 ;
        RECT 4.000 368.920 795.600 370.280 ;
        RECT 4.400 368.880 795.600 368.920 ;
        RECT 4.400 367.560 796.000 368.880 ;
        RECT 4.400 367.520 795.600 367.560 ;
        RECT 4.000 366.160 795.600 367.520 ;
        RECT 4.000 364.840 796.000 366.160 ;
        RECT 4.000 363.440 795.600 364.840 ;
        RECT 4.000 362.800 796.000 363.440 ;
        RECT 4.000 361.400 795.600 362.800 ;
        RECT 4.000 360.760 796.000 361.400 ;
        RECT 4.400 360.080 796.000 360.760 ;
        RECT 4.400 359.360 795.600 360.080 ;
        RECT 4.000 358.680 795.600 359.360 ;
        RECT 4.000 357.360 796.000 358.680 ;
        RECT 4.000 355.960 795.600 357.360 ;
        RECT 4.000 355.320 796.000 355.960 ;
        RECT 4.000 353.920 795.600 355.320 ;
        RECT 4.000 352.600 796.000 353.920 ;
        RECT 4.000 351.920 795.600 352.600 ;
        RECT 4.400 351.200 795.600 351.920 ;
        RECT 4.400 350.560 796.000 351.200 ;
        RECT 4.400 350.520 795.600 350.560 ;
        RECT 4.000 349.160 795.600 350.520 ;
        RECT 4.000 347.840 796.000 349.160 ;
        RECT 4.000 346.440 795.600 347.840 ;
        RECT 4.000 345.120 796.000 346.440 ;
        RECT 4.000 343.760 795.600 345.120 ;
        RECT 4.400 343.720 795.600 343.760 ;
        RECT 4.400 343.080 796.000 343.720 ;
        RECT 4.400 342.360 795.600 343.080 ;
        RECT 4.000 341.680 795.600 342.360 ;
        RECT 4.000 340.360 796.000 341.680 ;
        RECT 4.000 338.960 795.600 340.360 ;
        RECT 4.000 337.640 796.000 338.960 ;
        RECT 4.000 336.240 795.600 337.640 ;
        RECT 4.000 335.600 796.000 336.240 ;
        RECT 4.000 334.920 795.600 335.600 ;
        RECT 4.400 334.200 795.600 334.920 ;
        RECT 4.400 333.520 796.000 334.200 ;
        RECT 4.000 332.880 796.000 333.520 ;
        RECT 4.000 331.480 795.600 332.880 ;
        RECT 4.000 330.160 796.000 331.480 ;
        RECT 4.000 328.760 795.600 330.160 ;
        RECT 4.000 328.120 796.000 328.760 ;
        RECT 4.000 326.760 795.600 328.120 ;
        RECT 4.400 326.720 795.600 326.760 ;
        RECT 4.400 325.400 796.000 326.720 ;
        RECT 4.400 325.360 795.600 325.400 ;
        RECT 4.000 324.000 795.600 325.360 ;
        RECT 4.000 323.360 796.000 324.000 ;
        RECT 4.000 321.960 795.600 323.360 ;
        RECT 4.000 320.640 796.000 321.960 ;
        RECT 4.000 319.240 795.600 320.640 ;
        RECT 4.000 317.920 796.000 319.240 ;
        RECT 4.400 316.520 795.600 317.920 ;
        RECT 4.000 315.880 796.000 316.520 ;
        RECT 4.000 314.480 795.600 315.880 ;
        RECT 4.000 313.160 796.000 314.480 ;
        RECT 4.000 311.760 795.600 313.160 ;
        RECT 4.000 310.440 796.000 311.760 ;
        RECT 4.000 309.760 795.600 310.440 ;
        RECT 4.400 309.040 795.600 309.760 ;
        RECT 4.400 308.400 796.000 309.040 ;
        RECT 4.400 308.360 795.600 308.400 ;
        RECT 4.000 307.000 795.600 308.360 ;
        RECT 4.000 305.680 796.000 307.000 ;
        RECT 4.000 304.280 795.600 305.680 ;
        RECT 4.000 302.960 796.000 304.280 ;
        RECT 4.000 301.600 795.600 302.960 ;
        RECT 4.400 301.560 795.600 301.600 ;
        RECT 4.400 300.920 796.000 301.560 ;
        RECT 4.400 300.200 795.600 300.920 ;
        RECT 4.000 299.520 795.600 300.200 ;
        RECT 4.000 298.200 796.000 299.520 ;
        RECT 4.000 296.800 795.600 298.200 ;
        RECT 4.000 295.480 796.000 296.800 ;
        RECT 4.000 294.080 795.600 295.480 ;
        RECT 4.000 293.440 796.000 294.080 ;
        RECT 4.000 292.760 795.600 293.440 ;
        RECT 4.400 292.040 795.600 292.760 ;
        RECT 4.400 291.360 796.000 292.040 ;
        RECT 4.000 290.720 796.000 291.360 ;
        RECT 4.000 289.320 795.600 290.720 ;
        RECT 4.000 288.680 796.000 289.320 ;
        RECT 4.000 287.280 795.600 288.680 ;
        RECT 4.000 285.960 796.000 287.280 ;
        RECT 4.000 284.600 795.600 285.960 ;
        RECT 4.400 284.560 795.600 284.600 ;
        RECT 4.400 283.240 796.000 284.560 ;
        RECT 4.400 283.200 795.600 283.240 ;
        RECT 4.000 281.840 795.600 283.200 ;
        RECT 4.000 281.200 796.000 281.840 ;
        RECT 4.000 279.800 795.600 281.200 ;
        RECT 4.000 278.480 796.000 279.800 ;
        RECT 4.000 277.080 795.600 278.480 ;
        RECT 4.000 275.760 796.000 277.080 ;
        RECT 4.400 274.360 795.600 275.760 ;
        RECT 4.000 273.720 796.000 274.360 ;
        RECT 4.000 272.320 795.600 273.720 ;
        RECT 4.000 271.000 796.000 272.320 ;
        RECT 4.000 269.600 795.600 271.000 ;
        RECT 4.000 268.280 796.000 269.600 ;
        RECT 4.000 267.600 795.600 268.280 ;
        RECT 4.400 266.880 795.600 267.600 ;
        RECT 4.400 266.240 796.000 266.880 ;
        RECT 4.400 266.200 795.600 266.240 ;
        RECT 4.000 264.840 795.600 266.200 ;
        RECT 4.000 263.520 796.000 264.840 ;
        RECT 4.000 262.120 795.600 263.520 ;
        RECT 4.000 261.480 796.000 262.120 ;
        RECT 4.000 260.080 795.600 261.480 ;
        RECT 4.000 258.760 796.000 260.080 ;
        RECT 4.400 257.360 795.600 258.760 ;
        RECT 4.000 256.040 796.000 257.360 ;
        RECT 4.000 254.640 795.600 256.040 ;
        RECT 4.000 254.000 796.000 254.640 ;
        RECT 4.000 252.600 795.600 254.000 ;
        RECT 4.000 251.280 796.000 252.600 ;
        RECT 4.000 250.600 795.600 251.280 ;
        RECT 4.400 249.880 795.600 250.600 ;
        RECT 4.400 249.200 796.000 249.880 ;
        RECT 4.000 248.560 796.000 249.200 ;
        RECT 4.000 247.160 795.600 248.560 ;
        RECT 4.000 246.520 796.000 247.160 ;
        RECT 4.000 245.120 795.600 246.520 ;
        RECT 4.000 243.800 796.000 245.120 ;
        RECT 4.000 242.400 795.600 243.800 ;
        RECT 4.000 241.760 796.000 242.400 ;
        RECT 4.400 241.080 796.000 241.760 ;
        RECT 4.400 240.360 795.600 241.080 ;
        RECT 4.000 239.680 795.600 240.360 ;
        RECT 4.000 239.040 796.000 239.680 ;
        RECT 4.000 237.640 795.600 239.040 ;
        RECT 4.000 236.320 796.000 237.640 ;
        RECT 4.000 234.920 795.600 236.320 ;
        RECT 4.000 234.280 796.000 234.920 ;
        RECT 4.000 233.600 795.600 234.280 ;
        RECT 4.400 232.880 795.600 233.600 ;
        RECT 4.400 232.200 796.000 232.880 ;
        RECT 4.000 231.560 796.000 232.200 ;
        RECT 4.000 230.160 795.600 231.560 ;
        RECT 4.000 228.840 796.000 230.160 ;
        RECT 4.000 227.440 795.600 228.840 ;
        RECT 4.000 226.800 796.000 227.440 ;
        RECT 4.000 225.400 795.600 226.800 ;
        RECT 4.000 224.760 796.000 225.400 ;
        RECT 4.400 224.080 796.000 224.760 ;
        RECT 4.400 223.360 795.600 224.080 ;
        RECT 4.000 222.680 795.600 223.360 ;
        RECT 4.000 221.360 796.000 222.680 ;
        RECT 4.000 219.960 795.600 221.360 ;
        RECT 4.000 219.320 796.000 219.960 ;
        RECT 4.000 217.920 795.600 219.320 ;
        RECT 4.000 216.600 796.000 217.920 ;
        RECT 4.400 215.200 795.600 216.600 ;
        RECT 4.000 213.880 796.000 215.200 ;
        RECT 4.000 212.480 795.600 213.880 ;
        RECT 4.000 211.840 796.000 212.480 ;
        RECT 4.000 210.440 795.600 211.840 ;
        RECT 4.000 209.120 796.000 210.440 ;
        RECT 4.000 207.760 795.600 209.120 ;
        RECT 4.400 207.720 795.600 207.760 ;
        RECT 4.400 207.080 796.000 207.720 ;
        RECT 4.400 206.360 795.600 207.080 ;
        RECT 4.000 205.680 795.600 206.360 ;
        RECT 4.000 204.360 796.000 205.680 ;
        RECT 4.000 202.960 795.600 204.360 ;
        RECT 4.000 201.640 796.000 202.960 ;
        RECT 4.000 200.240 795.600 201.640 ;
        RECT 4.000 199.600 796.000 200.240 ;
        RECT 4.400 198.200 795.600 199.600 ;
        RECT 4.000 196.880 796.000 198.200 ;
        RECT 4.000 195.480 795.600 196.880 ;
        RECT 4.000 194.160 796.000 195.480 ;
        RECT 4.000 192.760 795.600 194.160 ;
        RECT 4.000 192.120 796.000 192.760 ;
        RECT 4.000 191.440 795.600 192.120 ;
        RECT 4.400 190.720 795.600 191.440 ;
        RECT 4.400 190.040 796.000 190.720 ;
        RECT 4.000 189.400 796.000 190.040 ;
        RECT 4.000 188.000 795.600 189.400 ;
        RECT 4.000 186.680 796.000 188.000 ;
        RECT 4.000 185.280 795.600 186.680 ;
        RECT 4.000 184.640 796.000 185.280 ;
        RECT 4.000 183.240 795.600 184.640 ;
        RECT 4.000 182.600 796.000 183.240 ;
        RECT 4.400 181.920 796.000 182.600 ;
        RECT 4.400 181.200 795.600 181.920 ;
        RECT 4.000 180.520 795.600 181.200 ;
        RECT 4.000 179.200 796.000 180.520 ;
        RECT 4.000 177.800 795.600 179.200 ;
        RECT 4.000 177.160 796.000 177.800 ;
        RECT 4.000 175.760 795.600 177.160 ;
        RECT 4.000 174.440 796.000 175.760 ;
        RECT 4.400 173.040 795.600 174.440 ;
        RECT 4.000 172.400 796.000 173.040 ;
        RECT 4.000 171.000 795.600 172.400 ;
        RECT 4.000 169.680 796.000 171.000 ;
        RECT 4.000 168.280 795.600 169.680 ;
        RECT 4.000 166.960 796.000 168.280 ;
        RECT 4.000 165.600 795.600 166.960 ;
        RECT 4.400 165.560 795.600 165.600 ;
        RECT 4.400 164.920 796.000 165.560 ;
        RECT 4.400 164.200 795.600 164.920 ;
        RECT 4.000 163.520 795.600 164.200 ;
        RECT 4.000 162.200 796.000 163.520 ;
        RECT 4.000 160.800 795.600 162.200 ;
        RECT 4.000 159.480 796.000 160.800 ;
        RECT 4.000 158.080 795.600 159.480 ;
        RECT 4.000 157.440 796.000 158.080 ;
        RECT 4.400 156.040 795.600 157.440 ;
        RECT 4.000 154.720 796.000 156.040 ;
        RECT 4.000 153.320 795.600 154.720 ;
        RECT 4.000 152.000 796.000 153.320 ;
        RECT 4.000 150.600 795.600 152.000 ;
        RECT 4.000 149.960 796.000 150.600 ;
        RECT 4.000 148.600 795.600 149.960 ;
        RECT 4.400 148.560 795.600 148.600 ;
        RECT 4.400 147.240 796.000 148.560 ;
        RECT 4.400 147.200 795.600 147.240 ;
        RECT 4.000 145.840 795.600 147.200 ;
        RECT 4.000 145.200 796.000 145.840 ;
        RECT 4.000 143.800 795.600 145.200 ;
        RECT 4.000 142.480 796.000 143.800 ;
        RECT 4.000 141.080 795.600 142.480 ;
        RECT 4.000 140.440 796.000 141.080 ;
        RECT 4.400 139.760 796.000 140.440 ;
        RECT 4.400 139.040 795.600 139.760 ;
        RECT 4.000 138.360 795.600 139.040 ;
        RECT 4.000 137.720 796.000 138.360 ;
        RECT 4.000 136.320 795.600 137.720 ;
        RECT 4.000 135.000 796.000 136.320 ;
        RECT 4.000 133.600 795.600 135.000 ;
        RECT 4.000 132.280 796.000 133.600 ;
        RECT 4.000 131.600 795.600 132.280 ;
        RECT 4.400 130.880 795.600 131.600 ;
        RECT 4.400 130.240 796.000 130.880 ;
        RECT 4.400 130.200 795.600 130.240 ;
        RECT 4.000 128.840 795.600 130.200 ;
        RECT 4.000 127.520 796.000 128.840 ;
        RECT 4.000 126.120 795.600 127.520 ;
        RECT 4.000 124.800 796.000 126.120 ;
        RECT 4.000 123.440 795.600 124.800 ;
        RECT 4.400 123.400 795.600 123.440 ;
        RECT 4.400 122.760 796.000 123.400 ;
        RECT 4.400 122.040 795.600 122.760 ;
        RECT 4.000 121.360 795.600 122.040 ;
        RECT 4.000 120.040 796.000 121.360 ;
        RECT 4.000 118.640 795.600 120.040 ;
        RECT 4.000 118.000 796.000 118.640 ;
        RECT 4.000 116.600 795.600 118.000 ;
        RECT 4.000 115.280 796.000 116.600 ;
        RECT 4.000 114.600 795.600 115.280 ;
        RECT 4.400 113.880 795.600 114.600 ;
        RECT 4.400 113.200 796.000 113.880 ;
        RECT 4.000 112.560 796.000 113.200 ;
        RECT 4.000 111.160 795.600 112.560 ;
        RECT 4.000 110.520 796.000 111.160 ;
        RECT 4.000 109.120 795.600 110.520 ;
        RECT 4.000 107.800 796.000 109.120 ;
        RECT 4.000 106.440 795.600 107.800 ;
        RECT 4.400 106.400 795.600 106.440 ;
        RECT 4.400 105.080 796.000 106.400 ;
        RECT 4.400 105.040 795.600 105.080 ;
        RECT 4.000 103.680 795.600 105.040 ;
        RECT 4.000 103.040 796.000 103.680 ;
        RECT 4.000 101.640 795.600 103.040 ;
        RECT 4.000 100.320 796.000 101.640 ;
        RECT 4.000 98.920 795.600 100.320 ;
        RECT 4.000 98.280 796.000 98.920 ;
        RECT 4.400 97.600 796.000 98.280 ;
        RECT 4.400 96.880 795.600 97.600 ;
        RECT 4.000 96.200 795.600 96.880 ;
        RECT 4.000 95.560 796.000 96.200 ;
        RECT 4.000 94.160 795.600 95.560 ;
        RECT 4.000 92.840 796.000 94.160 ;
        RECT 4.000 91.440 795.600 92.840 ;
        RECT 4.000 90.120 796.000 91.440 ;
        RECT 4.000 89.440 795.600 90.120 ;
        RECT 4.400 88.720 795.600 89.440 ;
        RECT 4.400 88.080 796.000 88.720 ;
        RECT 4.400 88.040 795.600 88.080 ;
        RECT 4.000 86.680 795.600 88.040 ;
        RECT 4.000 85.360 796.000 86.680 ;
        RECT 4.000 83.960 795.600 85.360 ;
        RECT 4.000 83.320 796.000 83.960 ;
        RECT 4.000 81.920 795.600 83.320 ;
        RECT 4.000 81.280 796.000 81.920 ;
        RECT 4.400 80.600 796.000 81.280 ;
        RECT 4.400 79.880 795.600 80.600 ;
        RECT 4.000 79.200 795.600 79.880 ;
        RECT 4.000 77.880 796.000 79.200 ;
        RECT 4.000 76.480 795.600 77.880 ;
        RECT 4.000 75.840 796.000 76.480 ;
        RECT 4.000 74.440 795.600 75.840 ;
        RECT 4.000 73.120 796.000 74.440 ;
        RECT 4.000 72.440 795.600 73.120 ;
        RECT 4.400 71.720 795.600 72.440 ;
        RECT 4.400 71.040 796.000 71.720 ;
        RECT 4.000 70.400 796.000 71.040 ;
        RECT 4.000 69.000 795.600 70.400 ;
        RECT 4.000 68.360 796.000 69.000 ;
        RECT 4.000 66.960 795.600 68.360 ;
        RECT 4.000 65.640 796.000 66.960 ;
        RECT 4.000 64.280 795.600 65.640 ;
        RECT 4.400 64.240 795.600 64.280 ;
        RECT 4.400 62.920 796.000 64.240 ;
        RECT 4.400 62.880 795.600 62.920 ;
        RECT 4.000 61.520 795.600 62.880 ;
        RECT 4.000 60.880 796.000 61.520 ;
        RECT 4.000 59.480 795.600 60.880 ;
        RECT 4.000 58.160 796.000 59.480 ;
        RECT 4.000 56.760 795.600 58.160 ;
        RECT 4.000 56.120 796.000 56.760 ;
        RECT 4.000 55.440 795.600 56.120 ;
        RECT 4.400 54.720 795.600 55.440 ;
        RECT 4.400 54.040 796.000 54.720 ;
        RECT 4.000 53.400 796.000 54.040 ;
        RECT 4.000 52.000 795.600 53.400 ;
        RECT 4.000 50.680 796.000 52.000 ;
        RECT 4.000 49.280 795.600 50.680 ;
        RECT 4.000 48.640 796.000 49.280 ;
        RECT 4.000 47.280 795.600 48.640 ;
        RECT 4.400 47.240 795.600 47.280 ;
        RECT 4.400 45.920 796.000 47.240 ;
        RECT 4.400 45.880 795.600 45.920 ;
        RECT 4.000 44.520 795.600 45.880 ;
        RECT 4.000 43.200 796.000 44.520 ;
        RECT 4.000 41.800 795.600 43.200 ;
        RECT 4.000 41.160 796.000 41.800 ;
        RECT 4.000 39.760 795.600 41.160 ;
        RECT 4.000 38.440 796.000 39.760 ;
        RECT 4.400 37.040 795.600 38.440 ;
        RECT 4.000 35.720 796.000 37.040 ;
        RECT 4.000 34.320 795.600 35.720 ;
        RECT 4.000 33.680 796.000 34.320 ;
        RECT 4.000 32.280 795.600 33.680 ;
        RECT 4.000 30.960 796.000 32.280 ;
        RECT 4.000 30.280 795.600 30.960 ;
        RECT 4.400 29.560 795.600 30.280 ;
        RECT 4.400 28.920 796.000 29.560 ;
        RECT 4.400 28.880 795.600 28.920 ;
        RECT 4.000 27.520 795.600 28.880 ;
        RECT 4.000 26.200 796.000 27.520 ;
        RECT 4.000 24.800 795.600 26.200 ;
        RECT 4.000 23.480 796.000 24.800 ;
        RECT 4.000 22.080 795.600 23.480 ;
        RECT 4.000 21.440 796.000 22.080 ;
        RECT 4.400 20.040 795.600 21.440 ;
        RECT 4.000 18.720 796.000 20.040 ;
        RECT 4.000 17.320 795.600 18.720 ;
        RECT 4.000 16.000 796.000 17.320 ;
        RECT 4.000 14.600 795.600 16.000 ;
        RECT 4.000 13.960 796.000 14.600 ;
        RECT 4.000 13.280 795.600 13.960 ;
        RECT 4.400 12.560 795.600 13.280 ;
        RECT 4.400 11.880 796.000 12.560 ;
        RECT 4.000 11.240 796.000 11.880 ;
        RECT 4.000 9.840 795.600 11.240 ;
        RECT 4.000 8.520 796.000 9.840 ;
        RECT 4.000 7.120 795.600 8.520 ;
        RECT 4.000 6.480 796.000 7.120 ;
        RECT 4.000 5.120 795.600 6.480 ;
        RECT 4.400 5.080 795.600 5.120 ;
        RECT 4.400 3.760 796.000 5.080 ;
        RECT 4.400 3.720 795.600 3.760 ;
        RECT 4.000 2.360 795.600 3.720 ;
        RECT 4.000 1.720 796.000 2.360 ;
        RECT 4.000 0.855 795.600 1.720 ;
      LAYER met4 ;
        RECT 778.615 440.815 778.945 462.905 ;
  END
END ExperiarCore
END LIBRARY

