magic
tech sky130A
magscale 1 2
timestamp 1654557799
<< obsli1 >>
rect 1104 2159 68816 97393
<< obsm1 >>
rect 290 1640 69722 97424
<< metal2 >>
rect 294 0 350 800
rect 846 0 902 800
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9126 0 9182 800
rect 9770 0 9826 800
rect 10414 0 10470 800
rect 11058 0 11114 800
rect 11702 0 11758 800
rect 12346 0 12402 800
rect 12990 0 13046 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 14922 0 14978 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23754 0 23810 800
rect 24398 0 24454 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26330 0 26386 800
rect 26974 0 27030 800
rect 27618 0 27674 800
rect 28262 0 28318 800
rect 28906 0 28962 800
rect 29550 0 29606 800
rect 30194 0 30250 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 32034 0 32090 800
rect 32678 0 32734 800
rect 33322 0 33378 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35898 0 35954 800
rect 36542 0 36598 800
rect 37186 0 37242 800
rect 37830 0 37886 800
rect 38474 0 38530 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40314 0 40370 800
rect 40958 0 41014 800
rect 41602 0 41658 800
rect 42246 0 42302 800
rect 42890 0 42946 800
rect 43534 0 43590 800
rect 44178 0 44234 800
rect 44822 0 44878 800
rect 45466 0 45522 800
rect 46110 0 46166 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47950 0 48006 800
rect 48594 0 48650 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51814 0 51870 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 54942 0 54998 800
rect 55586 0 55642 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57518 0 57574 800
rect 58162 0 58218 800
rect 58806 0 58862 800
rect 59450 0 59506 800
rect 60094 0 60150 800
rect 60738 0 60794 800
rect 61382 0 61438 800
rect 62026 0 62082 800
rect 62578 0 62634 800
rect 63222 0 63278 800
rect 63866 0 63922 800
rect 64510 0 64566 800
rect 65154 0 65210 800
rect 65798 0 65854 800
rect 66442 0 66498 800
rect 67086 0 67142 800
rect 67730 0 67786 800
rect 68374 0 68430 800
rect 69018 0 69074 800
rect 69662 0 69718 800
<< obsm2 >>
rect 296 856 69716 99657
rect 406 54 790 856
rect 958 54 1434 856
rect 1602 54 2078 856
rect 2246 54 2722 856
rect 2890 54 3366 856
rect 3534 54 4010 856
rect 4178 54 4654 856
rect 4822 54 5298 856
rect 5466 54 5942 856
rect 6110 54 6586 856
rect 6754 54 7230 856
rect 7398 54 7874 856
rect 8042 54 8426 856
rect 8594 54 9070 856
rect 9238 54 9714 856
rect 9882 54 10358 856
rect 10526 54 11002 856
rect 11170 54 11646 856
rect 11814 54 12290 856
rect 12458 54 12934 856
rect 13102 54 13578 856
rect 13746 54 14222 856
rect 14390 54 14866 856
rect 15034 54 15510 856
rect 15678 54 16062 856
rect 16230 54 16706 856
rect 16874 54 17350 856
rect 17518 54 17994 856
rect 18162 54 18638 856
rect 18806 54 19282 856
rect 19450 54 19926 856
rect 20094 54 20570 856
rect 20738 54 21214 856
rect 21382 54 21858 856
rect 22026 54 22502 856
rect 22670 54 23146 856
rect 23314 54 23698 856
rect 23866 54 24342 856
rect 24510 54 24986 856
rect 25154 54 25630 856
rect 25798 54 26274 856
rect 26442 54 26918 856
rect 27086 54 27562 856
rect 27730 54 28206 856
rect 28374 54 28850 856
rect 29018 54 29494 856
rect 29662 54 30138 856
rect 30306 54 30782 856
rect 30950 54 31334 856
rect 31502 54 31978 856
rect 32146 54 32622 856
rect 32790 54 33266 856
rect 33434 54 33910 856
rect 34078 54 34554 856
rect 34722 54 35198 856
rect 35366 54 35842 856
rect 36010 54 36486 856
rect 36654 54 37130 856
rect 37298 54 37774 856
rect 37942 54 38418 856
rect 38586 54 39062 856
rect 39230 54 39614 856
rect 39782 54 40258 856
rect 40426 54 40902 856
rect 41070 54 41546 856
rect 41714 54 42190 856
rect 42358 54 42834 856
rect 43002 54 43478 856
rect 43646 54 44122 856
rect 44290 54 44766 856
rect 44934 54 45410 856
rect 45578 54 46054 856
rect 46222 54 46698 856
rect 46866 54 47250 856
rect 47418 54 47894 856
rect 48062 54 48538 856
rect 48706 54 49182 856
rect 49350 54 49826 856
rect 49994 54 50470 856
rect 50638 54 51114 856
rect 51282 54 51758 856
rect 51926 54 52402 856
rect 52570 54 53046 856
rect 53214 54 53690 856
rect 53858 54 54334 856
rect 54502 54 54886 856
rect 55054 54 55530 856
rect 55698 54 56174 856
rect 56342 54 56818 856
rect 56986 54 57462 856
rect 57630 54 58106 856
rect 58274 54 58750 856
rect 58918 54 59394 856
rect 59562 54 60038 856
rect 60206 54 60682 856
rect 60850 54 61326 856
rect 61494 54 61970 856
rect 62138 54 62522 856
rect 62690 54 63166 856
rect 63334 54 63810 856
rect 63978 54 64454 856
rect 64622 54 65098 856
rect 65266 54 65742 856
rect 65910 54 66386 856
rect 66554 54 67030 856
rect 67198 54 67674 856
rect 67842 54 68318 856
rect 68486 54 68962 856
rect 69130 54 69606 856
<< metal3 >>
rect 0 99560 800 99680
rect 69200 99560 70000 99680
rect 0 99016 800 99136
rect 69200 99016 70000 99136
rect 0 98472 800 98592
rect 69200 98472 70000 98592
rect 0 97928 800 98048
rect 69200 97928 70000 98048
rect 0 97384 800 97504
rect 69200 97384 70000 97504
rect 0 96840 800 96960
rect 69200 96840 70000 96960
rect 0 96296 800 96416
rect 69200 96296 70000 96416
rect 0 95752 800 95872
rect 69200 95752 70000 95872
rect 0 95344 800 95464
rect 69200 95344 70000 95464
rect 0 94800 800 94920
rect 69200 94800 70000 94920
rect 0 94256 800 94376
rect 69200 94256 70000 94376
rect 0 93712 800 93832
rect 69200 93712 70000 93832
rect 0 93168 800 93288
rect 69200 93168 70000 93288
rect 0 92624 800 92744
rect 69200 92624 70000 92744
rect 0 92080 800 92200
rect 69200 92080 70000 92200
rect 0 91536 800 91656
rect 69200 91536 70000 91656
rect 0 90992 800 91112
rect 69200 90992 70000 91112
rect 0 90584 800 90704
rect 69200 90584 70000 90704
rect 0 90040 800 90160
rect 69200 90040 70000 90160
rect 0 89496 800 89616
rect 69200 89496 70000 89616
rect 0 88952 800 89072
rect 69200 88952 70000 89072
rect 0 88408 800 88528
rect 69200 88408 70000 88528
rect 0 87864 800 87984
rect 69200 87864 70000 87984
rect 0 87320 800 87440
rect 69200 87320 70000 87440
rect 0 86776 800 86896
rect 69200 86776 70000 86896
rect 0 86232 800 86352
rect 69200 86232 70000 86352
rect 0 85824 800 85944
rect 69200 85824 70000 85944
rect 0 85280 800 85400
rect 69200 85280 70000 85400
rect 0 84736 800 84856
rect 69200 84736 70000 84856
rect 0 84192 800 84312
rect 69200 84192 70000 84312
rect 0 83648 800 83768
rect 69200 83648 70000 83768
rect 0 83104 800 83224
rect 69200 83104 70000 83224
rect 0 82560 800 82680
rect 69200 82560 70000 82680
rect 0 82016 800 82136
rect 69200 82016 70000 82136
rect 0 81472 800 81592
rect 69200 81472 70000 81592
rect 0 81064 800 81184
rect 69200 81064 70000 81184
rect 0 80520 800 80640
rect 69200 80520 70000 80640
rect 0 79976 800 80096
rect 69200 79976 70000 80096
rect 0 79432 800 79552
rect 69200 79432 70000 79552
rect 0 78888 800 79008
rect 69200 78888 70000 79008
rect 0 78344 800 78464
rect 69200 78344 70000 78464
rect 0 77800 800 77920
rect 69200 77800 70000 77920
rect 0 77256 800 77376
rect 69200 77256 70000 77376
rect 0 76712 800 76832
rect 69200 76712 70000 76832
rect 0 76304 800 76424
rect 69200 76304 70000 76424
rect 0 75760 800 75880
rect 69200 75760 70000 75880
rect 0 75216 800 75336
rect 69200 75216 70000 75336
rect 0 74672 800 74792
rect 69200 74672 70000 74792
rect 0 74128 800 74248
rect 69200 74128 70000 74248
rect 0 73584 800 73704
rect 69200 73584 70000 73704
rect 0 73040 800 73160
rect 69200 73040 70000 73160
rect 0 72496 800 72616
rect 69200 72496 70000 72616
rect 0 71952 800 72072
rect 69200 71952 70000 72072
rect 0 71544 800 71664
rect 69200 71544 70000 71664
rect 0 71000 800 71120
rect 69200 71000 70000 71120
rect 0 70456 800 70576
rect 69200 70456 70000 70576
rect 0 69912 800 70032
rect 69200 69912 70000 70032
rect 0 69368 800 69488
rect 69200 69368 70000 69488
rect 0 68824 800 68944
rect 69200 68824 70000 68944
rect 0 68280 800 68400
rect 69200 68280 70000 68400
rect 0 67736 800 67856
rect 69200 67736 70000 67856
rect 0 67192 800 67312
rect 69200 67192 70000 67312
rect 0 66784 800 66904
rect 69200 66784 70000 66904
rect 0 66240 800 66360
rect 69200 66240 70000 66360
rect 0 65696 800 65816
rect 69200 65696 70000 65816
rect 0 65152 800 65272
rect 69200 65152 70000 65272
rect 0 64608 800 64728
rect 69200 64608 70000 64728
rect 0 64064 800 64184
rect 69200 64064 70000 64184
rect 0 63520 800 63640
rect 69200 63520 70000 63640
rect 0 62976 800 63096
rect 69200 62976 70000 63096
rect 0 62432 800 62552
rect 69200 62432 70000 62552
rect 0 62024 800 62144
rect 69200 62024 70000 62144
rect 0 61480 800 61600
rect 69200 61480 70000 61600
rect 0 60936 800 61056
rect 69200 60936 70000 61056
rect 0 60392 800 60512
rect 69200 60392 70000 60512
rect 0 59848 800 59968
rect 69200 59848 70000 59968
rect 0 59304 800 59424
rect 69200 59304 70000 59424
rect 0 58760 800 58880
rect 69200 58760 70000 58880
rect 0 58216 800 58336
rect 69200 58216 70000 58336
rect 0 57672 800 57792
rect 69200 57672 70000 57792
rect 0 57264 800 57384
rect 69200 57264 70000 57384
rect 0 56720 800 56840
rect 69200 56720 70000 56840
rect 0 56176 800 56296
rect 69200 56176 70000 56296
rect 0 55632 800 55752
rect 69200 55632 70000 55752
rect 0 55088 800 55208
rect 69200 55088 70000 55208
rect 0 54544 800 54664
rect 69200 54544 70000 54664
rect 0 54000 800 54120
rect 69200 54000 70000 54120
rect 0 53456 800 53576
rect 69200 53456 70000 53576
rect 0 52912 800 53032
rect 69200 52912 70000 53032
rect 0 52504 800 52624
rect 69200 52504 70000 52624
rect 0 51960 800 52080
rect 69200 51960 70000 52080
rect 0 51416 800 51536
rect 69200 51416 70000 51536
rect 0 50872 800 50992
rect 69200 50872 70000 50992
rect 0 50328 800 50448
rect 69200 50328 70000 50448
rect 0 49784 800 49904
rect 69200 49784 70000 49904
rect 0 49240 800 49360
rect 69200 49240 70000 49360
rect 0 48696 800 48816
rect 69200 48696 70000 48816
rect 0 48152 800 48272
rect 69200 48152 70000 48272
rect 0 47744 800 47864
rect 69200 47744 70000 47864
rect 0 47200 800 47320
rect 69200 47200 70000 47320
rect 0 46656 800 46776
rect 69200 46656 70000 46776
rect 0 46112 800 46232
rect 69200 46112 70000 46232
rect 0 45568 800 45688
rect 69200 45568 70000 45688
rect 0 45024 800 45144
rect 69200 45024 70000 45144
rect 0 44480 800 44600
rect 69200 44480 70000 44600
rect 0 43936 800 44056
rect 69200 43936 70000 44056
rect 0 43392 800 43512
rect 69200 43392 70000 43512
rect 0 42984 800 43104
rect 69200 42984 70000 43104
rect 0 42440 800 42560
rect 69200 42440 70000 42560
rect 0 41896 800 42016
rect 69200 41896 70000 42016
rect 0 41352 800 41472
rect 69200 41352 70000 41472
rect 0 40808 800 40928
rect 69200 40808 70000 40928
rect 0 40264 800 40384
rect 69200 40264 70000 40384
rect 0 39720 800 39840
rect 69200 39720 70000 39840
rect 0 39176 800 39296
rect 69200 39176 70000 39296
rect 0 38632 800 38752
rect 69200 38632 70000 38752
rect 0 38224 800 38344
rect 69200 38224 70000 38344
rect 0 37680 800 37800
rect 69200 37680 70000 37800
rect 0 37136 800 37256
rect 69200 37136 70000 37256
rect 0 36592 800 36712
rect 69200 36592 70000 36712
rect 0 36048 800 36168
rect 69200 36048 70000 36168
rect 0 35504 800 35624
rect 69200 35504 70000 35624
rect 0 34960 800 35080
rect 69200 34960 70000 35080
rect 0 34416 800 34536
rect 69200 34416 70000 34536
rect 0 33872 800 33992
rect 69200 33872 70000 33992
rect 0 33464 800 33584
rect 69200 33464 70000 33584
rect 0 32920 800 33040
rect 69200 32920 70000 33040
rect 0 32376 800 32496
rect 69200 32376 70000 32496
rect 0 31832 800 31952
rect 69200 31832 70000 31952
rect 0 31288 800 31408
rect 69200 31288 70000 31408
rect 0 30744 800 30864
rect 69200 30744 70000 30864
rect 0 30200 800 30320
rect 69200 30200 70000 30320
rect 0 29656 800 29776
rect 69200 29656 70000 29776
rect 0 29112 800 29232
rect 69200 29112 70000 29232
rect 0 28704 800 28824
rect 69200 28704 70000 28824
rect 0 28160 800 28280
rect 69200 28160 70000 28280
rect 0 27616 800 27736
rect 69200 27616 70000 27736
rect 0 27072 800 27192
rect 69200 27072 70000 27192
rect 0 26528 800 26648
rect 69200 26528 70000 26648
rect 0 25984 800 26104
rect 69200 25984 70000 26104
rect 0 25440 800 25560
rect 69200 25440 70000 25560
rect 0 24896 800 25016
rect 69200 24896 70000 25016
rect 0 24352 800 24472
rect 69200 24352 70000 24472
rect 0 23944 800 24064
rect 69200 23944 70000 24064
rect 0 23400 800 23520
rect 69200 23400 70000 23520
rect 0 22856 800 22976
rect 69200 22856 70000 22976
rect 0 22312 800 22432
rect 69200 22312 70000 22432
rect 0 21768 800 21888
rect 69200 21768 70000 21888
rect 0 21224 800 21344
rect 69200 21224 70000 21344
rect 0 20680 800 20800
rect 69200 20680 70000 20800
rect 0 20136 800 20256
rect 69200 20136 70000 20256
rect 0 19592 800 19712
rect 69200 19592 70000 19712
rect 0 19184 800 19304
rect 69200 19184 70000 19304
rect 0 18640 800 18760
rect 69200 18640 70000 18760
rect 0 18096 800 18216
rect 69200 18096 70000 18216
rect 0 17552 800 17672
rect 69200 17552 70000 17672
rect 0 17008 800 17128
rect 69200 17008 70000 17128
rect 0 16464 800 16584
rect 69200 16464 70000 16584
rect 0 15920 800 16040
rect 69200 15920 70000 16040
rect 0 15376 800 15496
rect 69200 15376 70000 15496
rect 0 14832 800 14952
rect 69200 14832 70000 14952
rect 0 14424 800 14544
rect 69200 14424 70000 14544
rect 0 13880 800 14000
rect 69200 13880 70000 14000
rect 0 13336 800 13456
rect 69200 13336 70000 13456
rect 0 12792 800 12912
rect 69200 12792 70000 12912
rect 0 12248 800 12368
rect 69200 12248 70000 12368
rect 0 11704 800 11824
rect 69200 11704 70000 11824
rect 0 11160 800 11280
rect 69200 11160 70000 11280
rect 0 10616 800 10736
rect 69200 10616 70000 10736
rect 0 10072 800 10192
rect 69200 10072 70000 10192
rect 0 9664 800 9784
rect 69200 9664 70000 9784
rect 0 9120 800 9240
rect 69200 9120 70000 9240
rect 0 8576 800 8696
rect 69200 8576 70000 8696
rect 0 8032 800 8152
rect 69200 8032 70000 8152
rect 0 7488 800 7608
rect 69200 7488 70000 7608
rect 0 6944 800 7064
rect 69200 6944 70000 7064
rect 0 6400 800 6520
rect 69200 6400 70000 6520
rect 0 5856 800 5976
rect 69200 5856 70000 5976
rect 0 5312 800 5432
rect 69200 5312 70000 5432
rect 0 4904 800 5024
rect 69200 4904 70000 5024
rect 0 4360 800 4480
rect 69200 4360 70000 4480
rect 0 3816 800 3936
rect 69200 3816 70000 3936
rect 0 3272 800 3392
rect 69200 3272 70000 3392
rect 0 2728 800 2848
rect 69200 2728 70000 2848
rect 0 2184 800 2304
rect 69200 2184 70000 2304
rect 0 1640 800 1760
rect 69200 1640 70000 1760
rect 0 1096 800 1216
rect 69200 1096 70000 1216
rect 0 552 800 672
rect 69200 552 70000 672
rect 0 144 800 264
rect 69200 144 70000 264
<< obsm3 >>
rect 880 99480 69120 99653
rect 798 99216 69200 99480
rect 880 98936 69120 99216
rect 798 98672 69200 98936
rect 880 98392 69120 98672
rect 798 98128 69200 98392
rect 880 97848 69120 98128
rect 798 97584 69200 97848
rect 880 97304 69120 97584
rect 798 97040 69200 97304
rect 880 96760 69120 97040
rect 798 96496 69200 96760
rect 880 96216 69120 96496
rect 798 95952 69200 96216
rect 880 95672 69120 95952
rect 798 95544 69200 95672
rect 880 95264 69120 95544
rect 798 95000 69200 95264
rect 880 94720 69120 95000
rect 798 94456 69200 94720
rect 880 94176 69120 94456
rect 798 93912 69200 94176
rect 880 93632 69120 93912
rect 798 93368 69200 93632
rect 880 93088 69120 93368
rect 798 92824 69200 93088
rect 880 92544 69120 92824
rect 798 92280 69200 92544
rect 880 92000 69120 92280
rect 798 91736 69200 92000
rect 880 91456 69120 91736
rect 798 91192 69200 91456
rect 880 90912 69120 91192
rect 798 90784 69200 90912
rect 880 90504 69120 90784
rect 798 90240 69200 90504
rect 880 89960 69120 90240
rect 798 89696 69200 89960
rect 880 89416 69120 89696
rect 798 89152 69200 89416
rect 880 88872 69120 89152
rect 798 88608 69200 88872
rect 880 88328 69120 88608
rect 798 88064 69200 88328
rect 880 87784 69120 88064
rect 798 87520 69200 87784
rect 880 87240 69120 87520
rect 798 86976 69200 87240
rect 880 86696 69120 86976
rect 798 86432 69200 86696
rect 880 86152 69120 86432
rect 798 86024 69200 86152
rect 880 85744 69120 86024
rect 798 85480 69200 85744
rect 880 85200 69120 85480
rect 798 84936 69200 85200
rect 880 84656 69120 84936
rect 798 84392 69200 84656
rect 880 84112 69120 84392
rect 798 83848 69200 84112
rect 880 83568 69120 83848
rect 798 83304 69200 83568
rect 880 83024 69120 83304
rect 798 82760 69200 83024
rect 880 82480 69120 82760
rect 798 82216 69200 82480
rect 880 81936 69120 82216
rect 798 81672 69200 81936
rect 880 81392 69120 81672
rect 798 81264 69200 81392
rect 880 80984 69120 81264
rect 798 80720 69200 80984
rect 880 80440 69120 80720
rect 798 80176 69200 80440
rect 880 79896 69120 80176
rect 798 79632 69200 79896
rect 880 79352 69120 79632
rect 798 79088 69200 79352
rect 880 78808 69120 79088
rect 798 78544 69200 78808
rect 880 78264 69120 78544
rect 798 78000 69200 78264
rect 880 77720 69120 78000
rect 798 77456 69200 77720
rect 880 77176 69120 77456
rect 798 76912 69200 77176
rect 880 76632 69120 76912
rect 798 76504 69200 76632
rect 880 76224 69120 76504
rect 798 75960 69200 76224
rect 880 75680 69120 75960
rect 798 75416 69200 75680
rect 880 75136 69120 75416
rect 798 74872 69200 75136
rect 880 74592 69120 74872
rect 798 74328 69200 74592
rect 880 74048 69120 74328
rect 798 73784 69200 74048
rect 880 73504 69120 73784
rect 798 73240 69200 73504
rect 880 72960 69120 73240
rect 798 72696 69200 72960
rect 880 72416 69120 72696
rect 798 72152 69200 72416
rect 880 71872 69120 72152
rect 798 71744 69200 71872
rect 880 71464 69120 71744
rect 798 71200 69200 71464
rect 880 70920 69120 71200
rect 798 70656 69200 70920
rect 880 70376 69120 70656
rect 798 70112 69200 70376
rect 880 69832 69120 70112
rect 798 69568 69200 69832
rect 880 69288 69120 69568
rect 798 69024 69200 69288
rect 880 68744 69120 69024
rect 798 68480 69200 68744
rect 880 68200 69120 68480
rect 798 67936 69200 68200
rect 880 67656 69120 67936
rect 798 67392 69200 67656
rect 880 67112 69120 67392
rect 798 66984 69200 67112
rect 880 66704 69120 66984
rect 798 66440 69200 66704
rect 880 66160 69120 66440
rect 798 65896 69200 66160
rect 880 65616 69120 65896
rect 798 65352 69200 65616
rect 880 65072 69120 65352
rect 798 64808 69200 65072
rect 880 64528 69120 64808
rect 798 64264 69200 64528
rect 880 63984 69120 64264
rect 798 63720 69200 63984
rect 880 63440 69120 63720
rect 798 63176 69200 63440
rect 880 62896 69120 63176
rect 798 62632 69200 62896
rect 880 62352 69120 62632
rect 798 62224 69200 62352
rect 880 61944 69120 62224
rect 798 61680 69200 61944
rect 880 61400 69120 61680
rect 798 61136 69200 61400
rect 880 60856 69120 61136
rect 798 60592 69200 60856
rect 880 60312 69120 60592
rect 798 60048 69200 60312
rect 880 59768 69120 60048
rect 798 59504 69200 59768
rect 880 59224 69120 59504
rect 798 58960 69200 59224
rect 880 58680 69120 58960
rect 798 58416 69200 58680
rect 880 58136 69120 58416
rect 798 57872 69200 58136
rect 880 57592 69120 57872
rect 798 57464 69200 57592
rect 880 57184 69120 57464
rect 798 56920 69200 57184
rect 880 56640 69120 56920
rect 798 56376 69200 56640
rect 880 56096 69120 56376
rect 798 55832 69200 56096
rect 880 55552 69120 55832
rect 798 55288 69200 55552
rect 880 55008 69120 55288
rect 798 54744 69200 55008
rect 880 54464 69120 54744
rect 798 54200 69200 54464
rect 880 53920 69120 54200
rect 798 53656 69200 53920
rect 880 53376 69120 53656
rect 798 53112 69200 53376
rect 880 52832 69120 53112
rect 798 52704 69200 52832
rect 880 52424 69120 52704
rect 798 52160 69200 52424
rect 880 51880 69120 52160
rect 798 51616 69200 51880
rect 880 51336 69120 51616
rect 798 51072 69200 51336
rect 880 50792 69120 51072
rect 798 50528 69200 50792
rect 880 50248 69120 50528
rect 798 49984 69200 50248
rect 880 49704 69120 49984
rect 798 49440 69200 49704
rect 880 49160 69120 49440
rect 798 48896 69200 49160
rect 880 48616 69120 48896
rect 798 48352 69200 48616
rect 880 48072 69120 48352
rect 798 47944 69200 48072
rect 880 47664 69120 47944
rect 798 47400 69200 47664
rect 880 47120 69120 47400
rect 798 46856 69200 47120
rect 880 46576 69120 46856
rect 798 46312 69200 46576
rect 880 46032 69120 46312
rect 798 45768 69200 46032
rect 880 45488 69120 45768
rect 798 45224 69200 45488
rect 880 44944 69120 45224
rect 798 44680 69200 44944
rect 880 44400 69120 44680
rect 798 44136 69200 44400
rect 880 43856 69120 44136
rect 798 43592 69200 43856
rect 880 43312 69120 43592
rect 798 43184 69200 43312
rect 880 42904 69120 43184
rect 798 42640 69200 42904
rect 880 42360 69120 42640
rect 798 42096 69200 42360
rect 880 41816 69120 42096
rect 798 41552 69200 41816
rect 880 41272 69120 41552
rect 798 41008 69200 41272
rect 880 40728 69120 41008
rect 798 40464 69200 40728
rect 880 40184 69120 40464
rect 798 39920 69200 40184
rect 880 39640 69120 39920
rect 798 39376 69200 39640
rect 880 39096 69120 39376
rect 798 38832 69200 39096
rect 880 38552 69120 38832
rect 798 38424 69200 38552
rect 880 38144 69120 38424
rect 798 37880 69200 38144
rect 880 37600 69120 37880
rect 798 37336 69200 37600
rect 880 37056 69120 37336
rect 798 36792 69200 37056
rect 880 36512 69120 36792
rect 798 36248 69200 36512
rect 880 35968 69120 36248
rect 798 35704 69200 35968
rect 880 35424 69120 35704
rect 798 35160 69200 35424
rect 880 34880 69120 35160
rect 798 34616 69200 34880
rect 880 34336 69120 34616
rect 798 34072 69200 34336
rect 880 33792 69120 34072
rect 798 33664 69200 33792
rect 880 33384 69120 33664
rect 798 33120 69200 33384
rect 880 32840 69120 33120
rect 798 32576 69200 32840
rect 880 32296 69120 32576
rect 798 32032 69200 32296
rect 880 31752 69120 32032
rect 798 31488 69200 31752
rect 880 31208 69120 31488
rect 798 30944 69200 31208
rect 880 30664 69120 30944
rect 798 30400 69200 30664
rect 880 30120 69120 30400
rect 798 29856 69200 30120
rect 880 29576 69120 29856
rect 798 29312 69200 29576
rect 880 29032 69120 29312
rect 798 28904 69200 29032
rect 880 28624 69120 28904
rect 798 28360 69200 28624
rect 880 28080 69120 28360
rect 798 27816 69200 28080
rect 880 27536 69120 27816
rect 798 27272 69200 27536
rect 880 26992 69120 27272
rect 798 26728 69200 26992
rect 880 26448 69120 26728
rect 798 26184 69200 26448
rect 880 25904 69120 26184
rect 798 25640 69200 25904
rect 880 25360 69120 25640
rect 798 25096 69200 25360
rect 880 24816 69120 25096
rect 798 24552 69200 24816
rect 880 24272 69120 24552
rect 798 24144 69200 24272
rect 880 23864 69120 24144
rect 798 23600 69200 23864
rect 880 23320 69120 23600
rect 798 23056 69200 23320
rect 880 22776 69120 23056
rect 798 22512 69200 22776
rect 880 22232 69120 22512
rect 798 21968 69200 22232
rect 880 21688 69120 21968
rect 798 21424 69200 21688
rect 880 21144 69120 21424
rect 798 20880 69200 21144
rect 880 20600 69120 20880
rect 798 20336 69200 20600
rect 880 20056 69120 20336
rect 798 19792 69200 20056
rect 880 19512 69120 19792
rect 798 19384 69200 19512
rect 880 19104 69120 19384
rect 798 18840 69200 19104
rect 880 18560 69120 18840
rect 798 18296 69200 18560
rect 880 18016 69120 18296
rect 798 17752 69200 18016
rect 880 17472 69120 17752
rect 798 17208 69200 17472
rect 880 16928 69120 17208
rect 798 16664 69200 16928
rect 880 16384 69120 16664
rect 798 16120 69200 16384
rect 880 15840 69120 16120
rect 798 15576 69200 15840
rect 880 15296 69120 15576
rect 798 15032 69200 15296
rect 880 14752 69120 15032
rect 798 14624 69200 14752
rect 880 14344 69120 14624
rect 798 14080 69200 14344
rect 880 13800 69120 14080
rect 798 13536 69200 13800
rect 880 13256 69120 13536
rect 798 12992 69200 13256
rect 880 12712 69120 12992
rect 798 12448 69200 12712
rect 880 12168 69120 12448
rect 798 11904 69200 12168
rect 880 11624 69120 11904
rect 798 11360 69200 11624
rect 880 11080 69120 11360
rect 798 10816 69200 11080
rect 880 10536 69120 10816
rect 798 10272 69200 10536
rect 880 9992 69120 10272
rect 798 9864 69200 9992
rect 880 9584 69120 9864
rect 798 9320 69200 9584
rect 880 9040 69120 9320
rect 798 8776 69200 9040
rect 880 8496 69120 8776
rect 798 8232 69200 8496
rect 880 7952 69120 8232
rect 798 7688 69200 7952
rect 880 7408 69120 7688
rect 798 7144 69200 7408
rect 880 6864 69120 7144
rect 798 6600 69200 6864
rect 880 6320 69120 6600
rect 798 6056 69200 6320
rect 880 5776 69120 6056
rect 798 5512 69200 5776
rect 880 5232 69120 5512
rect 798 5104 69200 5232
rect 880 4824 69120 5104
rect 798 4560 69200 4824
rect 880 4280 69120 4560
rect 798 4016 69200 4280
rect 880 3736 69120 4016
rect 798 3472 69200 3736
rect 880 3192 69120 3472
rect 798 2928 69200 3192
rect 880 2648 69120 2928
rect 798 2384 69200 2648
rect 880 2104 69120 2384
rect 798 1840 69200 2104
rect 880 1560 69120 1840
rect 798 1296 69200 1560
rect 880 1016 69120 1296
rect 798 752 69200 1016
rect 880 472 69120 752
rect 798 344 69200 472
rect 880 171 69120 344
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
<< obsm4 >>
rect 7971 8875 19488 84829
rect 19968 8875 34848 84829
rect 35328 8875 50208 84829
rect 50688 8875 65568 84829
rect 66048 8875 67101 84829
<< labels >>
rlabel metal3 s 0 44480 800 44600 6 sram0_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 sram0_addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 sram0_addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 sram0_addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 sram0_addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 sram0_addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 sram0_addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 sram0_addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 sram0_addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 sram0_addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 sram0_addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 sram0_addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 sram0_addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 sram0_addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 sram0_addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 sram0_addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 sram0_addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 sram0_addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 sram0_clk0
port 19 nsew signal output
rlabel metal3 s 0 144 800 264 6 sram0_clk1
port 20 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 sram0_csb0[0]
port 21 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 sram0_csb0[1]
port 22 nsew signal output
rlabel metal3 s 0 552 800 672 6 sram0_csb1[0]
port 23 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 sram0_csb1[1]
port 24 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 sram0_din0[0]
port 25 nsew signal output
rlabel metal3 s 0 54544 800 54664 6 sram0_din0[10]
port 26 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 sram0_din0[11]
port 27 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 sram0_din0[12]
port 28 nsew signal output
rlabel metal3 s 0 56176 800 56296 6 sram0_din0[13]
port 29 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 sram0_din0[14]
port 30 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 sram0_din0[15]
port 31 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 sram0_din0[16]
port 32 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 sram0_din0[17]
port 33 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 sram0_din0[18]
port 34 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 sram0_din0[19]
port 35 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 sram0_din0[1]
port 36 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 sram0_din0[20]
port 37 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 sram0_din0[21]
port 38 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 sram0_din0[22]
port 39 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 sram0_din0[23]
port 40 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 sram0_din0[24]
port 41 nsew signal output
rlabel metal3 s 0 62432 800 62552 6 sram0_din0[25]
port 42 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 sram0_din0[26]
port 43 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 sram0_din0[27]
port 44 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 sram0_din0[28]
port 45 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 sram0_din0[29]
port 46 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 sram0_din0[2]
port 47 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 sram0_din0[30]
port 48 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 sram0_din0[31]
port 49 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 sram0_din0[3]
port 50 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 sram0_din0[4]
port 51 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 sram0_din0[5]
port 52 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 sram0_din0[6]
port 53 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 sram0_din0[7]
port 54 nsew signal output
rlabel metal3 s 0 53456 800 53576 6 sram0_din0[8]
port 55 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 sram0_din0[9]
port 56 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 sram0_dout0[0]
port 57 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 sram0_dout0[10]
port 58 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 sram0_dout0[11]
port 59 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 sram0_dout0[12]
port 60 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 sram0_dout0[13]
port 61 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 sram0_dout0[14]
port 62 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 sram0_dout0[15]
port 63 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 sram0_dout0[16]
port 64 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 sram0_dout0[17]
port 65 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 sram0_dout0[18]
port 66 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 sram0_dout0[19]
port 67 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 sram0_dout0[1]
port 68 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 sram0_dout0[20]
port 69 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 sram0_dout0[21]
port 70 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 sram0_dout0[22]
port 71 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 sram0_dout0[23]
port 72 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 sram0_dout0[24]
port 73 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 sram0_dout0[25]
port 74 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 sram0_dout0[26]
port 75 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 sram0_dout0[27]
port 76 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 sram0_dout0[28]
port 77 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 sram0_dout0[29]
port 78 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 sram0_dout0[2]
port 79 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 sram0_dout0[30]
port 80 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 sram0_dout0[31]
port 81 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 sram0_dout0[32]
port 82 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 sram0_dout0[33]
port 83 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 sram0_dout0[34]
port 84 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 sram0_dout0[35]
port 85 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 sram0_dout0[36]
port 86 nsew signal input
rlabel metal3 s 0 85824 800 85944 6 sram0_dout0[37]
port 87 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 sram0_dout0[38]
port 88 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 sram0_dout0[39]
port 89 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 sram0_dout0[3]
port 90 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 sram0_dout0[40]
port 91 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 sram0_dout0[41]
port 92 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 sram0_dout0[42]
port 93 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 sram0_dout0[43]
port 94 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 sram0_dout0[44]
port 95 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 sram0_dout0[45]
port 96 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 sram0_dout0[46]
port 97 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 sram0_dout0[47]
port 98 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 sram0_dout0[48]
port 99 nsew signal input
rlabel metal3 s 0 92080 800 92200 6 sram0_dout0[49]
port 100 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 sram0_dout0[4]
port 101 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 sram0_dout0[50]
port 102 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 sram0_dout0[51]
port 103 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 sram0_dout0[52]
port 104 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 sram0_dout0[53]
port 105 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 sram0_dout0[54]
port 106 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 sram0_dout0[55]
port 107 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 sram0_dout0[56]
port 108 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 sram0_dout0[57]
port 109 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 sram0_dout0[58]
port 110 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 sram0_dout0[59]
port 111 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 sram0_dout0[5]
port 112 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 sram0_dout0[60]
port 113 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 sram0_dout0[61]
port 114 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 sram0_dout0[62]
port 115 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 sram0_dout0[63]
port 116 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 sram0_dout0[6]
port 117 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 sram0_dout0[7]
port 118 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 sram0_dout0[8]
port 119 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 sram0_dout0[9]
port 120 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 sram0_dout1[0]
port 121 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 sram0_dout1[10]
port 122 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 sram0_dout1[11]
port 123 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 sram0_dout1[12]
port 124 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 sram0_dout1[13]
port 125 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 sram0_dout1[14]
port 126 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 sram0_dout1[15]
port 127 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 sram0_dout1[16]
port 128 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 sram0_dout1[17]
port 129 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 sram0_dout1[18]
port 130 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 sram0_dout1[19]
port 131 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 sram0_dout1[1]
port 132 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 sram0_dout1[20]
port 133 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 sram0_dout1[21]
port 134 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 sram0_dout1[22]
port 135 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 sram0_dout1[23]
port 136 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 sram0_dout1[24]
port 137 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 sram0_dout1[25]
port 138 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 sram0_dout1[26]
port 139 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 sram0_dout1[27]
port 140 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 sram0_dout1[28]
port 141 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 sram0_dout1[29]
port 142 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 sram0_dout1[2]
port 143 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 sram0_dout1[30]
port 144 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 sram0_dout1[31]
port 145 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 sram0_dout1[32]
port 146 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 sram0_dout1[33]
port 147 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 sram0_dout1[34]
port 148 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 sram0_dout1[35]
port 149 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 sram0_dout1[36]
port 150 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 sram0_dout1[37]
port 151 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 sram0_dout1[38]
port 152 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 sram0_dout1[39]
port 153 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 sram0_dout1[3]
port 154 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 sram0_dout1[40]
port 155 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 sram0_dout1[41]
port 156 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 sram0_dout1[42]
port 157 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 sram0_dout1[43]
port 158 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 sram0_dout1[44]
port 159 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 sram0_dout1[45]
port 160 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 sram0_dout1[46]
port 161 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 sram0_dout1[47]
port 162 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 sram0_dout1[48]
port 163 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 sram0_dout1[49]
port 164 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 sram0_dout1[4]
port 165 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 sram0_dout1[50]
port 166 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 sram0_dout1[51]
port 167 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 sram0_dout1[52]
port 168 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 sram0_dout1[53]
port 169 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 sram0_dout1[54]
port 170 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 sram0_dout1[55]
port 171 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 sram0_dout1[56]
port 172 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 sram0_dout1[57]
port 173 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 sram0_dout1[58]
port 174 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 sram0_dout1[59]
port 175 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 sram0_dout1[5]
port 176 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 sram0_dout1[60]
port 177 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 sram0_dout1[61]
port 178 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 sram0_dout1[62]
port 179 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 sram0_dout1[63]
port 180 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 sram0_dout1[6]
port 181 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 sram0_dout1[7]
port 182 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 sram0_dout1[8]
port 183 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 sram0_dout1[9]
port 184 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 sram0_web0
port 185 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 sram0_wmask0[0]
port 186 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 sram0_wmask0[1]
port 187 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 sram0_wmask0[2]
port 188 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 sram0_wmask0[3]
port 189 nsew signal output
rlabel metal3 s 69200 44480 70000 44600 6 sram1_addr0[0]
port 190 nsew signal output
rlabel metal3 s 69200 45024 70000 45144 6 sram1_addr0[1]
port 191 nsew signal output
rlabel metal3 s 69200 45568 70000 45688 6 sram1_addr0[2]
port 192 nsew signal output
rlabel metal3 s 69200 46112 70000 46232 6 sram1_addr0[3]
port 193 nsew signal output
rlabel metal3 s 69200 46656 70000 46776 6 sram1_addr0[4]
port 194 nsew signal output
rlabel metal3 s 69200 47200 70000 47320 6 sram1_addr0[5]
port 195 nsew signal output
rlabel metal3 s 69200 47744 70000 47864 6 sram1_addr0[6]
port 196 nsew signal output
rlabel metal3 s 69200 48152 70000 48272 6 sram1_addr0[7]
port 197 nsew signal output
rlabel metal3 s 69200 48696 70000 48816 6 sram1_addr0[8]
port 198 nsew signal output
rlabel metal3 s 69200 1640 70000 1760 6 sram1_addr1[0]
port 199 nsew signal output
rlabel metal3 s 69200 2184 70000 2304 6 sram1_addr1[1]
port 200 nsew signal output
rlabel metal3 s 69200 2728 70000 2848 6 sram1_addr1[2]
port 201 nsew signal output
rlabel metal3 s 69200 3272 70000 3392 6 sram1_addr1[3]
port 202 nsew signal output
rlabel metal3 s 69200 3816 70000 3936 6 sram1_addr1[4]
port 203 nsew signal output
rlabel metal3 s 69200 4360 70000 4480 6 sram1_addr1[5]
port 204 nsew signal output
rlabel metal3 s 69200 4904 70000 5024 6 sram1_addr1[6]
port 205 nsew signal output
rlabel metal3 s 69200 5312 70000 5432 6 sram1_addr1[7]
port 206 nsew signal output
rlabel metal3 s 69200 5856 70000 5976 6 sram1_addr1[8]
port 207 nsew signal output
rlabel metal3 s 69200 40264 70000 40384 6 sram1_clk0
port 208 nsew signal output
rlabel metal3 s 69200 144 70000 264 6 sram1_clk1
port 209 nsew signal output
rlabel metal3 s 69200 40808 70000 40928 6 sram1_csb0[0]
port 210 nsew signal output
rlabel metal3 s 69200 41352 70000 41472 6 sram1_csb0[1]
port 211 nsew signal output
rlabel metal3 s 69200 552 70000 672 6 sram1_csb1[0]
port 212 nsew signal output
rlabel metal3 s 69200 1096 70000 1216 6 sram1_csb1[1]
port 213 nsew signal output
rlabel metal3 s 69200 49240 70000 49360 6 sram1_din0[0]
port 214 nsew signal output
rlabel metal3 s 69200 54544 70000 54664 6 sram1_din0[10]
port 215 nsew signal output
rlabel metal3 s 69200 55088 70000 55208 6 sram1_din0[11]
port 216 nsew signal output
rlabel metal3 s 69200 55632 70000 55752 6 sram1_din0[12]
port 217 nsew signal output
rlabel metal3 s 69200 56176 70000 56296 6 sram1_din0[13]
port 218 nsew signal output
rlabel metal3 s 69200 56720 70000 56840 6 sram1_din0[14]
port 219 nsew signal output
rlabel metal3 s 69200 57264 70000 57384 6 sram1_din0[15]
port 220 nsew signal output
rlabel metal3 s 69200 57672 70000 57792 6 sram1_din0[16]
port 221 nsew signal output
rlabel metal3 s 69200 58216 70000 58336 6 sram1_din0[17]
port 222 nsew signal output
rlabel metal3 s 69200 58760 70000 58880 6 sram1_din0[18]
port 223 nsew signal output
rlabel metal3 s 69200 59304 70000 59424 6 sram1_din0[19]
port 224 nsew signal output
rlabel metal3 s 69200 49784 70000 49904 6 sram1_din0[1]
port 225 nsew signal output
rlabel metal3 s 69200 59848 70000 59968 6 sram1_din0[20]
port 226 nsew signal output
rlabel metal3 s 69200 60392 70000 60512 6 sram1_din0[21]
port 227 nsew signal output
rlabel metal3 s 69200 60936 70000 61056 6 sram1_din0[22]
port 228 nsew signal output
rlabel metal3 s 69200 61480 70000 61600 6 sram1_din0[23]
port 229 nsew signal output
rlabel metal3 s 69200 62024 70000 62144 6 sram1_din0[24]
port 230 nsew signal output
rlabel metal3 s 69200 62432 70000 62552 6 sram1_din0[25]
port 231 nsew signal output
rlabel metal3 s 69200 62976 70000 63096 6 sram1_din0[26]
port 232 nsew signal output
rlabel metal3 s 69200 63520 70000 63640 6 sram1_din0[27]
port 233 nsew signal output
rlabel metal3 s 69200 64064 70000 64184 6 sram1_din0[28]
port 234 nsew signal output
rlabel metal3 s 69200 64608 70000 64728 6 sram1_din0[29]
port 235 nsew signal output
rlabel metal3 s 69200 50328 70000 50448 6 sram1_din0[2]
port 236 nsew signal output
rlabel metal3 s 69200 65152 70000 65272 6 sram1_din0[30]
port 237 nsew signal output
rlabel metal3 s 69200 65696 70000 65816 6 sram1_din0[31]
port 238 nsew signal output
rlabel metal3 s 69200 50872 70000 50992 6 sram1_din0[3]
port 239 nsew signal output
rlabel metal3 s 69200 51416 70000 51536 6 sram1_din0[4]
port 240 nsew signal output
rlabel metal3 s 69200 51960 70000 52080 6 sram1_din0[5]
port 241 nsew signal output
rlabel metal3 s 69200 52504 70000 52624 6 sram1_din0[6]
port 242 nsew signal output
rlabel metal3 s 69200 52912 70000 53032 6 sram1_din0[7]
port 243 nsew signal output
rlabel metal3 s 69200 53456 70000 53576 6 sram1_din0[8]
port 244 nsew signal output
rlabel metal3 s 69200 54000 70000 54120 6 sram1_din0[9]
port 245 nsew signal output
rlabel metal3 s 69200 66240 70000 66360 6 sram1_dout0[0]
port 246 nsew signal input
rlabel metal3 s 69200 71544 70000 71664 6 sram1_dout0[10]
port 247 nsew signal input
rlabel metal3 s 69200 71952 70000 72072 6 sram1_dout0[11]
port 248 nsew signal input
rlabel metal3 s 69200 72496 70000 72616 6 sram1_dout0[12]
port 249 nsew signal input
rlabel metal3 s 69200 73040 70000 73160 6 sram1_dout0[13]
port 250 nsew signal input
rlabel metal3 s 69200 73584 70000 73704 6 sram1_dout0[14]
port 251 nsew signal input
rlabel metal3 s 69200 74128 70000 74248 6 sram1_dout0[15]
port 252 nsew signal input
rlabel metal3 s 69200 74672 70000 74792 6 sram1_dout0[16]
port 253 nsew signal input
rlabel metal3 s 69200 75216 70000 75336 6 sram1_dout0[17]
port 254 nsew signal input
rlabel metal3 s 69200 75760 70000 75880 6 sram1_dout0[18]
port 255 nsew signal input
rlabel metal3 s 69200 76304 70000 76424 6 sram1_dout0[19]
port 256 nsew signal input
rlabel metal3 s 69200 66784 70000 66904 6 sram1_dout0[1]
port 257 nsew signal input
rlabel metal3 s 69200 76712 70000 76832 6 sram1_dout0[20]
port 258 nsew signal input
rlabel metal3 s 69200 77256 70000 77376 6 sram1_dout0[21]
port 259 nsew signal input
rlabel metal3 s 69200 77800 70000 77920 6 sram1_dout0[22]
port 260 nsew signal input
rlabel metal3 s 69200 78344 70000 78464 6 sram1_dout0[23]
port 261 nsew signal input
rlabel metal3 s 69200 78888 70000 79008 6 sram1_dout0[24]
port 262 nsew signal input
rlabel metal3 s 69200 79432 70000 79552 6 sram1_dout0[25]
port 263 nsew signal input
rlabel metal3 s 69200 79976 70000 80096 6 sram1_dout0[26]
port 264 nsew signal input
rlabel metal3 s 69200 80520 70000 80640 6 sram1_dout0[27]
port 265 nsew signal input
rlabel metal3 s 69200 81064 70000 81184 6 sram1_dout0[28]
port 266 nsew signal input
rlabel metal3 s 69200 81472 70000 81592 6 sram1_dout0[29]
port 267 nsew signal input
rlabel metal3 s 69200 67192 70000 67312 6 sram1_dout0[2]
port 268 nsew signal input
rlabel metal3 s 69200 82016 70000 82136 6 sram1_dout0[30]
port 269 nsew signal input
rlabel metal3 s 69200 82560 70000 82680 6 sram1_dout0[31]
port 270 nsew signal input
rlabel metal3 s 69200 83104 70000 83224 6 sram1_dout0[32]
port 271 nsew signal input
rlabel metal3 s 69200 83648 70000 83768 6 sram1_dout0[33]
port 272 nsew signal input
rlabel metal3 s 69200 84192 70000 84312 6 sram1_dout0[34]
port 273 nsew signal input
rlabel metal3 s 69200 84736 70000 84856 6 sram1_dout0[35]
port 274 nsew signal input
rlabel metal3 s 69200 85280 70000 85400 6 sram1_dout0[36]
port 275 nsew signal input
rlabel metal3 s 69200 85824 70000 85944 6 sram1_dout0[37]
port 276 nsew signal input
rlabel metal3 s 69200 86232 70000 86352 6 sram1_dout0[38]
port 277 nsew signal input
rlabel metal3 s 69200 86776 70000 86896 6 sram1_dout0[39]
port 278 nsew signal input
rlabel metal3 s 69200 67736 70000 67856 6 sram1_dout0[3]
port 279 nsew signal input
rlabel metal3 s 69200 87320 70000 87440 6 sram1_dout0[40]
port 280 nsew signal input
rlabel metal3 s 69200 87864 70000 87984 6 sram1_dout0[41]
port 281 nsew signal input
rlabel metal3 s 69200 88408 70000 88528 6 sram1_dout0[42]
port 282 nsew signal input
rlabel metal3 s 69200 88952 70000 89072 6 sram1_dout0[43]
port 283 nsew signal input
rlabel metal3 s 69200 89496 70000 89616 6 sram1_dout0[44]
port 284 nsew signal input
rlabel metal3 s 69200 90040 70000 90160 6 sram1_dout0[45]
port 285 nsew signal input
rlabel metal3 s 69200 90584 70000 90704 6 sram1_dout0[46]
port 286 nsew signal input
rlabel metal3 s 69200 90992 70000 91112 6 sram1_dout0[47]
port 287 nsew signal input
rlabel metal3 s 69200 91536 70000 91656 6 sram1_dout0[48]
port 288 nsew signal input
rlabel metal3 s 69200 92080 70000 92200 6 sram1_dout0[49]
port 289 nsew signal input
rlabel metal3 s 69200 68280 70000 68400 6 sram1_dout0[4]
port 290 nsew signal input
rlabel metal3 s 69200 92624 70000 92744 6 sram1_dout0[50]
port 291 nsew signal input
rlabel metal3 s 69200 93168 70000 93288 6 sram1_dout0[51]
port 292 nsew signal input
rlabel metal3 s 69200 93712 70000 93832 6 sram1_dout0[52]
port 293 nsew signal input
rlabel metal3 s 69200 94256 70000 94376 6 sram1_dout0[53]
port 294 nsew signal input
rlabel metal3 s 69200 94800 70000 94920 6 sram1_dout0[54]
port 295 nsew signal input
rlabel metal3 s 69200 95344 70000 95464 6 sram1_dout0[55]
port 296 nsew signal input
rlabel metal3 s 69200 95752 70000 95872 6 sram1_dout0[56]
port 297 nsew signal input
rlabel metal3 s 69200 96296 70000 96416 6 sram1_dout0[57]
port 298 nsew signal input
rlabel metal3 s 69200 96840 70000 96960 6 sram1_dout0[58]
port 299 nsew signal input
rlabel metal3 s 69200 97384 70000 97504 6 sram1_dout0[59]
port 300 nsew signal input
rlabel metal3 s 69200 68824 70000 68944 6 sram1_dout0[5]
port 301 nsew signal input
rlabel metal3 s 69200 97928 70000 98048 6 sram1_dout0[60]
port 302 nsew signal input
rlabel metal3 s 69200 98472 70000 98592 6 sram1_dout0[61]
port 303 nsew signal input
rlabel metal3 s 69200 99016 70000 99136 6 sram1_dout0[62]
port 304 nsew signal input
rlabel metal3 s 69200 99560 70000 99680 6 sram1_dout0[63]
port 305 nsew signal input
rlabel metal3 s 69200 69368 70000 69488 6 sram1_dout0[6]
port 306 nsew signal input
rlabel metal3 s 69200 69912 70000 70032 6 sram1_dout0[7]
port 307 nsew signal input
rlabel metal3 s 69200 70456 70000 70576 6 sram1_dout0[8]
port 308 nsew signal input
rlabel metal3 s 69200 71000 70000 71120 6 sram1_dout0[9]
port 309 nsew signal input
rlabel metal3 s 69200 6400 70000 6520 6 sram1_dout1[0]
port 310 nsew signal input
rlabel metal3 s 69200 11704 70000 11824 6 sram1_dout1[10]
port 311 nsew signal input
rlabel metal3 s 69200 12248 70000 12368 6 sram1_dout1[11]
port 312 nsew signal input
rlabel metal3 s 69200 12792 70000 12912 6 sram1_dout1[12]
port 313 nsew signal input
rlabel metal3 s 69200 13336 70000 13456 6 sram1_dout1[13]
port 314 nsew signal input
rlabel metal3 s 69200 13880 70000 14000 6 sram1_dout1[14]
port 315 nsew signal input
rlabel metal3 s 69200 14424 70000 14544 6 sram1_dout1[15]
port 316 nsew signal input
rlabel metal3 s 69200 14832 70000 14952 6 sram1_dout1[16]
port 317 nsew signal input
rlabel metal3 s 69200 15376 70000 15496 6 sram1_dout1[17]
port 318 nsew signal input
rlabel metal3 s 69200 15920 70000 16040 6 sram1_dout1[18]
port 319 nsew signal input
rlabel metal3 s 69200 16464 70000 16584 6 sram1_dout1[19]
port 320 nsew signal input
rlabel metal3 s 69200 6944 70000 7064 6 sram1_dout1[1]
port 321 nsew signal input
rlabel metal3 s 69200 17008 70000 17128 6 sram1_dout1[20]
port 322 nsew signal input
rlabel metal3 s 69200 17552 70000 17672 6 sram1_dout1[21]
port 323 nsew signal input
rlabel metal3 s 69200 18096 70000 18216 6 sram1_dout1[22]
port 324 nsew signal input
rlabel metal3 s 69200 18640 70000 18760 6 sram1_dout1[23]
port 325 nsew signal input
rlabel metal3 s 69200 19184 70000 19304 6 sram1_dout1[24]
port 326 nsew signal input
rlabel metal3 s 69200 19592 70000 19712 6 sram1_dout1[25]
port 327 nsew signal input
rlabel metal3 s 69200 20136 70000 20256 6 sram1_dout1[26]
port 328 nsew signal input
rlabel metal3 s 69200 20680 70000 20800 6 sram1_dout1[27]
port 329 nsew signal input
rlabel metal3 s 69200 21224 70000 21344 6 sram1_dout1[28]
port 330 nsew signal input
rlabel metal3 s 69200 21768 70000 21888 6 sram1_dout1[29]
port 331 nsew signal input
rlabel metal3 s 69200 7488 70000 7608 6 sram1_dout1[2]
port 332 nsew signal input
rlabel metal3 s 69200 22312 70000 22432 6 sram1_dout1[30]
port 333 nsew signal input
rlabel metal3 s 69200 22856 70000 22976 6 sram1_dout1[31]
port 334 nsew signal input
rlabel metal3 s 69200 23400 70000 23520 6 sram1_dout1[32]
port 335 nsew signal input
rlabel metal3 s 69200 23944 70000 24064 6 sram1_dout1[33]
port 336 nsew signal input
rlabel metal3 s 69200 24352 70000 24472 6 sram1_dout1[34]
port 337 nsew signal input
rlabel metal3 s 69200 24896 70000 25016 6 sram1_dout1[35]
port 338 nsew signal input
rlabel metal3 s 69200 25440 70000 25560 6 sram1_dout1[36]
port 339 nsew signal input
rlabel metal3 s 69200 25984 70000 26104 6 sram1_dout1[37]
port 340 nsew signal input
rlabel metal3 s 69200 26528 70000 26648 6 sram1_dout1[38]
port 341 nsew signal input
rlabel metal3 s 69200 27072 70000 27192 6 sram1_dout1[39]
port 342 nsew signal input
rlabel metal3 s 69200 8032 70000 8152 6 sram1_dout1[3]
port 343 nsew signal input
rlabel metal3 s 69200 27616 70000 27736 6 sram1_dout1[40]
port 344 nsew signal input
rlabel metal3 s 69200 28160 70000 28280 6 sram1_dout1[41]
port 345 nsew signal input
rlabel metal3 s 69200 28704 70000 28824 6 sram1_dout1[42]
port 346 nsew signal input
rlabel metal3 s 69200 29112 70000 29232 6 sram1_dout1[43]
port 347 nsew signal input
rlabel metal3 s 69200 29656 70000 29776 6 sram1_dout1[44]
port 348 nsew signal input
rlabel metal3 s 69200 30200 70000 30320 6 sram1_dout1[45]
port 349 nsew signal input
rlabel metal3 s 69200 30744 70000 30864 6 sram1_dout1[46]
port 350 nsew signal input
rlabel metal3 s 69200 31288 70000 31408 6 sram1_dout1[47]
port 351 nsew signal input
rlabel metal3 s 69200 31832 70000 31952 6 sram1_dout1[48]
port 352 nsew signal input
rlabel metal3 s 69200 32376 70000 32496 6 sram1_dout1[49]
port 353 nsew signal input
rlabel metal3 s 69200 8576 70000 8696 6 sram1_dout1[4]
port 354 nsew signal input
rlabel metal3 s 69200 32920 70000 33040 6 sram1_dout1[50]
port 355 nsew signal input
rlabel metal3 s 69200 33464 70000 33584 6 sram1_dout1[51]
port 356 nsew signal input
rlabel metal3 s 69200 33872 70000 33992 6 sram1_dout1[52]
port 357 nsew signal input
rlabel metal3 s 69200 34416 70000 34536 6 sram1_dout1[53]
port 358 nsew signal input
rlabel metal3 s 69200 34960 70000 35080 6 sram1_dout1[54]
port 359 nsew signal input
rlabel metal3 s 69200 35504 70000 35624 6 sram1_dout1[55]
port 360 nsew signal input
rlabel metal3 s 69200 36048 70000 36168 6 sram1_dout1[56]
port 361 nsew signal input
rlabel metal3 s 69200 36592 70000 36712 6 sram1_dout1[57]
port 362 nsew signal input
rlabel metal3 s 69200 37136 70000 37256 6 sram1_dout1[58]
port 363 nsew signal input
rlabel metal3 s 69200 37680 70000 37800 6 sram1_dout1[59]
port 364 nsew signal input
rlabel metal3 s 69200 9120 70000 9240 6 sram1_dout1[5]
port 365 nsew signal input
rlabel metal3 s 69200 38224 70000 38344 6 sram1_dout1[60]
port 366 nsew signal input
rlabel metal3 s 69200 38632 70000 38752 6 sram1_dout1[61]
port 367 nsew signal input
rlabel metal3 s 69200 39176 70000 39296 6 sram1_dout1[62]
port 368 nsew signal input
rlabel metal3 s 69200 39720 70000 39840 6 sram1_dout1[63]
port 369 nsew signal input
rlabel metal3 s 69200 9664 70000 9784 6 sram1_dout1[6]
port 370 nsew signal input
rlabel metal3 s 69200 10072 70000 10192 6 sram1_dout1[7]
port 371 nsew signal input
rlabel metal3 s 69200 10616 70000 10736 6 sram1_dout1[8]
port 372 nsew signal input
rlabel metal3 s 69200 11160 70000 11280 6 sram1_dout1[9]
port 373 nsew signal input
rlabel metal3 s 69200 41896 70000 42016 6 sram1_web0
port 374 nsew signal output
rlabel metal3 s 69200 42440 70000 42560 6 sram1_wmask0[0]
port 375 nsew signal output
rlabel metal3 s 69200 42984 70000 43104 6 sram1_wmask0[1]
port 376 nsew signal output
rlabel metal3 s 69200 43392 70000 43512 6 sram1_wmask0[2]
port 377 nsew signal output
rlabel metal3 s 69200 43936 70000 44056 6 sram1_wmask0[3]
port 378 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 379 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 379 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 379 nsew power input
rlabel metal2 s 66442 0 66498 800 6 vga_b[0]
port 380 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 vga_b[1]
port 381 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 vga_g[0]
port 382 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 vga_g[1]
port 383 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 vga_hsync
port 384 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 vga_r[0]
port 385 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 vga_r[1]
port 386 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 vga_vsync
port 387 nsew signal output
rlabel metal2 s 294 0 350 800 6 video_irq[0]
port 388 nsew signal output
rlabel metal2 s 846 0 902 800 6 video_irq[1]
port 389 nsew signal output
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 390 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 390 nsew ground input
rlabel metal2 s 1490 0 1546 800 6 wb_ack_o
port 391 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wb_adr_i[0]
port 392 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wb_adr_i[10]
port 393 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wb_adr_i[11]
port 394 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wb_adr_i[12]
port 395 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wb_adr_i[13]
port 396 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wb_adr_i[14]
port 397 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wb_adr_i[15]
port 398 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wb_adr_i[16]
port 399 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wb_adr_i[17]
port 400 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wb_adr_i[18]
port 401 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wb_adr_i[19]
port 402 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wb_adr_i[1]
port 403 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wb_adr_i[20]
port 404 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wb_adr_i[21]
port 405 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wb_adr_i[22]
port 406 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wb_adr_i[23]
port 407 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wb_adr_i[2]
port 408 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wb_adr_i[3]
port 409 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wb_adr_i[4]
port 410 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wb_adr_i[5]
port 411 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wb_adr_i[6]
port 412 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wb_adr_i[7]
port 413 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb_adr_i[8]
port 414 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wb_adr_i[9]
port 415 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wb_clk_i
port 416 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wb_cyc_i
port 417 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_data_i[0]
port 418 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wb_data_i[10]
port 419 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wb_data_i[11]
port 420 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wb_data_i[12]
port 421 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wb_data_i[13]
port 422 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wb_data_i[14]
port 423 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wb_data_i[15]
port 424 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wb_data_i[16]
port 425 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wb_data_i[17]
port 426 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wb_data_i[18]
port 427 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wb_data_i[19]
port 428 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wb_data_i[1]
port 429 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wb_data_i[20]
port 430 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wb_data_i[21]
port 431 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wb_data_i[22]
port 432 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wb_data_i[23]
port 433 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wb_data_i[24]
port 434 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wb_data_i[25]
port 435 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wb_data_i[26]
port 436 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 wb_data_i[27]
port 437 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wb_data_i[28]
port 438 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 wb_data_i[29]
port 439 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wb_data_i[2]
port 440 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wb_data_i[30]
port 441 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 wb_data_i[31]
port 442 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wb_data_i[3]
port 443 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wb_data_i[4]
port 444 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wb_data_i[5]
port 445 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wb_data_i[6]
port 446 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wb_data_i[7]
port 447 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wb_data_i[8]
port 448 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wb_data_i[9]
port 449 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wb_data_o[0]
port 450 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wb_data_o[10]
port 451 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wb_data_o[11]
port 452 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wb_data_o[12]
port 453 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wb_data_o[13]
port 454 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 wb_data_o[14]
port 455 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wb_data_o[15]
port 456 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wb_data_o[16]
port 457 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wb_data_o[17]
port 458 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wb_data_o[18]
port 459 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 wb_data_o[19]
port 460 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wb_data_o[1]
port 461 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wb_data_o[20]
port 462 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wb_data_o[21]
port 463 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 wb_data_o[22]
port 464 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 wb_data_o[23]
port 465 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wb_data_o[24]
port 466 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wb_data_o[25]
port 467 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 wb_data_o[26]
port 468 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 wb_data_o[27]
port 469 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 wb_data_o[28]
port 470 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 wb_data_o[29]
port 471 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wb_data_o[2]
port 472 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 wb_data_o[30]
port 473 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 wb_data_o[31]
port 474 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wb_data_o[3]
port 475 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wb_data_o[4]
port 476 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wb_data_o[5]
port 477 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wb_data_o[6]
port 478 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wb_data_o[7]
port 479 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wb_data_o[8]
port 480 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wb_data_o[9]
port 481 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 wb_error_o
port 482 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wb_rst_i
port 483 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wb_sel_i[0]
port 484 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wb_sel_i[1]
port 485 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wb_sel_i[2]
port 486 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wb_sel_i[3]
port 487 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wb_stall_o
port 488 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wb_stb_i
port 489 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb_we_i
port 490 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9073506
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Video/runs/Video/results/finishing/Video.magic.gds
string GDS_START 892618
<< end >>

