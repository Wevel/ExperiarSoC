magic
tech sky130A
magscale 1 2
timestamp 1654557611
<< obsli1 >>
rect 1104 2159 58880 39729
<< obsm1 >>
rect 198 1028 59694 39760
<< metal2 >>
rect 3698 41200 3754 42000
rect 11150 41200 11206 42000
rect 18694 41200 18750 42000
rect 26146 41200 26202 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48686 41200 48742 42000
rect 56138 41200 56194 42000
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
<< obsm2 >>
rect 204 41144 3642 41721
rect 3810 41144 11094 41721
rect 11262 41144 18638 41721
rect 18806 41144 26090 41721
rect 26258 41144 33634 41721
rect 33802 41144 41086 41721
rect 41254 41144 48630 41721
rect 48798 41144 56082 41721
rect 56250 41144 59688 41721
rect 204 856 59688 41144
rect 314 167 606 856
rect 774 167 1066 856
rect 1234 167 1526 856
rect 1694 167 2078 856
rect 2246 167 2538 856
rect 2706 167 2998 856
rect 3166 167 3550 856
rect 3718 167 4010 856
rect 4178 167 4470 856
rect 4638 167 5022 856
rect 5190 167 5482 856
rect 5650 167 5942 856
rect 6110 167 6402 856
rect 6570 167 6954 856
rect 7122 167 7414 856
rect 7582 167 7874 856
rect 8042 167 8426 856
rect 8594 167 8886 856
rect 9054 167 9346 856
rect 9514 167 9898 856
rect 10066 167 10358 856
rect 10526 167 10818 856
rect 10986 167 11278 856
rect 11446 167 11830 856
rect 11998 167 12290 856
rect 12458 167 12750 856
rect 12918 167 13302 856
rect 13470 167 13762 856
rect 13930 167 14222 856
rect 14390 167 14774 856
rect 14942 167 15234 856
rect 15402 167 15694 856
rect 15862 167 16154 856
rect 16322 167 16706 856
rect 16874 167 17166 856
rect 17334 167 17626 856
rect 17794 167 18178 856
rect 18346 167 18638 856
rect 18806 167 19098 856
rect 19266 167 19650 856
rect 19818 167 20110 856
rect 20278 167 20570 856
rect 20738 167 21030 856
rect 21198 167 21582 856
rect 21750 167 22042 856
rect 22210 167 22502 856
rect 22670 167 23054 856
rect 23222 167 23514 856
rect 23682 167 23974 856
rect 24142 167 24526 856
rect 24694 167 24986 856
rect 25154 167 25446 856
rect 25614 167 25906 856
rect 26074 167 26458 856
rect 26626 167 26918 856
rect 27086 167 27378 856
rect 27546 167 27930 856
rect 28098 167 28390 856
rect 28558 167 28850 856
rect 29018 167 29402 856
rect 29570 167 29862 856
rect 30030 167 30322 856
rect 30490 167 30782 856
rect 30950 167 31334 856
rect 31502 167 31794 856
rect 31962 167 32254 856
rect 32422 167 32806 856
rect 32974 167 33266 856
rect 33434 167 33726 856
rect 33894 167 34278 856
rect 34446 167 34738 856
rect 34906 167 35198 856
rect 35366 167 35658 856
rect 35826 167 36210 856
rect 36378 167 36670 856
rect 36838 167 37130 856
rect 37298 167 37682 856
rect 37850 167 38142 856
rect 38310 167 38602 856
rect 38770 167 39154 856
rect 39322 167 39614 856
rect 39782 167 40074 856
rect 40242 167 40534 856
rect 40702 167 41086 856
rect 41254 167 41546 856
rect 41714 167 42006 856
rect 42174 167 42558 856
rect 42726 167 43018 856
rect 43186 167 43478 856
rect 43646 167 44030 856
rect 44198 167 44490 856
rect 44658 167 44950 856
rect 45118 167 45410 856
rect 45578 167 45962 856
rect 46130 167 46422 856
rect 46590 167 46882 856
rect 47050 167 47434 856
rect 47602 167 47894 856
rect 48062 167 48354 856
rect 48522 167 48906 856
rect 49074 167 49366 856
rect 49534 167 49826 856
rect 49994 167 50286 856
rect 50454 167 50838 856
rect 51006 167 51298 856
rect 51466 167 51758 856
rect 51926 167 52310 856
rect 52478 167 52770 856
rect 52938 167 53230 856
rect 53398 167 53782 856
rect 53950 167 54242 856
rect 54410 167 54702 856
rect 54870 167 55162 856
rect 55330 167 55714 856
rect 55882 167 56174 856
rect 56342 167 56634 856
rect 56802 167 57186 856
rect 57354 167 57646 856
rect 57814 167 58106 856
rect 58274 167 58658 856
rect 58826 167 59118 856
rect 59286 167 59578 856
<< metal3 >>
rect 0 41624 800 41744
rect 0 41216 800 41336
rect 0 40808 800 40928
rect 0 40400 800 40520
rect 0 39992 800 40112
rect 0 39584 800 39704
rect 0 39176 800 39296
rect 0 38768 800 38888
rect 0 38360 800 38480
rect 0 37952 800 38072
rect 0 37544 800 37664
rect 0 37000 800 37120
rect 0 36592 800 36712
rect 0 36184 800 36304
rect 0 35776 800 35896
rect 0 35368 800 35488
rect 0 34960 800 35080
rect 0 34552 800 34672
rect 0 34144 800 34264
rect 0 33736 800 33856
rect 0 33328 800 33448
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 0 31968 800 32088
rect 0 31560 800 31680
rect 0 31152 800 31272
rect 0 30744 800 30864
rect 0 30336 800 30456
rect 0 29928 800 30048
rect 0 29520 800 29640
rect 0 29112 800 29232
rect 0 28704 800 28824
rect 0 28296 800 28416
rect 0 27752 800 27872
rect 0 27344 800 27464
rect 0 26936 800 27056
rect 0 26528 800 26648
rect 0 26120 800 26240
rect 0 25712 800 25832
rect 0 25304 800 25424
rect 0 24896 800 25016
rect 0 24488 800 24608
rect 0 24080 800 24200
rect 0 23672 800 23792
rect 0 23128 800 23248
rect 0 22720 800 22840
rect 0 22312 800 22432
rect 0 21904 800 22024
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 0 20680 800 20800
rect 0 20272 800 20392
rect 0 19864 800 19984
rect 0 19456 800 19576
rect 0 19048 800 19168
rect 0 18504 800 18624
rect 0 18096 800 18216
rect 0 17688 800 17808
rect 0 17280 800 17400
rect 0 16872 800 16992
rect 0 16464 800 16584
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 0 15240 800 15360
rect 0 14832 800 14952
rect 0 14424 800 14544
rect 0 13880 800 14000
rect 0 13472 800 13592
rect 0 13064 800 13184
rect 0 12656 800 12776
rect 0 12248 800 12368
rect 0 11840 800 11960
rect 0 11432 800 11552
rect 0 11024 800 11144
rect 0 10616 800 10736
rect 0 10208 800 10328
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 0 8848 800 8968
rect 0 8440 800 8560
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6808 800 6928
rect 0 6400 800 6520
rect 0 5992 800 6112
rect 0 5584 800 5704
rect 0 5176 800 5296
rect 0 4632 800 4752
rect 0 4224 800 4344
rect 0 3816 800 3936
rect 0 3408 800 3528
rect 0 3000 800 3120
rect 0 2592 800 2712
rect 0 2184 800 2304
rect 0 1776 800 1896
rect 0 1368 800 1488
rect 0 960 800 1080
rect 0 552 800 672
rect 0 144 800 264
<< obsm3 >>
rect 880 41544 55923 41717
rect 800 41416 55923 41544
rect 880 41136 55923 41416
rect 800 41008 55923 41136
rect 880 40728 55923 41008
rect 800 40600 55923 40728
rect 880 40320 55923 40600
rect 800 40192 55923 40320
rect 880 39912 55923 40192
rect 800 39784 55923 39912
rect 880 39504 55923 39784
rect 800 39376 55923 39504
rect 880 39096 55923 39376
rect 800 38968 55923 39096
rect 880 38688 55923 38968
rect 800 38560 55923 38688
rect 880 38280 55923 38560
rect 800 38152 55923 38280
rect 880 37872 55923 38152
rect 800 37744 55923 37872
rect 880 37464 55923 37744
rect 800 37200 55923 37464
rect 880 36920 55923 37200
rect 800 36792 55923 36920
rect 880 36512 55923 36792
rect 800 36384 55923 36512
rect 880 36104 55923 36384
rect 800 35976 55923 36104
rect 880 35696 55923 35976
rect 800 35568 55923 35696
rect 880 35288 55923 35568
rect 800 35160 55923 35288
rect 880 34880 55923 35160
rect 800 34752 55923 34880
rect 880 34472 55923 34752
rect 800 34344 55923 34472
rect 880 34064 55923 34344
rect 800 33936 55923 34064
rect 880 33656 55923 33936
rect 800 33528 55923 33656
rect 880 33248 55923 33528
rect 800 33120 55923 33248
rect 880 32840 55923 33120
rect 800 32576 55923 32840
rect 880 32296 55923 32576
rect 800 32168 55923 32296
rect 880 31888 55923 32168
rect 800 31760 55923 31888
rect 880 31480 55923 31760
rect 800 31352 55923 31480
rect 880 31072 55923 31352
rect 800 30944 55923 31072
rect 880 30664 55923 30944
rect 800 30536 55923 30664
rect 880 30256 55923 30536
rect 800 30128 55923 30256
rect 880 29848 55923 30128
rect 800 29720 55923 29848
rect 880 29440 55923 29720
rect 800 29312 55923 29440
rect 880 29032 55923 29312
rect 800 28904 55923 29032
rect 880 28624 55923 28904
rect 800 28496 55923 28624
rect 880 28216 55923 28496
rect 800 27952 55923 28216
rect 880 27672 55923 27952
rect 800 27544 55923 27672
rect 880 27264 55923 27544
rect 800 27136 55923 27264
rect 880 26856 55923 27136
rect 800 26728 55923 26856
rect 880 26448 55923 26728
rect 800 26320 55923 26448
rect 880 26040 55923 26320
rect 800 25912 55923 26040
rect 880 25632 55923 25912
rect 800 25504 55923 25632
rect 880 25224 55923 25504
rect 800 25096 55923 25224
rect 880 24816 55923 25096
rect 800 24688 55923 24816
rect 880 24408 55923 24688
rect 800 24280 55923 24408
rect 880 24000 55923 24280
rect 800 23872 55923 24000
rect 880 23592 55923 23872
rect 800 23328 55923 23592
rect 880 23048 55923 23328
rect 800 22920 55923 23048
rect 880 22640 55923 22920
rect 800 22512 55923 22640
rect 880 22232 55923 22512
rect 800 22104 55923 22232
rect 880 21824 55923 22104
rect 800 21696 55923 21824
rect 880 21416 55923 21696
rect 800 21288 55923 21416
rect 880 21008 55923 21288
rect 800 20880 55923 21008
rect 880 20600 55923 20880
rect 800 20472 55923 20600
rect 880 20192 55923 20472
rect 800 20064 55923 20192
rect 880 19784 55923 20064
rect 800 19656 55923 19784
rect 880 19376 55923 19656
rect 800 19248 55923 19376
rect 880 18968 55923 19248
rect 800 18704 55923 18968
rect 880 18424 55923 18704
rect 800 18296 55923 18424
rect 880 18016 55923 18296
rect 800 17888 55923 18016
rect 880 17608 55923 17888
rect 800 17480 55923 17608
rect 880 17200 55923 17480
rect 800 17072 55923 17200
rect 880 16792 55923 17072
rect 800 16664 55923 16792
rect 880 16384 55923 16664
rect 800 16256 55923 16384
rect 880 15976 55923 16256
rect 800 15848 55923 15976
rect 880 15568 55923 15848
rect 800 15440 55923 15568
rect 880 15160 55923 15440
rect 800 15032 55923 15160
rect 880 14752 55923 15032
rect 800 14624 55923 14752
rect 880 14344 55923 14624
rect 800 14080 55923 14344
rect 880 13800 55923 14080
rect 800 13672 55923 13800
rect 880 13392 55923 13672
rect 800 13264 55923 13392
rect 880 12984 55923 13264
rect 800 12856 55923 12984
rect 880 12576 55923 12856
rect 800 12448 55923 12576
rect 880 12168 55923 12448
rect 800 12040 55923 12168
rect 880 11760 55923 12040
rect 800 11632 55923 11760
rect 880 11352 55923 11632
rect 800 11224 55923 11352
rect 880 10944 55923 11224
rect 800 10816 55923 10944
rect 880 10536 55923 10816
rect 800 10408 55923 10536
rect 880 10128 55923 10408
rect 800 10000 55923 10128
rect 880 9720 55923 10000
rect 800 9456 55923 9720
rect 880 9176 55923 9456
rect 800 9048 55923 9176
rect 880 8768 55923 9048
rect 800 8640 55923 8768
rect 880 8360 55923 8640
rect 800 8232 55923 8360
rect 880 7952 55923 8232
rect 800 7824 55923 7952
rect 880 7544 55923 7824
rect 800 7416 55923 7544
rect 880 7136 55923 7416
rect 800 7008 55923 7136
rect 880 6728 55923 7008
rect 800 6600 55923 6728
rect 880 6320 55923 6600
rect 800 6192 55923 6320
rect 880 5912 55923 6192
rect 800 5784 55923 5912
rect 880 5504 55923 5784
rect 800 5376 55923 5504
rect 880 5096 55923 5376
rect 800 4832 55923 5096
rect 880 4552 55923 4832
rect 800 4424 55923 4552
rect 880 4144 55923 4424
rect 800 4016 55923 4144
rect 880 3736 55923 4016
rect 800 3608 55923 3736
rect 880 3328 55923 3608
rect 800 3200 55923 3328
rect 880 2920 55923 3200
rect 800 2792 55923 2920
rect 880 2512 55923 2792
rect 800 2384 55923 2512
rect 880 2104 55923 2384
rect 800 1976 55923 2104
rect 880 1696 55923 1976
rect 800 1568 55923 1696
rect 880 1288 55923 1568
rect 800 1160 55923 1288
rect 880 880 55923 1160
rect 800 752 55923 880
rect 880 472 55923 752
rect 800 344 55923 472
rect 880 171 55923 344
<< metal4 >>
rect 4208 2128 4528 39760
rect 19568 2128 19888 39760
rect 34928 2128 35248 39760
rect 50288 2128 50608 39760
<< obsm4 >>
rect 9811 2347 10613 23493
<< labels >>
rlabel metal2 s 3698 41200 3754 42000 6 flash_csb
port 1 nsew signal output
rlabel metal2 s 11150 41200 11206 42000 6 flash_io0_read
port 2 nsew signal input
rlabel metal2 s 18694 41200 18750 42000 6 flash_io0_we
port 3 nsew signal output
rlabel metal2 s 26146 41200 26202 42000 6 flash_io0_write
port 4 nsew signal output
rlabel metal2 s 33690 41200 33746 42000 6 flash_io1_read
port 5 nsew signal input
rlabel metal2 s 41142 41200 41198 42000 6 flash_io1_we
port 6 nsew signal output
rlabel metal2 s 48686 41200 48742 42000 6 flash_io1_write
port 7 nsew signal output
rlabel metal2 s 56138 41200 56194 42000 6 flash_sck
port 8 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 sram_addr0[0]
port 9 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 sram_addr0[1]
port 10 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 sram_addr0[2]
port 11 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 sram_addr0[3]
port 12 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[4]
port 13 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 sram_addr0[5]
port 14 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 sram_addr0[6]
port 15 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 sram_addr0[7]
port 16 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 sram_addr0[8]
port 17 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 sram_addr1[0]
port 18 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 sram_addr1[1]
port 19 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 sram_addr1[2]
port 20 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 sram_addr1[3]
port 21 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 sram_addr1[4]
port 22 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 sram_addr1[5]
port 23 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 sram_addr1[6]
port 24 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 sram_addr1[7]
port 25 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 sram_addr1[8]
port 26 nsew signal output
rlabel metal2 s 202 0 258 800 6 sram_clk0
port 27 nsew signal output
rlabel metal2 s 662 0 718 800 6 sram_clk1
port 28 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 sram_csb0
port 29 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 sram_csb1
port 30 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 sram_din0[0]
port 31 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 sram_din0[10]
port 32 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 33 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 34 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 sram_din0[13]
port 35 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 sram_din0[14]
port 36 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 sram_din0[15]
port 37 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 sram_din0[16]
port 38 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 sram_din0[17]
port 39 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 sram_din0[18]
port 40 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 sram_din0[19]
port 41 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 sram_din0[1]
port 42 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 sram_din0[20]
port 43 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 sram_din0[21]
port 44 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 sram_din0[22]
port 45 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 sram_din0[23]
port 46 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 sram_din0[24]
port 47 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 sram_din0[25]
port 48 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 sram_din0[26]
port 49 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 sram_din0[27]
port 50 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 sram_din0[28]
port 51 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 sram_din0[29]
port 52 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 sram_din0[2]
port 53 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 sram_din0[30]
port 54 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 sram_din0[31]
port 55 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 sram_din0[3]
port 56 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 sram_din0[4]
port 57 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 sram_din0[5]
port 58 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 sram_din0[6]
port 59 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 sram_din0[7]
port 60 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 sram_din0[8]
port 61 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 sram_din0[9]
port 62 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 sram_dout0[0]
port 63 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 sram_dout0[10]
port 64 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 65 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 sram_dout0[12]
port 66 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sram_dout0[13]
port 67 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 sram_dout0[14]
port 68 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout0[15]
port 69 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 sram_dout0[16]
port 70 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout0[17]
port 71 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 sram_dout0[18]
port 72 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 sram_dout0[19]
port 73 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 sram_dout0[1]
port 74 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[20]
port 75 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 sram_dout0[21]
port 76 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 sram_dout0[22]
port 77 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout0[23]
port 78 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 sram_dout0[24]
port 79 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 sram_dout0[25]
port 80 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 sram_dout0[26]
port 81 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 sram_dout0[27]
port 82 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[28]
port 83 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout0[29]
port 84 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 sram_dout0[2]
port 85 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 sram_dout0[30]
port 86 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 sram_dout0[31]
port 87 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 sram_dout0[3]
port 88 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 sram_dout0[4]
port 89 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 sram_dout0[5]
port 90 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 sram_dout0[6]
port 91 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 sram_dout0[7]
port 92 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 sram_dout0[8]
port 93 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 sram_dout0[9]
port 94 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 sram_dout1[0]
port 95 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 sram_dout1[10]
port 96 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 97 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 sram_dout1[12]
port 98 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 sram_dout1[13]
port 99 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 sram_dout1[14]
port 100 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 sram_dout1[15]
port 101 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 sram_dout1[16]
port 102 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 sram_dout1[17]
port 103 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 sram_dout1[18]
port 104 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 sram_dout1[19]
port 105 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 sram_dout1[1]
port 106 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 sram_dout1[20]
port 107 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 sram_dout1[21]
port 108 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout1[22]
port 109 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 sram_dout1[23]
port 110 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 sram_dout1[24]
port 111 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 sram_dout1[25]
port 112 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[26]
port 113 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[27]
port 114 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[28]
port 115 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 sram_dout1[29]
port 116 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 sram_dout1[2]
port 117 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 sram_dout1[30]
port 118 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 sram_dout1[31]
port 119 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 sram_dout1[3]
port 120 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 sram_dout1[4]
port 121 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 sram_dout1[5]
port 122 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 sram_dout1[6]
port 123 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 sram_dout1[7]
port 124 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout1[8]
port 125 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[9]
port 126 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 sram_web0
port 127 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 sram_wmask0[0]
port 128 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 sram_wmask0[1]
port 129 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 sram_wmask0[2]
port 130 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 sram_wmask0[3]
port 131 nsew signal output
rlabel metal4 s 4208 2128 4528 39760 6 vccd1
port 132 nsew power input
rlabel metal4 s 34928 2128 35248 39760 6 vccd1
port 132 nsew power input
rlabel metal4 s 19568 2128 19888 39760 6 vssd1
port 133 nsew ground input
rlabel metal4 s 50288 2128 50608 39760 6 vssd1
port 133 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 134 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 wb_adr_i[0]
port 135 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wb_adr_i[10]
port 136 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[11]
port 137 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[12]
port 138 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[13]
port 139 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[14]
port 140 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wb_adr_i[15]
port 141 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wb_adr_i[16]
port 142 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wb_adr_i[17]
port 143 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wb_adr_i[18]
port 144 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_adr_i[19]
port 145 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wb_adr_i[1]
port 146 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_adr_i[20]
port 147 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_adr_i[21]
port 148 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_adr_i[22]
port 149 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[23]
port 150 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_adr_i[2]
port 151 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_adr_i[3]
port 152 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wb_adr_i[4]
port 153 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 wb_adr_i[5]
port 154 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wb_adr_i[6]
port 155 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wb_adr_i[7]
port 156 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wb_adr_i[8]
port 157 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wb_adr_i[9]
port 158 nsew signal input
rlabel metal3 s 0 552 800 672 6 wb_clk_i
port 159 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wb_cyc_i
port 160 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 wb_data_i[0]
port 161 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_data_i[10]
port 162 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[11]
port 163 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[12]
port 164 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[13]
port 165 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[14]
port 166 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[15]
port 167 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[16]
port 168 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wb_data_i[17]
port 169 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wb_data_i[18]
port 170 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wb_data_i[19]
port 171 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wb_data_i[1]
port 172 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[20]
port 173 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wb_data_i[21]
port 174 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wb_data_i[22]
port 175 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_data_i[23]
port 176 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wb_data_i[24]
port 177 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 wb_data_i[25]
port 178 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 wb_data_i[26]
port 179 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 wb_data_i[27]
port 180 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_data_i[28]
port 181 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 wb_data_i[29]
port 182 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wb_data_i[2]
port 183 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 wb_data_i[30]
port 184 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 wb_data_i[31]
port 185 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wb_data_i[3]
port 186 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_data_i[4]
port 187 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_data_i[5]
port 188 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_data_i[6]
port 189 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wb_data_i[7]
port 190 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wb_data_i[8]
port 191 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wb_data_i[9]
port 192 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 wb_data_o[0]
port 193 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 wb_data_o[10]
port 194 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[11]
port 195 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[12]
port 196 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[13]
port 197 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 wb_data_o[14]
port 198 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 wb_data_o[15]
port 199 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 wb_data_o[16]
port 200 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 wb_data_o[17]
port 201 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 wb_data_o[18]
port 202 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 wb_data_o[19]
port 203 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 wb_data_o[1]
port 204 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 wb_data_o[20]
port 205 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[21]
port 206 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 wb_data_o[22]
port 207 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 wb_data_o[23]
port 208 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 wb_data_o[24]
port 209 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 wb_data_o[25]
port 210 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 wb_data_o[26]
port 211 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 wb_data_o[27]
port 212 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 wb_data_o[28]
port 213 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 wb_data_o[29]
port 214 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 wb_data_o[2]
port 215 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 wb_data_o[30]
port 216 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 wb_data_o[31]
port 217 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 wb_data_o[3]
port 218 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 wb_data_o[4]
port 219 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 wb_data_o[5]
port 220 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 wb_data_o[6]
port 221 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 wb_data_o[7]
port 222 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 wb_data_o[8]
port 223 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 wb_data_o[9]
port 224 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 wb_error_o
port 225 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 wb_rst_i
port 226 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wb_sel_i[0]
port 227 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wb_sel_i[1]
port 228 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 wb_sel_i[2]
port 229 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_sel_i[3]
port 230 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_stall_o
port 231 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 wb_stb_i
port 232 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 wb_we_i
port 233 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3537982
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Flash/runs/Flash/results/finishing/Flash.magic.gds
string GDS_START 532464
<< end >>

