magic
tech sky130A
magscale 1 2
timestamp 1652654224
<< viali >>
rect 7481 22185 7515 22219
rect 6837 22049 6871 22083
rect 8125 21913 8159 21947
rect 8125 21641 8159 21675
rect 6837 21505 6871 21539
rect 7481 21369 7515 21403
rect 7481 21097 7515 21131
rect 8125 20893 8159 20927
rect 8125 20349 8159 20383
rect 8125 19737 8159 19771
rect 8125 19329 8159 19363
rect 7481 19193 7515 19227
rect 8125 18717 8159 18751
rect 8125 18173 8159 18207
rect 8125 17629 8159 17663
rect 8125 17085 8159 17119
rect 8125 16609 8159 16643
rect 8125 15997 8159 16031
rect 8125 15453 8159 15487
rect 8125 14909 8159 14943
rect 8125 14365 8159 14399
rect 8125 13821 8159 13855
rect 8125 13277 8159 13311
rect 8125 12597 8159 12631
rect 8125 12189 8159 12223
rect 8125 11509 8159 11543
rect 8125 11101 8159 11135
rect 8125 10421 8159 10455
rect 8125 10013 8159 10047
rect 8125 9333 8159 9367
rect 8125 8925 8159 8959
rect 8125 8313 8159 8347
rect 8125 7837 8159 7871
rect 8125 7157 8159 7191
rect 8125 6749 8159 6783
rect 8125 6069 8159 6103
rect 8125 5661 8159 5695
rect 8125 4981 8159 5015
rect 8125 4437 8159 4471
rect 7481 3893 7515 3927
rect 8125 3893 8159 3927
rect 7481 3485 7515 3519
rect 8125 3485 8159 3519
rect 7481 2805 7515 2839
rect 8125 2805 8159 2839
rect 7481 2397 7515 2431
rect 8125 2397 8159 2431
<< metal1 >>
rect 1104 22330 8832 22352
rect 1104 22278 2248 22330
rect 2300 22278 2312 22330
rect 2364 22278 2376 22330
rect 2428 22278 2440 22330
rect 2492 22278 2504 22330
rect 2556 22278 4846 22330
rect 4898 22278 4910 22330
rect 4962 22278 4974 22330
rect 5026 22278 5038 22330
rect 5090 22278 5102 22330
rect 5154 22278 7443 22330
rect 7495 22278 7507 22330
rect 7559 22278 7571 22330
rect 7623 22278 7635 22330
rect 7687 22278 7699 22330
rect 7751 22278 8832 22330
rect 1104 22256 8832 22278
rect 6822 22176 6828 22228
rect 6880 22216 6886 22228
rect 7469 22219 7527 22225
rect 7469 22216 7481 22219
rect 6880 22188 7481 22216
rect 6880 22176 6886 22188
rect 7469 22185 7481 22188
rect 7515 22185 7527 22219
rect 7469 22179 7527 22185
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 6788 22120 6868 22148
rect 6788 22108 6794 22120
rect 6840 22089 6868 22120
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22049 6883 22083
rect 6825 22043 6883 22049
rect 8110 21944 8116 21956
rect 8071 21916 8116 21944
rect 8110 21904 8116 21916
rect 8168 21904 8174 21956
rect 1104 21786 8832 21808
rect 1104 21734 3547 21786
rect 3599 21734 3611 21786
rect 3663 21734 3675 21786
rect 3727 21734 3739 21786
rect 3791 21734 3803 21786
rect 3855 21734 6144 21786
rect 6196 21734 6208 21786
rect 6260 21734 6272 21786
rect 6324 21734 6336 21786
rect 6388 21734 6400 21786
rect 6452 21734 8832 21786
rect 1104 21712 8832 21734
rect 8113 21675 8171 21681
rect 8113 21641 8125 21675
rect 8159 21672 8171 21675
rect 8202 21672 8208 21684
rect 8159 21644 8208 21672
rect 8159 21641 8171 21644
rect 8113 21635 8171 21641
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 6638 21496 6644 21548
rect 6696 21536 6702 21548
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 6696 21508 6837 21536
rect 6696 21496 6702 21508
rect 6825 21505 6837 21508
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 7466 21400 7472 21412
rect 7427 21372 7472 21400
rect 7466 21360 7472 21372
rect 7524 21360 7530 21412
rect 1104 21242 8832 21264
rect 1104 21190 2248 21242
rect 2300 21190 2312 21242
rect 2364 21190 2376 21242
rect 2428 21190 2440 21242
rect 2492 21190 2504 21242
rect 2556 21190 4846 21242
rect 4898 21190 4910 21242
rect 4962 21190 4974 21242
rect 5026 21190 5038 21242
rect 5090 21190 5102 21242
rect 5154 21190 7443 21242
rect 7495 21190 7507 21242
rect 7559 21190 7571 21242
rect 7623 21190 7635 21242
rect 7687 21190 7699 21242
rect 7751 21190 8832 21242
rect 1104 21168 8832 21190
rect 7469 21131 7527 21137
rect 7469 21097 7481 21131
rect 7515 21128 7527 21131
rect 7834 21128 7840 21140
rect 7515 21100 7840 21128
rect 7515 21097 7527 21100
rect 7469 21091 7527 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 8110 20924 8116 20936
rect 8071 20896 8116 20924
rect 8110 20884 8116 20896
rect 8168 20884 8174 20936
rect 1104 20698 8832 20720
rect 1104 20646 3547 20698
rect 3599 20646 3611 20698
rect 3663 20646 3675 20698
rect 3727 20646 3739 20698
rect 3791 20646 3803 20698
rect 3855 20646 6144 20698
rect 6196 20646 6208 20698
rect 6260 20646 6272 20698
rect 6324 20646 6336 20698
rect 6388 20646 6400 20698
rect 6452 20646 8832 20698
rect 1104 20624 8832 20646
rect 8110 20380 8116 20392
rect 8071 20352 8116 20380
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 1104 20154 8832 20176
rect 1104 20102 2248 20154
rect 2300 20102 2312 20154
rect 2364 20102 2376 20154
rect 2428 20102 2440 20154
rect 2492 20102 2504 20154
rect 2556 20102 4846 20154
rect 4898 20102 4910 20154
rect 4962 20102 4974 20154
rect 5026 20102 5038 20154
rect 5090 20102 5102 20154
rect 5154 20102 7443 20154
rect 7495 20102 7507 20154
rect 7559 20102 7571 20154
rect 7623 20102 7635 20154
rect 7687 20102 7699 20154
rect 7751 20102 8832 20154
rect 1104 20080 8832 20102
rect 8110 19768 8116 19780
rect 8071 19740 8116 19768
rect 8110 19728 8116 19740
rect 8168 19728 8174 19780
rect 1104 19610 8832 19632
rect 1104 19558 3547 19610
rect 3599 19558 3611 19610
rect 3663 19558 3675 19610
rect 3727 19558 3739 19610
rect 3791 19558 3803 19610
rect 3855 19558 6144 19610
rect 6196 19558 6208 19610
rect 6260 19558 6272 19610
rect 6324 19558 6336 19610
rect 6388 19558 6400 19610
rect 6452 19558 8832 19610
rect 1104 19536 8832 19558
rect 8110 19360 8116 19372
rect 8071 19332 8116 19360
rect 8110 19320 8116 19332
rect 8168 19320 8174 19372
rect 7466 19224 7472 19236
rect 7427 19196 7472 19224
rect 7466 19184 7472 19196
rect 7524 19184 7530 19236
rect 1104 19066 8832 19088
rect 1104 19014 2248 19066
rect 2300 19014 2312 19066
rect 2364 19014 2376 19066
rect 2428 19014 2440 19066
rect 2492 19014 2504 19066
rect 2556 19014 4846 19066
rect 4898 19014 4910 19066
rect 4962 19014 4974 19066
rect 5026 19014 5038 19066
rect 5090 19014 5102 19066
rect 5154 19014 7443 19066
rect 7495 19014 7507 19066
rect 7559 19014 7571 19066
rect 7623 19014 7635 19066
rect 7687 19014 7699 19066
rect 7751 19014 8832 19066
rect 1104 18992 8832 19014
rect 8110 18748 8116 18760
rect 8071 18720 8116 18748
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 1104 18522 8832 18544
rect 1104 18470 3547 18522
rect 3599 18470 3611 18522
rect 3663 18470 3675 18522
rect 3727 18470 3739 18522
rect 3791 18470 3803 18522
rect 3855 18470 6144 18522
rect 6196 18470 6208 18522
rect 6260 18470 6272 18522
rect 6324 18470 6336 18522
rect 6388 18470 6400 18522
rect 6452 18470 8832 18522
rect 1104 18448 8832 18470
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 1104 17978 8832 18000
rect 1104 17926 2248 17978
rect 2300 17926 2312 17978
rect 2364 17926 2376 17978
rect 2428 17926 2440 17978
rect 2492 17926 2504 17978
rect 2556 17926 4846 17978
rect 4898 17926 4910 17978
rect 4962 17926 4974 17978
rect 5026 17926 5038 17978
rect 5090 17926 5102 17978
rect 5154 17926 7443 17978
rect 7495 17926 7507 17978
rect 7559 17926 7571 17978
rect 7623 17926 7635 17978
rect 7687 17926 7699 17978
rect 7751 17926 8832 17978
rect 1104 17904 8832 17926
rect 8110 17660 8116 17672
rect 8071 17632 8116 17660
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 1104 17434 8832 17456
rect 1104 17382 3547 17434
rect 3599 17382 3611 17434
rect 3663 17382 3675 17434
rect 3727 17382 3739 17434
rect 3791 17382 3803 17434
rect 3855 17382 6144 17434
rect 6196 17382 6208 17434
rect 6260 17382 6272 17434
rect 6324 17382 6336 17434
rect 6388 17382 6400 17434
rect 6452 17382 8832 17434
rect 1104 17360 8832 17382
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17116 8171 17119
rect 8202 17116 8208 17128
rect 8159 17088 8208 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 1104 16890 8832 16912
rect 1104 16838 2248 16890
rect 2300 16838 2312 16890
rect 2364 16838 2376 16890
rect 2428 16838 2440 16890
rect 2492 16838 2504 16890
rect 2556 16838 4846 16890
rect 4898 16838 4910 16890
rect 4962 16838 4974 16890
rect 5026 16838 5038 16890
rect 5090 16838 5102 16890
rect 5154 16838 7443 16890
rect 7495 16838 7507 16890
rect 7559 16838 7571 16890
rect 7623 16838 7635 16890
rect 7687 16838 7699 16890
rect 7751 16838 8832 16890
rect 1104 16816 8832 16838
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 1104 16346 8832 16368
rect 1104 16294 3547 16346
rect 3599 16294 3611 16346
rect 3663 16294 3675 16346
rect 3727 16294 3739 16346
rect 3791 16294 3803 16346
rect 3855 16294 6144 16346
rect 6196 16294 6208 16346
rect 6260 16294 6272 16346
rect 6324 16294 6336 16346
rect 6388 16294 6400 16346
rect 6452 16294 8832 16346
rect 1104 16272 8832 16294
rect 8110 16028 8116 16040
rect 8071 16000 8116 16028
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 1104 15802 8832 15824
rect 1104 15750 2248 15802
rect 2300 15750 2312 15802
rect 2364 15750 2376 15802
rect 2428 15750 2440 15802
rect 2492 15750 2504 15802
rect 2556 15750 4846 15802
rect 4898 15750 4910 15802
rect 4962 15750 4974 15802
rect 5026 15750 5038 15802
rect 5090 15750 5102 15802
rect 5154 15750 7443 15802
rect 7495 15750 7507 15802
rect 7559 15750 7571 15802
rect 7623 15750 7635 15802
rect 7687 15750 7699 15802
rect 7751 15750 8832 15802
rect 1104 15728 8832 15750
rect 8110 15484 8116 15496
rect 8071 15456 8116 15484
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 1104 15258 8832 15280
rect 1104 15206 3547 15258
rect 3599 15206 3611 15258
rect 3663 15206 3675 15258
rect 3727 15206 3739 15258
rect 3791 15206 3803 15258
rect 3855 15206 6144 15258
rect 6196 15206 6208 15258
rect 6260 15206 6272 15258
rect 6324 15206 6336 15258
rect 6388 15206 6400 15258
rect 6452 15206 8832 15258
rect 1104 15184 8832 15206
rect 8110 14940 8116 14952
rect 8071 14912 8116 14940
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 1104 14714 8832 14736
rect 1104 14662 2248 14714
rect 2300 14662 2312 14714
rect 2364 14662 2376 14714
rect 2428 14662 2440 14714
rect 2492 14662 2504 14714
rect 2556 14662 4846 14714
rect 4898 14662 4910 14714
rect 4962 14662 4974 14714
rect 5026 14662 5038 14714
rect 5090 14662 5102 14714
rect 5154 14662 7443 14714
rect 7495 14662 7507 14714
rect 7559 14662 7571 14714
rect 7623 14662 7635 14714
rect 7687 14662 7699 14714
rect 7751 14662 8832 14714
rect 1104 14640 8832 14662
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 1104 14170 8832 14192
rect 1104 14118 3547 14170
rect 3599 14118 3611 14170
rect 3663 14118 3675 14170
rect 3727 14118 3739 14170
rect 3791 14118 3803 14170
rect 3855 14118 6144 14170
rect 6196 14118 6208 14170
rect 6260 14118 6272 14170
rect 6324 14118 6336 14170
rect 6388 14118 6400 14170
rect 6452 14118 8832 14170
rect 1104 14096 8832 14118
rect 8110 13852 8116 13864
rect 8071 13824 8116 13852
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 1104 13626 8832 13648
rect 1104 13574 2248 13626
rect 2300 13574 2312 13626
rect 2364 13574 2376 13626
rect 2428 13574 2440 13626
rect 2492 13574 2504 13626
rect 2556 13574 4846 13626
rect 4898 13574 4910 13626
rect 4962 13574 4974 13626
rect 5026 13574 5038 13626
rect 5090 13574 5102 13626
rect 5154 13574 7443 13626
rect 7495 13574 7507 13626
rect 7559 13574 7571 13626
rect 7623 13574 7635 13626
rect 7687 13574 7699 13626
rect 7751 13574 8832 13626
rect 1104 13552 8832 13574
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 1104 13082 8832 13104
rect 1104 13030 3547 13082
rect 3599 13030 3611 13082
rect 3663 13030 3675 13082
rect 3727 13030 3739 13082
rect 3791 13030 3803 13082
rect 3855 13030 6144 13082
rect 6196 13030 6208 13082
rect 6260 13030 6272 13082
rect 6324 13030 6336 13082
rect 6388 13030 6400 13082
rect 6452 13030 8832 13082
rect 1104 13008 8832 13030
rect 8110 12628 8116 12640
rect 8071 12600 8116 12628
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 1104 12538 8832 12560
rect 1104 12486 2248 12538
rect 2300 12486 2312 12538
rect 2364 12486 2376 12538
rect 2428 12486 2440 12538
rect 2492 12486 2504 12538
rect 2556 12486 4846 12538
rect 4898 12486 4910 12538
rect 4962 12486 4974 12538
rect 5026 12486 5038 12538
rect 5090 12486 5102 12538
rect 5154 12486 7443 12538
rect 7495 12486 7507 12538
rect 7559 12486 7571 12538
rect 7623 12486 7635 12538
rect 7687 12486 7699 12538
rect 7751 12486 8832 12538
rect 1104 12464 8832 12486
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 1104 11994 8832 12016
rect 1104 11942 3547 11994
rect 3599 11942 3611 11994
rect 3663 11942 3675 11994
rect 3727 11942 3739 11994
rect 3791 11942 3803 11994
rect 3855 11942 6144 11994
rect 6196 11942 6208 11994
rect 6260 11942 6272 11994
rect 6324 11942 6336 11994
rect 6388 11942 6400 11994
rect 6452 11942 8832 11994
rect 1104 11920 8832 11942
rect 8110 11540 8116 11552
rect 8071 11512 8116 11540
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 1104 11450 8832 11472
rect 1104 11398 2248 11450
rect 2300 11398 2312 11450
rect 2364 11398 2376 11450
rect 2428 11398 2440 11450
rect 2492 11398 2504 11450
rect 2556 11398 4846 11450
rect 4898 11398 4910 11450
rect 4962 11398 4974 11450
rect 5026 11398 5038 11450
rect 5090 11398 5102 11450
rect 5154 11398 7443 11450
rect 7495 11398 7507 11450
rect 7559 11398 7571 11450
rect 7623 11398 7635 11450
rect 7687 11398 7699 11450
rect 7751 11398 8832 11450
rect 1104 11376 8832 11398
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 1104 10906 8832 10928
rect 1104 10854 3547 10906
rect 3599 10854 3611 10906
rect 3663 10854 3675 10906
rect 3727 10854 3739 10906
rect 3791 10854 3803 10906
rect 3855 10854 6144 10906
rect 6196 10854 6208 10906
rect 6260 10854 6272 10906
rect 6324 10854 6336 10906
rect 6388 10854 6400 10906
rect 6452 10854 8832 10906
rect 1104 10832 8832 10854
rect 8110 10452 8116 10464
rect 8071 10424 8116 10452
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 1104 10362 8832 10384
rect 1104 10310 2248 10362
rect 2300 10310 2312 10362
rect 2364 10310 2376 10362
rect 2428 10310 2440 10362
rect 2492 10310 2504 10362
rect 2556 10310 4846 10362
rect 4898 10310 4910 10362
rect 4962 10310 4974 10362
rect 5026 10310 5038 10362
rect 5090 10310 5102 10362
rect 5154 10310 7443 10362
rect 7495 10310 7507 10362
rect 7559 10310 7571 10362
rect 7623 10310 7635 10362
rect 7687 10310 7699 10362
rect 7751 10310 8832 10362
rect 1104 10288 8832 10310
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 1104 9818 8832 9840
rect 1104 9766 3547 9818
rect 3599 9766 3611 9818
rect 3663 9766 3675 9818
rect 3727 9766 3739 9818
rect 3791 9766 3803 9818
rect 3855 9766 6144 9818
rect 6196 9766 6208 9818
rect 6260 9766 6272 9818
rect 6324 9766 6336 9818
rect 6388 9766 6400 9818
rect 6452 9766 8832 9818
rect 1104 9744 8832 9766
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 1104 9274 8832 9296
rect 1104 9222 2248 9274
rect 2300 9222 2312 9274
rect 2364 9222 2376 9274
rect 2428 9222 2440 9274
rect 2492 9222 2504 9274
rect 2556 9222 4846 9274
rect 4898 9222 4910 9274
rect 4962 9222 4974 9274
rect 5026 9222 5038 9274
rect 5090 9222 5102 9274
rect 5154 9222 7443 9274
rect 7495 9222 7507 9274
rect 7559 9222 7571 9274
rect 7623 9222 7635 9274
rect 7687 9222 7699 9274
rect 7751 9222 8832 9274
rect 1104 9200 8832 9222
rect 8110 8956 8116 8968
rect 8071 8928 8116 8956
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 1104 8730 8832 8752
rect 1104 8678 3547 8730
rect 3599 8678 3611 8730
rect 3663 8678 3675 8730
rect 3727 8678 3739 8730
rect 3791 8678 3803 8730
rect 3855 8678 6144 8730
rect 6196 8678 6208 8730
rect 6260 8678 6272 8730
rect 6324 8678 6336 8730
rect 6388 8678 6400 8730
rect 6452 8678 8832 8730
rect 1104 8656 8832 8678
rect 8110 8344 8116 8356
rect 8071 8316 8116 8344
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 1104 8186 8832 8208
rect 1104 8134 2248 8186
rect 2300 8134 2312 8186
rect 2364 8134 2376 8186
rect 2428 8134 2440 8186
rect 2492 8134 2504 8186
rect 2556 8134 4846 8186
rect 4898 8134 4910 8186
rect 4962 8134 4974 8186
rect 5026 8134 5038 8186
rect 5090 8134 5102 8186
rect 5154 8134 7443 8186
rect 7495 8134 7507 8186
rect 7559 8134 7571 8186
rect 7623 8134 7635 8186
rect 7687 8134 7699 8186
rect 7751 8134 8832 8186
rect 1104 8112 8832 8134
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 1104 7642 8832 7664
rect 1104 7590 3547 7642
rect 3599 7590 3611 7642
rect 3663 7590 3675 7642
rect 3727 7590 3739 7642
rect 3791 7590 3803 7642
rect 3855 7590 6144 7642
rect 6196 7590 6208 7642
rect 6260 7590 6272 7642
rect 6324 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 8832 7642
rect 1104 7568 8832 7590
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 1104 7098 8832 7120
rect 1104 7046 2248 7098
rect 2300 7046 2312 7098
rect 2364 7046 2376 7098
rect 2428 7046 2440 7098
rect 2492 7046 2504 7098
rect 2556 7046 4846 7098
rect 4898 7046 4910 7098
rect 4962 7046 4974 7098
rect 5026 7046 5038 7098
rect 5090 7046 5102 7098
rect 5154 7046 7443 7098
rect 7495 7046 7507 7098
rect 7559 7046 7571 7098
rect 7623 7046 7635 7098
rect 7687 7046 7699 7098
rect 7751 7046 8832 7098
rect 1104 7024 8832 7046
rect 8110 6780 8116 6792
rect 8071 6752 8116 6780
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 1104 6554 8832 6576
rect 1104 6502 3547 6554
rect 3599 6502 3611 6554
rect 3663 6502 3675 6554
rect 3727 6502 3739 6554
rect 3791 6502 3803 6554
rect 3855 6502 6144 6554
rect 6196 6502 6208 6554
rect 6260 6502 6272 6554
rect 6324 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 8832 6554
rect 1104 6480 8832 6502
rect 8110 6100 8116 6112
rect 8071 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 1104 6010 8832 6032
rect 1104 5958 2248 6010
rect 2300 5958 2312 6010
rect 2364 5958 2376 6010
rect 2428 5958 2440 6010
rect 2492 5958 2504 6010
rect 2556 5958 4846 6010
rect 4898 5958 4910 6010
rect 4962 5958 4974 6010
rect 5026 5958 5038 6010
rect 5090 5958 5102 6010
rect 5154 5958 7443 6010
rect 7495 5958 7507 6010
rect 7559 5958 7571 6010
rect 7623 5958 7635 6010
rect 7687 5958 7699 6010
rect 7751 5958 8832 6010
rect 1104 5936 8832 5958
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 1104 5466 8832 5488
rect 1104 5414 3547 5466
rect 3599 5414 3611 5466
rect 3663 5414 3675 5466
rect 3727 5414 3739 5466
rect 3791 5414 3803 5466
rect 3855 5414 6144 5466
rect 6196 5414 6208 5466
rect 6260 5414 6272 5466
rect 6324 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 8832 5466
rect 1104 5392 8832 5414
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 1104 4922 8832 4944
rect 1104 4870 2248 4922
rect 2300 4870 2312 4922
rect 2364 4870 2376 4922
rect 2428 4870 2440 4922
rect 2492 4870 2504 4922
rect 2556 4870 4846 4922
rect 4898 4870 4910 4922
rect 4962 4870 4974 4922
rect 5026 4870 5038 4922
rect 5090 4870 5102 4922
rect 5154 4870 7443 4922
rect 7495 4870 7507 4922
rect 7559 4870 7571 4922
rect 7623 4870 7635 4922
rect 7687 4870 7699 4922
rect 7751 4870 8832 4922
rect 1104 4848 8832 4870
rect 8110 4468 8116 4480
rect 8071 4440 8116 4468
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 1104 4378 8832 4400
rect 1104 4326 3547 4378
rect 3599 4326 3611 4378
rect 3663 4326 3675 4378
rect 3727 4326 3739 4378
rect 3791 4326 3803 4378
rect 3855 4326 6144 4378
rect 6196 4326 6208 4378
rect 6260 4326 6272 4378
rect 6324 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 8832 4378
rect 1104 4304 8832 4326
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 7834 3924 7840 3936
rect 7515 3896 7840 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 1104 3834 8832 3856
rect 1104 3782 2248 3834
rect 2300 3782 2312 3834
rect 2364 3782 2376 3834
rect 2428 3782 2440 3834
rect 2492 3782 2504 3834
rect 2556 3782 4846 3834
rect 4898 3782 4910 3834
rect 4962 3782 4974 3834
rect 5026 3782 5038 3834
rect 5090 3782 5102 3834
rect 5154 3782 7443 3834
rect 7495 3782 7507 3834
rect 7559 3782 7571 3834
rect 7623 3782 7635 3834
rect 7687 3782 7699 3834
rect 7751 3782 8832 3834
rect 1104 3760 8832 3782
rect 7466 3516 7472 3528
rect 7427 3488 7472 3516
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8202 3516 8208 3528
rect 8159 3488 8208 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 1104 3290 8832 3312
rect 1104 3238 3547 3290
rect 3599 3238 3611 3290
rect 3663 3238 3675 3290
rect 3727 3238 3739 3290
rect 3791 3238 3803 3290
rect 3855 3238 6144 3290
rect 6196 3238 6208 3290
rect 6260 3238 6272 3290
rect 6324 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 8832 3290
rect 1104 3216 8832 3238
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 7834 2836 7840 2848
rect 7515 2808 7840 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 8076 2808 8125 2836
rect 8076 2796 8082 2808
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8113 2799 8171 2805
rect 1104 2746 8832 2768
rect 1104 2694 2248 2746
rect 2300 2694 2312 2746
rect 2364 2694 2376 2746
rect 2428 2694 2440 2746
rect 2492 2694 2504 2746
rect 2556 2694 4846 2746
rect 4898 2694 4910 2746
rect 4962 2694 4974 2746
rect 5026 2694 5038 2746
rect 5090 2694 5102 2746
rect 5154 2694 7443 2746
rect 7495 2694 7507 2746
rect 7559 2694 7571 2746
rect 7623 2694 7635 2746
rect 7687 2694 7699 2746
rect 7751 2694 8832 2746
rect 1104 2672 8832 2694
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8110 2428 8116 2440
rect 8071 2400 8116 2428
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 1104 2202 8832 2224
rect 1104 2150 3547 2202
rect 3599 2150 3611 2202
rect 3663 2150 3675 2202
rect 3727 2150 3739 2202
rect 3791 2150 3803 2202
rect 3855 2150 6144 2202
rect 6196 2150 6208 2202
rect 6260 2150 6272 2202
rect 6324 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 2248 22278 2300 22330
rect 2312 22278 2364 22330
rect 2376 22278 2428 22330
rect 2440 22278 2492 22330
rect 2504 22278 2556 22330
rect 4846 22278 4898 22330
rect 4910 22278 4962 22330
rect 4974 22278 5026 22330
rect 5038 22278 5090 22330
rect 5102 22278 5154 22330
rect 7443 22278 7495 22330
rect 7507 22278 7559 22330
rect 7571 22278 7623 22330
rect 7635 22278 7687 22330
rect 7699 22278 7751 22330
rect 6828 22176 6880 22228
rect 6736 22108 6788 22160
rect 8116 21947 8168 21956
rect 8116 21913 8125 21947
rect 8125 21913 8159 21947
rect 8159 21913 8168 21947
rect 8116 21904 8168 21913
rect 3547 21734 3599 21786
rect 3611 21734 3663 21786
rect 3675 21734 3727 21786
rect 3739 21734 3791 21786
rect 3803 21734 3855 21786
rect 6144 21734 6196 21786
rect 6208 21734 6260 21786
rect 6272 21734 6324 21786
rect 6336 21734 6388 21786
rect 6400 21734 6452 21786
rect 8208 21632 8260 21684
rect 6644 21496 6696 21548
rect 7472 21403 7524 21412
rect 7472 21369 7481 21403
rect 7481 21369 7515 21403
rect 7515 21369 7524 21403
rect 7472 21360 7524 21369
rect 2248 21190 2300 21242
rect 2312 21190 2364 21242
rect 2376 21190 2428 21242
rect 2440 21190 2492 21242
rect 2504 21190 2556 21242
rect 4846 21190 4898 21242
rect 4910 21190 4962 21242
rect 4974 21190 5026 21242
rect 5038 21190 5090 21242
rect 5102 21190 5154 21242
rect 7443 21190 7495 21242
rect 7507 21190 7559 21242
rect 7571 21190 7623 21242
rect 7635 21190 7687 21242
rect 7699 21190 7751 21242
rect 7840 21088 7892 21140
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 3547 20646 3599 20698
rect 3611 20646 3663 20698
rect 3675 20646 3727 20698
rect 3739 20646 3791 20698
rect 3803 20646 3855 20698
rect 6144 20646 6196 20698
rect 6208 20646 6260 20698
rect 6272 20646 6324 20698
rect 6336 20646 6388 20698
rect 6400 20646 6452 20698
rect 8116 20383 8168 20392
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 2248 20102 2300 20154
rect 2312 20102 2364 20154
rect 2376 20102 2428 20154
rect 2440 20102 2492 20154
rect 2504 20102 2556 20154
rect 4846 20102 4898 20154
rect 4910 20102 4962 20154
rect 4974 20102 5026 20154
rect 5038 20102 5090 20154
rect 5102 20102 5154 20154
rect 7443 20102 7495 20154
rect 7507 20102 7559 20154
rect 7571 20102 7623 20154
rect 7635 20102 7687 20154
rect 7699 20102 7751 20154
rect 8116 19771 8168 19780
rect 8116 19737 8125 19771
rect 8125 19737 8159 19771
rect 8159 19737 8168 19771
rect 8116 19728 8168 19737
rect 3547 19558 3599 19610
rect 3611 19558 3663 19610
rect 3675 19558 3727 19610
rect 3739 19558 3791 19610
rect 3803 19558 3855 19610
rect 6144 19558 6196 19610
rect 6208 19558 6260 19610
rect 6272 19558 6324 19610
rect 6336 19558 6388 19610
rect 6400 19558 6452 19610
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 8116 19320 8168 19329
rect 7472 19227 7524 19236
rect 7472 19193 7481 19227
rect 7481 19193 7515 19227
rect 7515 19193 7524 19227
rect 7472 19184 7524 19193
rect 2248 19014 2300 19066
rect 2312 19014 2364 19066
rect 2376 19014 2428 19066
rect 2440 19014 2492 19066
rect 2504 19014 2556 19066
rect 4846 19014 4898 19066
rect 4910 19014 4962 19066
rect 4974 19014 5026 19066
rect 5038 19014 5090 19066
rect 5102 19014 5154 19066
rect 7443 19014 7495 19066
rect 7507 19014 7559 19066
rect 7571 19014 7623 19066
rect 7635 19014 7687 19066
rect 7699 19014 7751 19066
rect 8116 18751 8168 18760
rect 8116 18717 8125 18751
rect 8125 18717 8159 18751
rect 8159 18717 8168 18751
rect 8116 18708 8168 18717
rect 3547 18470 3599 18522
rect 3611 18470 3663 18522
rect 3675 18470 3727 18522
rect 3739 18470 3791 18522
rect 3803 18470 3855 18522
rect 6144 18470 6196 18522
rect 6208 18470 6260 18522
rect 6272 18470 6324 18522
rect 6336 18470 6388 18522
rect 6400 18470 6452 18522
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 2248 17926 2300 17978
rect 2312 17926 2364 17978
rect 2376 17926 2428 17978
rect 2440 17926 2492 17978
rect 2504 17926 2556 17978
rect 4846 17926 4898 17978
rect 4910 17926 4962 17978
rect 4974 17926 5026 17978
rect 5038 17926 5090 17978
rect 5102 17926 5154 17978
rect 7443 17926 7495 17978
rect 7507 17926 7559 17978
rect 7571 17926 7623 17978
rect 7635 17926 7687 17978
rect 7699 17926 7751 17978
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 3547 17382 3599 17434
rect 3611 17382 3663 17434
rect 3675 17382 3727 17434
rect 3739 17382 3791 17434
rect 3803 17382 3855 17434
rect 6144 17382 6196 17434
rect 6208 17382 6260 17434
rect 6272 17382 6324 17434
rect 6336 17382 6388 17434
rect 6400 17382 6452 17434
rect 8208 17076 8260 17128
rect 2248 16838 2300 16890
rect 2312 16838 2364 16890
rect 2376 16838 2428 16890
rect 2440 16838 2492 16890
rect 2504 16838 2556 16890
rect 4846 16838 4898 16890
rect 4910 16838 4962 16890
rect 4974 16838 5026 16890
rect 5038 16838 5090 16890
rect 5102 16838 5154 16890
rect 7443 16838 7495 16890
rect 7507 16838 7559 16890
rect 7571 16838 7623 16890
rect 7635 16838 7687 16890
rect 7699 16838 7751 16890
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 3547 16294 3599 16346
rect 3611 16294 3663 16346
rect 3675 16294 3727 16346
rect 3739 16294 3791 16346
rect 3803 16294 3855 16346
rect 6144 16294 6196 16346
rect 6208 16294 6260 16346
rect 6272 16294 6324 16346
rect 6336 16294 6388 16346
rect 6400 16294 6452 16346
rect 8116 16031 8168 16040
rect 8116 15997 8125 16031
rect 8125 15997 8159 16031
rect 8159 15997 8168 16031
rect 8116 15988 8168 15997
rect 2248 15750 2300 15802
rect 2312 15750 2364 15802
rect 2376 15750 2428 15802
rect 2440 15750 2492 15802
rect 2504 15750 2556 15802
rect 4846 15750 4898 15802
rect 4910 15750 4962 15802
rect 4974 15750 5026 15802
rect 5038 15750 5090 15802
rect 5102 15750 5154 15802
rect 7443 15750 7495 15802
rect 7507 15750 7559 15802
rect 7571 15750 7623 15802
rect 7635 15750 7687 15802
rect 7699 15750 7751 15802
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 3547 15206 3599 15258
rect 3611 15206 3663 15258
rect 3675 15206 3727 15258
rect 3739 15206 3791 15258
rect 3803 15206 3855 15258
rect 6144 15206 6196 15258
rect 6208 15206 6260 15258
rect 6272 15206 6324 15258
rect 6336 15206 6388 15258
rect 6400 15206 6452 15258
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 2248 14662 2300 14714
rect 2312 14662 2364 14714
rect 2376 14662 2428 14714
rect 2440 14662 2492 14714
rect 2504 14662 2556 14714
rect 4846 14662 4898 14714
rect 4910 14662 4962 14714
rect 4974 14662 5026 14714
rect 5038 14662 5090 14714
rect 5102 14662 5154 14714
rect 7443 14662 7495 14714
rect 7507 14662 7559 14714
rect 7571 14662 7623 14714
rect 7635 14662 7687 14714
rect 7699 14662 7751 14714
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 3547 14118 3599 14170
rect 3611 14118 3663 14170
rect 3675 14118 3727 14170
rect 3739 14118 3791 14170
rect 3803 14118 3855 14170
rect 6144 14118 6196 14170
rect 6208 14118 6260 14170
rect 6272 14118 6324 14170
rect 6336 14118 6388 14170
rect 6400 14118 6452 14170
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 2248 13574 2300 13626
rect 2312 13574 2364 13626
rect 2376 13574 2428 13626
rect 2440 13574 2492 13626
rect 2504 13574 2556 13626
rect 4846 13574 4898 13626
rect 4910 13574 4962 13626
rect 4974 13574 5026 13626
rect 5038 13574 5090 13626
rect 5102 13574 5154 13626
rect 7443 13574 7495 13626
rect 7507 13574 7559 13626
rect 7571 13574 7623 13626
rect 7635 13574 7687 13626
rect 7699 13574 7751 13626
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 3547 13030 3599 13082
rect 3611 13030 3663 13082
rect 3675 13030 3727 13082
rect 3739 13030 3791 13082
rect 3803 13030 3855 13082
rect 6144 13030 6196 13082
rect 6208 13030 6260 13082
rect 6272 13030 6324 13082
rect 6336 13030 6388 13082
rect 6400 13030 6452 13082
rect 8116 12631 8168 12640
rect 8116 12597 8125 12631
rect 8125 12597 8159 12631
rect 8159 12597 8168 12631
rect 8116 12588 8168 12597
rect 2248 12486 2300 12538
rect 2312 12486 2364 12538
rect 2376 12486 2428 12538
rect 2440 12486 2492 12538
rect 2504 12486 2556 12538
rect 4846 12486 4898 12538
rect 4910 12486 4962 12538
rect 4974 12486 5026 12538
rect 5038 12486 5090 12538
rect 5102 12486 5154 12538
rect 7443 12486 7495 12538
rect 7507 12486 7559 12538
rect 7571 12486 7623 12538
rect 7635 12486 7687 12538
rect 7699 12486 7751 12538
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 3547 11942 3599 11994
rect 3611 11942 3663 11994
rect 3675 11942 3727 11994
rect 3739 11942 3791 11994
rect 3803 11942 3855 11994
rect 6144 11942 6196 11994
rect 6208 11942 6260 11994
rect 6272 11942 6324 11994
rect 6336 11942 6388 11994
rect 6400 11942 6452 11994
rect 8116 11543 8168 11552
rect 8116 11509 8125 11543
rect 8125 11509 8159 11543
rect 8159 11509 8168 11543
rect 8116 11500 8168 11509
rect 2248 11398 2300 11450
rect 2312 11398 2364 11450
rect 2376 11398 2428 11450
rect 2440 11398 2492 11450
rect 2504 11398 2556 11450
rect 4846 11398 4898 11450
rect 4910 11398 4962 11450
rect 4974 11398 5026 11450
rect 5038 11398 5090 11450
rect 5102 11398 5154 11450
rect 7443 11398 7495 11450
rect 7507 11398 7559 11450
rect 7571 11398 7623 11450
rect 7635 11398 7687 11450
rect 7699 11398 7751 11450
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 3547 10854 3599 10906
rect 3611 10854 3663 10906
rect 3675 10854 3727 10906
rect 3739 10854 3791 10906
rect 3803 10854 3855 10906
rect 6144 10854 6196 10906
rect 6208 10854 6260 10906
rect 6272 10854 6324 10906
rect 6336 10854 6388 10906
rect 6400 10854 6452 10906
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 2248 10310 2300 10362
rect 2312 10310 2364 10362
rect 2376 10310 2428 10362
rect 2440 10310 2492 10362
rect 2504 10310 2556 10362
rect 4846 10310 4898 10362
rect 4910 10310 4962 10362
rect 4974 10310 5026 10362
rect 5038 10310 5090 10362
rect 5102 10310 5154 10362
rect 7443 10310 7495 10362
rect 7507 10310 7559 10362
rect 7571 10310 7623 10362
rect 7635 10310 7687 10362
rect 7699 10310 7751 10362
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 3547 9766 3599 9818
rect 3611 9766 3663 9818
rect 3675 9766 3727 9818
rect 3739 9766 3791 9818
rect 3803 9766 3855 9818
rect 6144 9766 6196 9818
rect 6208 9766 6260 9818
rect 6272 9766 6324 9818
rect 6336 9766 6388 9818
rect 6400 9766 6452 9818
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 2248 9222 2300 9274
rect 2312 9222 2364 9274
rect 2376 9222 2428 9274
rect 2440 9222 2492 9274
rect 2504 9222 2556 9274
rect 4846 9222 4898 9274
rect 4910 9222 4962 9274
rect 4974 9222 5026 9274
rect 5038 9222 5090 9274
rect 5102 9222 5154 9274
rect 7443 9222 7495 9274
rect 7507 9222 7559 9274
rect 7571 9222 7623 9274
rect 7635 9222 7687 9274
rect 7699 9222 7751 9274
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 3547 8678 3599 8730
rect 3611 8678 3663 8730
rect 3675 8678 3727 8730
rect 3739 8678 3791 8730
rect 3803 8678 3855 8730
rect 6144 8678 6196 8730
rect 6208 8678 6260 8730
rect 6272 8678 6324 8730
rect 6336 8678 6388 8730
rect 6400 8678 6452 8730
rect 8116 8347 8168 8356
rect 8116 8313 8125 8347
rect 8125 8313 8159 8347
rect 8159 8313 8168 8347
rect 8116 8304 8168 8313
rect 2248 8134 2300 8186
rect 2312 8134 2364 8186
rect 2376 8134 2428 8186
rect 2440 8134 2492 8186
rect 2504 8134 2556 8186
rect 4846 8134 4898 8186
rect 4910 8134 4962 8186
rect 4974 8134 5026 8186
rect 5038 8134 5090 8186
rect 5102 8134 5154 8186
rect 7443 8134 7495 8186
rect 7507 8134 7559 8186
rect 7571 8134 7623 8186
rect 7635 8134 7687 8186
rect 7699 8134 7751 8186
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 3547 7590 3599 7642
rect 3611 7590 3663 7642
rect 3675 7590 3727 7642
rect 3739 7590 3791 7642
rect 3803 7590 3855 7642
rect 6144 7590 6196 7642
rect 6208 7590 6260 7642
rect 6272 7590 6324 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 2248 7046 2300 7098
rect 2312 7046 2364 7098
rect 2376 7046 2428 7098
rect 2440 7046 2492 7098
rect 2504 7046 2556 7098
rect 4846 7046 4898 7098
rect 4910 7046 4962 7098
rect 4974 7046 5026 7098
rect 5038 7046 5090 7098
rect 5102 7046 5154 7098
rect 7443 7046 7495 7098
rect 7507 7046 7559 7098
rect 7571 7046 7623 7098
rect 7635 7046 7687 7098
rect 7699 7046 7751 7098
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 3547 6502 3599 6554
rect 3611 6502 3663 6554
rect 3675 6502 3727 6554
rect 3739 6502 3791 6554
rect 3803 6502 3855 6554
rect 6144 6502 6196 6554
rect 6208 6502 6260 6554
rect 6272 6502 6324 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 2248 5958 2300 6010
rect 2312 5958 2364 6010
rect 2376 5958 2428 6010
rect 2440 5958 2492 6010
rect 2504 5958 2556 6010
rect 4846 5958 4898 6010
rect 4910 5958 4962 6010
rect 4974 5958 5026 6010
rect 5038 5958 5090 6010
rect 5102 5958 5154 6010
rect 7443 5958 7495 6010
rect 7507 5958 7559 6010
rect 7571 5958 7623 6010
rect 7635 5958 7687 6010
rect 7699 5958 7751 6010
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 3547 5414 3599 5466
rect 3611 5414 3663 5466
rect 3675 5414 3727 5466
rect 3739 5414 3791 5466
rect 3803 5414 3855 5466
rect 6144 5414 6196 5466
rect 6208 5414 6260 5466
rect 6272 5414 6324 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 2248 4870 2300 4922
rect 2312 4870 2364 4922
rect 2376 4870 2428 4922
rect 2440 4870 2492 4922
rect 2504 4870 2556 4922
rect 4846 4870 4898 4922
rect 4910 4870 4962 4922
rect 4974 4870 5026 4922
rect 5038 4870 5090 4922
rect 5102 4870 5154 4922
rect 7443 4870 7495 4922
rect 7507 4870 7559 4922
rect 7571 4870 7623 4922
rect 7635 4870 7687 4922
rect 7699 4870 7751 4922
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 3547 4326 3599 4378
rect 3611 4326 3663 4378
rect 3675 4326 3727 4378
rect 3739 4326 3791 4378
rect 3803 4326 3855 4378
rect 6144 4326 6196 4378
rect 6208 4326 6260 4378
rect 6272 4326 6324 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 7840 3884 7892 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 2248 3782 2300 3834
rect 2312 3782 2364 3834
rect 2376 3782 2428 3834
rect 2440 3782 2492 3834
rect 2504 3782 2556 3834
rect 4846 3782 4898 3834
rect 4910 3782 4962 3834
rect 4974 3782 5026 3834
rect 5038 3782 5090 3834
rect 5102 3782 5154 3834
rect 7443 3782 7495 3834
rect 7507 3782 7559 3834
rect 7571 3782 7623 3834
rect 7635 3782 7687 3834
rect 7699 3782 7751 3834
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 8208 3476 8260 3528
rect 3547 3238 3599 3290
rect 3611 3238 3663 3290
rect 3675 3238 3727 3290
rect 3739 3238 3791 3290
rect 3803 3238 3855 3290
rect 6144 3238 6196 3290
rect 6208 3238 6260 3290
rect 6272 3238 6324 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 7840 2796 7892 2848
rect 8024 2796 8076 2848
rect 2248 2694 2300 2746
rect 2312 2694 2364 2746
rect 2376 2694 2428 2746
rect 2440 2694 2492 2746
rect 2504 2694 2556 2746
rect 4846 2694 4898 2746
rect 4910 2694 4962 2746
rect 4974 2694 5026 2746
rect 5038 2694 5090 2746
rect 5102 2694 5154 2746
rect 7443 2694 7495 2746
rect 7507 2694 7559 2746
rect 7571 2694 7623 2746
rect 7635 2694 7687 2746
rect 7699 2694 7751 2746
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 3547 2150 3599 2202
rect 3611 2150 3663 2202
rect 3675 2150 3727 2202
rect 3739 2150 3791 2202
rect 3803 2150 3855 2202
rect 6144 2150 6196 2202
rect 6208 2150 6260 2202
rect 6272 2150 6324 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
<< metal2 >>
rect 6642 24712 6698 24721
rect 6642 24647 6698 24656
rect 2248 22332 2556 22352
rect 2248 22330 2254 22332
rect 2310 22330 2334 22332
rect 2390 22330 2414 22332
rect 2470 22330 2494 22332
rect 2550 22330 2556 22332
rect 2310 22278 2312 22330
rect 2492 22278 2494 22330
rect 2248 22276 2254 22278
rect 2310 22276 2334 22278
rect 2390 22276 2414 22278
rect 2470 22276 2494 22278
rect 2550 22276 2556 22278
rect 2248 22256 2556 22276
rect 4846 22332 5154 22352
rect 4846 22330 4852 22332
rect 4908 22330 4932 22332
rect 4988 22330 5012 22332
rect 5068 22330 5092 22332
rect 5148 22330 5154 22332
rect 4908 22278 4910 22330
rect 5090 22278 5092 22330
rect 4846 22276 4852 22278
rect 4908 22276 4932 22278
rect 4988 22276 5012 22278
rect 5068 22276 5092 22278
rect 5148 22276 5154 22278
rect 4846 22256 5154 22276
rect 3547 21788 3855 21808
rect 3547 21786 3553 21788
rect 3609 21786 3633 21788
rect 3689 21786 3713 21788
rect 3769 21786 3793 21788
rect 3849 21786 3855 21788
rect 3609 21734 3611 21786
rect 3791 21734 3793 21786
rect 3547 21732 3553 21734
rect 3609 21732 3633 21734
rect 3689 21732 3713 21734
rect 3769 21732 3793 21734
rect 3849 21732 3855 21734
rect 3547 21712 3855 21732
rect 6144 21788 6452 21808
rect 6144 21786 6150 21788
rect 6206 21786 6230 21788
rect 6286 21786 6310 21788
rect 6366 21786 6390 21788
rect 6446 21786 6452 21788
rect 6206 21734 6208 21786
rect 6388 21734 6390 21786
rect 6144 21732 6150 21734
rect 6206 21732 6230 21734
rect 6286 21732 6310 21734
rect 6366 21732 6390 21734
rect 6446 21732 6452 21734
rect 6144 21712 6452 21732
rect 6656 21554 6684 24647
rect 7838 24168 7894 24177
rect 7838 24103 7894 24112
rect 6734 23624 6790 23633
rect 6734 23559 6790 23568
rect 6748 22166 6776 23559
rect 6826 23080 6882 23089
rect 6826 23015 6882 23024
rect 6840 22234 6868 23015
rect 7443 22332 7751 22352
rect 7443 22330 7449 22332
rect 7505 22330 7529 22332
rect 7585 22330 7609 22332
rect 7665 22330 7689 22332
rect 7745 22330 7751 22332
rect 7505 22278 7507 22330
rect 7687 22278 7689 22330
rect 7443 22276 7449 22278
rect 7505 22276 7529 22278
rect 7585 22276 7609 22278
rect 7665 22276 7689 22278
rect 7745 22276 7751 22278
rect 7443 22256 7751 22276
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 7470 21448 7526 21457
rect 7470 21383 7472 21392
rect 7524 21383 7526 21392
rect 7472 21354 7524 21360
rect 2248 21244 2556 21264
rect 2248 21242 2254 21244
rect 2310 21242 2334 21244
rect 2390 21242 2414 21244
rect 2470 21242 2494 21244
rect 2550 21242 2556 21244
rect 2310 21190 2312 21242
rect 2492 21190 2494 21242
rect 2248 21188 2254 21190
rect 2310 21188 2334 21190
rect 2390 21188 2414 21190
rect 2470 21188 2494 21190
rect 2550 21188 2556 21190
rect 2248 21168 2556 21188
rect 4846 21244 5154 21264
rect 4846 21242 4852 21244
rect 4908 21242 4932 21244
rect 4988 21242 5012 21244
rect 5068 21242 5092 21244
rect 5148 21242 5154 21244
rect 4908 21190 4910 21242
rect 5090 21190 5092 21242
rect 4846 21188 4852 21190
rect 4908 21188 4932 21190
rect 4988 21188 5012 21190
rect 5068 21188 5092 21190
rect 5148 21188 5154 21190
rect 4846 21168 5154 21188
rect 7443 21244 7751 21264
rect 7443 21242 7449 21244
rect 7505 21242 7529 21244
rect 7585 21242 7609 21244
rect 7665 21242 7689 21244
rect 7745 21242 7751 21244
rect 7505 21190 7507 21242
rect 7687 21190 7689 21242
rect 7443 21188 7449 21190
rect 7505 21188 7529 21190
rect 7585 21188 7609 21190
rect 7665 21188 7689 21190
rect 7745 21188 7751 21190
rect 7443 21168 7751 21188
rect 7852 21146 7880 24103
rect 8206 22536 8262 22545
rect 8206 22471 8262 22480
rect 8114 21992 8170 22001
rect 8114 21927 8116 21936
rect 8168 21927 8170 21936
rect 8116 21898 8168 21904
rect 8220 21690 8248 22471
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 8116 20936 8168 20942
rect 8114 20904 8116 20913
rect 8168 20904 8170 20913
rect 8114 20839 8170 20848
rect 3547 20700 3855 20720
rect 3547 20698 3553 20700
rect 3609 20698 3633 20700
rect 3689 20698 3713 20700
rect 3769 20698 3793 20700
rect 3849 20698 3855 20700
rect 3609 20646 3611 20698
rect 3791 20646 3793 20698
rect 3547 20644 3553 20646
rect 3609 20644 3633 20646
rect 3689 20644 3713 20646
rect 3769 20644 3793 20646
rect 3849 20644 3855 20646
rect 3547 20624 3855 20644
rect 6144 20700 6452 20720
rect 6144 20698 6150 20700
rect 6206 20698 6230 20700
rect 6286 20698 6310 20700
rect 6366 20698 6390 20700
rect 6446 20698 6452 20700
rect 6206 20646 6208 20698
rect 6388 20646 6390 20698
rect 6144 20644 6150 20646
rect 6206 20644 6230 20646
rect 6286 20644 6310 20646
rect 6366 20644 6390 20646
rect 6446 20644 6452 20646
rect 6144 20624 6452 20644
rect 8116 20392 8168 20398
rect 8114 20360 8116 20369
rect 8168 20360 8170 20369
rect 8114 20295 8170 20304
rect 2248 20156 2556 20176
rect 2248 20154 2254 20156
rect 2310 20154 2334 20156
rect 2390 20154 2414 20156
rect 2470 20154 2494 20156
rect 2550 20154 2556 20156
rect 2310 20102 2312 20154
rect 2492 20102 2494 20154
rect 2248 20100 2254 20102
rect 2310 20100 2334 20102
rect 2390 20100 2414 20102
rect 2470 20100 2494 20102
rect 2550 20100 2556 20102
rect 2248 20080 2556 20100
rect 4846 20156 5154 20176
rect 4846 20154 4852 20156
rect 4908 20154 4932 20156
rect 4988 20154 5012 20156
rect 5068 20154 5092 20156
rect 5148 20154 5154 20156
rect 4908 20102 4910 20154
rect 5090 20102 5092 20154
rect 4846 20100 4852 20102
rect 4908 20100 4932 20102
rect 4988 20100 5012 20102
rect 5068 20100 5092 20102
rect 5148 20100 5154 20102
rect 4846 20080 5154 20100
rect 7443 20156 7751 20176
rect 7443 20154 7449 20156
rect 7505 20154 7529 20156
rect 7585 20154 7609 20156
rect 7665 20154 7689 20156
rect 7745 20154 7751 20156
rect 7505 20102 7507 20154
rect 7687 20102 7689 20154
rect 7443 20100 7449 20102
rect 7505 20100 7529 20102
rect 7585 20100 7609 20102
rect 7665 20100 7689 20102
rect 7745 20100 7751 20102
rect 7443 20080 7751 20100
rect 8114 19816 8170 19825
rect 8114 19751 8116 19760
rect 8168 19751 8170 19760
rect 8116 19722 8168 19728
rect 3547 19612 3855 19632
rect 3547 19610 3553 19612
rect 3609 19610 3633 19612
rect 3689 19610 3713 19612
rect 3769 19610 3793 19612
rect 3849 19610 3855 19612
rect 3609 19558 3611 19610
rect 3791 19558 3793 19610
rect 3547 19556 3553 19558
rect 3609 19556 3633 19558
rect 3689 19556 3713 19558
rect 3769 19556 3793 19558
rect 3849 19556 3855 19558
rect 3547 19536 3855 19556
rect 6144 19612 6452 19632
rect 6144 19610 6150 19612
rect 6206 19610 6230 19612
rect 6286 19610 6310 19612
rect 6366 19610 6390 19612
rect 6446 19610 6452 19612
rect 6206 19558 6208 19610
rect 6388 19558 6390 19610
rect 6144 19556 6150 19558
rect 6206 19556 6230 19558
rect 6286 19556 6310 19558
rect 6366 19556 6390 19558
rect 6446 19556 6452 19558
rect 6144 19536 6452 19556
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 7470 19272 7526 19281
rect 7470 19207 7472 19216
rect 7524 19207 7526 19216
rect 7472 19178 7524 19184
rect 2248 19068 2556 19088
rect 2248 19066 2254 19068
rect 2310 19066 2334 19068
rect 2390 19066 2414 19068
rect 2470 19066 2494 19068
rect 2550 19066 2556 19068
rect 2310 19014 2312 19066
rect 2492 19014 2494 19066
rect 2248 19012 2254 19014
rect 2310 19012 2334 19014
rect 2390 19012 2414 19014
rect 2470 19012 2494 19014
rect 2550 19012 2556 19014
rect 2248 18992 2556 19012
rect 4846 19068 5154 19088
rect 4846 19066 4852 19068
rect 4908 19066 4932 19068
rect 4988 19066 5012 19068
rect 5068 19066 5092 19068
rect 5148 19066 5154 19068
rect 4908 19014 4910 19066
rect 5090 19014 5092 19066
rect 4846 19012 4852 19014
rect 4908 19012 4932 19014
rect 4988 19012 5012 19014
rect 5068 19012 5092 19014
rect 5148 19012 5154 19014
rect 4846 18992 5154 19012
rect 7443 19068 7751 19088
rect 7443 19066 7449 19068
rect 7505 19066 7529 19068
rect 7585 19066 7609 19068
rect 7665 19066 7689 19068
rect 7745 19066 7751 19068
rect 7505 19014 7507 19066
rect 7687 19014 7689 19066
rect 7443 19012 7449 19014
rect 7505 19012 7529 19014
rect 7585 19012 7609 19014
rect 7665 19012 7689 19014
rect 7745 19012 7751 19014
rect 7443 18992 7751 19012
rect 8128 18873 8156 19314
rect 8114 18864 8170 18873
rect 8114 18799 8170 18808
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 3547 18524 3855 18544
rect 3547 18522 3553 18524
rect 3609 18522 3633 18524
rect 3689 18522 3713 18524
rect 3769 18522 3793 18524
rect 3849 18522 3855 18524
rect 3609 18470 3611 18522
rect 3791 18470 3793 18522
rect 3547 18468 3553 18470
rect 3609 18468 3633 18470
rect 3689 18468 3713 18470
rect 3769 18468 3793 18470
rect 3849 18468 3855 18470
rect 3547 18448 3855 18468
rect 6144 18524 6452 18544
rect 6144 18522 6150 18524
rect 6206 18522 6230 18524
rect 6286 18522 6310 18524
rect 6366 18522 6390 18524
rect 6446 18522 6452 18524
rect 6206 18470 6208 18522
rect 6388 18470 6390 18522
rect 6144 18468 6150 18470
rect 6206 18468 6230 18470
rect 6286 18468 6310 18470
rect 6366 18468 6390 18470
rect 6446 18468 6452 18470
rect 6144 18448 6452 18468
rect 8128 18329 8156 18702
rect 8114 18320 8170 18329
rect 8114 18255 8170 18264
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 2248 17980 2556 18000
rect 2248 17978 2254 17980
rect 2310 17978 2334 17980
rect 2390 17978 2414 17980
rect 2470 17978 2494 17980
rect 2550 17978 2556 17980
rect 2310 17926 2312 17978
rect 2492 17926 2494 17978
rect 2248 17924 2254 17926
rect 2310 17924 2334 17926
rect 2390 17924 2414 17926
rect 2470 17924 2494 17926
rect 2550 17924 2556 17926
rect 2248 17904 2556 17924
rect 4846 17980 5154 18000
rect 4846 17978 4852 17980
rect 4908 17978 4932 17980
rect 4988 17978 5012 17980
rect 5068 17978 5092 17980
rect 5148 17978 5154 17980
rect 4908 17926 4910 17978
rect 5090 17926 5092 17978
rect 4846 17924 4852 17926
rect 4908 17924 4932 17926
rect 4988 17924 5012 17926
rect 5068 17924 5092 17926
rect 5148 17924 5154 17926
rect 4846 17904 5154 17924
rect 7443 17980 7751 18000
rect 7443 17978 7449 17980
rect 7505 17978 7529 17980
rect 7585 17978 7609 17980
rect 7665 17978 7689 17980
rect 7745 17978 7751 17980
rect 7505 17926 7507 17978
rect 7687 17926 7689 17978
rect 7443 17924 7449 17926
rect 7505 17924 7529 17926
rect 7585 17924 7609 17926
rect 7665 17924 7689 17926
rect 7745 17924 7751 17926
rect 7443 17904 7751 17924
rect 8128 17785 8156 18158
rect 8114 17776 8170 17785
rect 8114 17711 8170 17720
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 3547 17436 3855 17456
rect 3547 17434 3553 17436
rect 3609 17434 3633 17436
rect 3689 17434 3713 17436
rect 3769 17434 3793 17436
rect 3849 17434 3855 17436
rect 3609 17382 3611 17434
rect 3791 17382 3793 17434
rect 3547 17380 3553 17382
rect 3609 17380 3633 17382
rect 3689 17380 3713 17382
rect 3769 17380 3793 17382
rect 3849 17380 3855 17382
rect 3547 17360 3855 17380
rect 6144 17436 6452 17456
rect 6144 17434 6150 17436
rect 6206 17434 6230 17436
rect 6286 17434 6310 17436
rect 6366 17434 6390 17436
rect 6446 17434 6452 17436
rect 6206 17382 6208 17434
rect 6388 17382 6390 17434
rect 6144 17380 6150 17382
rect 6206 17380 6230 17382
rect 6286 17380 6310 17382
rect 6366 17380 6390 17382
rect 6446 17380 6452 17382
rect 6144 17360 6452 17380
rect 8128 17241 8156 17614
rect 8114 17232 8170 17241
rect 8114 17167 8170 17176
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 2248 16892 2556 16912
rect 2248 16890 2254 16892
rect 2310 16890 2334 16892
rect 2390 16890 2414 16892
rect 2470 16890 2494 16892
rect 2550 16890 2556 16892
rect 2310 16838 2312 16890
rect 2492 16838 2494 16890
rect 2248 16836 2254 16838
rect 2310 16836 2334 16838
rect 2390 16836 2414 16838
rect 2470 16836 2494 16838
rect 2550 16836 2556 16838
rect 2248 16816 2556 16836
rect 4846 16892 5154 16912
rect 4846 16890 4852 16892
rect 4908 16890 4932 16892
rect 4988 16890 5012 16892
rect 5068 16890 5092 16892
rect 5148 16890 5154 16892
rect 4908 16838 4910 16890
rect 5090 16838 5092 16890
rect 4846 16836 4852 16838
rect 4908 16836 4932 16838
rect 4988 16836 5012 16838
rect 5068 16836 5092 16838
rect 5148 16836 5154 16838
rect 4846 16816 5154 16836
rect 7443 16892 7751 16912
rect 7443 16890 7449 16892
rect 7505 16890 7529 16892
rect 7585 16890 7609 16892
rect 7665 16890 7689 16892
rect 7745 16890 7751 16892
rect 7505 16838 7507 16890
rect 7687 16838 7689 16890
rect 7443 16836 7449 16838
rect 7505 16836 7529 16838
rect 7585 16836 7609 16838
rect 7665 16836 7689 16838
rect 7745 16836 7751 16838
rect 7443 16816 7751 16836
rect 8220 16697 8248 17070
rect 8206 16688 8262 16697
rect 8116 16652 8168 16658
rect 8206 16623 8262 16632
rect 8116 16594 8168 16600
rect 3547 16348 3855 16368
rect 3547 16346 3553 16348
rect 3609 16346 3633 16348
rect 3689 16346 3713 16348
rect 3769 16346 3793 16348
rect 3849 16346 3855 16348
rect 3609 16294 3611 16346
rect 3791 16294 3793 16346
rect 3547 16292 3553 16294
rect 3609 16292 3633 16294
rect 3689 16292 3713 16294
rect 3769 16292 3793 16294
rect 3849 16292 3855 16294
rect 3547 16272 3855 16292
rect 6144 16348 6452 16368
rect 6144 16346 6150 16348
rect 6206 16346 6230 16348
rect 6286 16346 6310 16348
rect 6366 16346 6390 16348
rect 6446 16346 6452 16348
rect 6206 16294 6208 16346
rect 6388 16294 6390 16346
rect 6144 16292 6150 16294
rect 6206 16292 6230 16294
rect 6286 16292 6310 16294
rect 6366 16292 6390 16294
rect 6446 16292 6452 16294
rect 6144 16272 6452 16292
rect 8128 16153 8156 16594
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 2248 15804 2556 15824
rect 2248 15802 2254 15804
rect 2310 15802 2334 15804
rect 2390 15802 2414 15804
rect 2470 15802 2494 15804
rect 2550 15802 2556 15804
rect 2310 15750 2312 15802
rect 2492 15750 2494 15802
rect 2248 15748 2254 15750
rect 2310 15748 2334 15750
rect 2390 15748 2414 15750
rect 2470 15748 2494 15750
rect 2550 15748 2556 15750
rect 2248 15728 2556 15748
rect 4846 15804 5154 15824
rect 4846 15802 4852 15804
rect 4908 15802 4932 15804
rect 4988 15802 5012 15804
rect 5068 15802 5092 15804
rect 5148 15802 5154 15804
rect 4908 15750 4910 15802
rect 5090 15750 5092 15802
rect 4846 15748 4852 15750
rect 4908 15748 4932 15750
rect 4988 15748 5012 15750
rect 5068 15748 5092 15750
rect 5148 15748 5154 15750
rect 4846 15728 5154 15748
rect 7443 15804 7751 15824
rect 7443 15802 7449 15804
rect 7505 15802 7529 15804
rect 7585 15802 7609 15804
rect 7665 15802 7689 15804
rect 7745 15802 7751 15804
rect 7505 15750 7507 15802
rect 7687 15750 7689 15802
rect 7443 15748 7449 15750
rect 7505 15748 7529 15750
rect 7585 15748 7609 15750
rect 7665 15748 7689 15750
rect 7745 15748 7751 15750
rect 7443 15728 7751 15748
rect 8128 15609 8156 15982
rect 8114 15600 8170 15609
rect 8114 15535 8170 15544
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 3547 15260 3855 15280
rect 3547 15258 3553 15260
rect 3609 15258 3633 15260
rect 3689 15258 3713 15260
rect 3769 15258 3793 15260
rect 3849 15258 3855 15260
rect 3609 15206 3611 15258
rect 3791 15206 3793 15258
rect 3547 15204 3553 15206
rect 3609 15204 3633 15206
rect 3689 15204 3713 15206
rect 3769 15204 3793 15206
rect 3849 15204 3855 15206
rect 3547 15184 3855 15204
rect 6144 15260 6452 15280
rect 6144 15258 6150 15260
rect 6206 15258 6230 15260
rect 6286 15258 6310 15260
rect 6366 15258 6390 15260
rect 6446 15258 6452 15260
rect 6206 15206 6208 15258
rect 6388 15206 6390 15258
rect 6144 15204 6150 15206
rect 6206 15204 6230 15206
rect 6286 15204 6310 15206
rect 6366 15204 6390 15206
rect 6446 15204 6452 15206
rect 6144 15184 6452 15204
rect 8128 15065 8156 15438
rect 8114 15056 8170 15065
rect 8114 14991 8170 15000
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 2248 14716 2556 14736
rect 2248 14714 2254 14716
rect 2310 14714 2334 14716
rect 2390 14714 2414 14716
rect 2470 14714 2494 14716
rect 2550 14714 2556 14716
rect 2310 14662 2312 14714
rect 2492 14662 2494 14714
rect 2248 14660 2254 14662
rect 2310 14660 2334 14662
rect 2390 14660 2414 14662
rect 2470 14660 2494 14662
rect 2550 14660 2556 14662
rect 2248 14640 2556 14660
rect 4846 14716 5154 14736
rect 4846 14714 4852 14716
rect 4908 14714 4932 14716
rect 4988 14714 5012 14716
rect 5068 14714 5092 14716
rect 5148 14714 5154 14716
rect 4908 14662 4910 14714
rect 5090 14662 5092 14714
rect 4846 14660 4852 14662
rect 4908 14660 4932 14662
rect 4988 14660 5012 14662
rect 5068 14660 5092 14662
rect 5148 14660 5154 14662
rect 4846 14640 5154 14660
rect 7443 14716 7751 14736
rect 7443 14714 7449 14716
rect 7505 14714 7529 14716
rect 7585 14714 7609 14716
rect 7665 14714 7689 14716
rect 7745 14714 7751 14716
rect 7505 14662 7507 14714
rect 7687 14662 7689 14714
rect 7443 14660 7449 14662
rect 7505 14660 7529 14662
rect 7585 14660 7609 14662
rect 7665 14660 7689 14662
rect 7745 14660 7751 14662
rect 7443 14640 7751 14660
rect 8128 14521 8156 14894
rect 8114 14512 8170 14521
rect 8114 14447 8170 14456
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 3547 14172 3855 14192
rect 3547 14170 3553 14172
rect 3609 14170 3633 14172
rect 3689 14170 3713 14172
rect 3769 14170 3793 14172
rect 3849 14170 3855 14172
rect 3609 14118 3611 14170
rect 3791 14118 3793 14170
rect 3547 14116 3553 14118
rect 3609 14116 3633 14118
rect 3689 14116 3713 14118
rect 3769 14116 3793 14118
rect 3849 14116 3855 14118
rect 3547 14096 3855 14116
rect 6144 14172 6452 14192
rect 6144 14170 6150 14172
rect 6206 14170 6230 14172
rect 6286 14170 6310 14172
rect 6366 14170 6390 14172
rect 6446 14170 6452 14172
rect 6206 14118 6208 14170
rect 6388 14118 6390 14170
rect 6144 14116 6150 14118
rect 6206 14116 6230 14118
rect 6286 14116 6310 14118
rect 6366 14116 6390 14118
rect 6446 14116 6452 14118
rect 6144 14096 6452 14116
rect 8128 13977 8156 14350
rect 8114 13968 8170 13977
rect 8114 13903 8170 13912
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 2248 13628 2556 13648
rect 2248 13626 2254 13628
rect 2310 13626 2334 13628
rect 2390 13626 2414 13628
rect 2470 13626 2494 13628
rect 2550 13626 2556 13628
rect 2310 13574 2312 13626
rect 2492 13574 2494 13626
rect 2248 13572 2254 13574
rect 2310 13572 2334 13574
rect 2390 13572 2414 13574
rect 2470 13572 2494 13574
rect 2550 13572 2556 13574
rect 2248 13552 2556 13572
rect 4846 13628 5154 13648
rect 4846 13626 4852 13628
rect 4908 13626 4932 13628
rect 4988 13626 5012 13628
rect 5068 13626 5092 13628
rect 5148 13626 5154 13628
rect 4908 13574 4910 13626
rect 5090 13574 5092 13626
rect 4846 13572 4852 13574
rect 4908 13572 4932 13574
rect 4988 13572 5012 13574
rect 5068 13572 5092 13574
rect 5148 13572 5154 13574
rect 4846 13552 5154 13572
rect 7443 13628 7751 13648
rect 7443 13626 7449 13628
rect 7505 13626 7529 13628
rect 7585 13626 7609 13628
rect 7665 13626 7689 13628
rect 7745 13626 7751 13628
rect 7505 13574 7507 13626
rect 7687 13574 7689 13626
rect 7443 13572 7449 13574
rect 7505 13572 7529 13574
rect 7585 13572 7609 13574
rect 7665 13572 7689 13574
rect 7745 13572 7751 13574
rect 7443 13552 7751 13572
rect 8128 13433 8156 13806
rect 8114 13424 8170 13433
rect 8114 13359 8170 13368
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 3547 13084 3855 13104
rect 3547 13082 3553 13084
rect 3609 13082 3633 13084
rect 3689 13082 3713 13084
rect 3769 13082 3793 13084
rect 3849 13082 3855 13084
rect 3609 13030 3611 13082
rect 3791 13030 3793 13082
rect 3547 13028 3553 13030
rect 3609 13028 3633 13030
rect 3689 13028 3713 13030
rect 3769 13028 3793 13030
rect 3849 13028 3855 13030
rect 3547 13008 3855 13028
rect 6144 13084 6452 13104
rect 6144 13082 6150 13084
rect 6206 13082 6230 13084
rect 6286 13082 6310 13084
rect 6366 13082 6390 13084
rect 6446 13082 6452 13084
rect 6206 13030 6208 13082
rect 6388 13030 6390 13082
rect 6144 13028 6150 13030
rect 6206 13028 6230 13030
rect 6286 13028 6310 13030
rect 6366 13028 6390 13030
rect 6446 13028 6452 13030
rect 6144 13008 6452 13028
rect 8128 12889 8156 13262
rect 8114 12880 8170 12889
rect 8114 12815 8170 12824
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 2248 12540 2556 12560
rect 2248 12538 2254 12540
rect 2310 12538 2334 12540
rect 2390 12538 2414 12540
rect 2470 12538 2494 12540
rect 2550 12538 2556 12540
rect 2310 12486 2312 12538
rect 2492 12486 2494 12538
rect 2248 12484 2254 12486
rect 2310 12484 2334 12486
rect 2390 12484 2414 12486
rect 2470 12484 2494 12486
rect 2550 12484 2556 12486
rect 2248 12464 2556 12484
rect 4846 12540 5154 12560
rect 4846 12538 4852 12540
rect 4908 12538 4932 12540
rect 4988 12538 5012 12540
rect 5068 12538 5092 12540
rect 5148 12538 5154 12540
rect 4908 12486 4910 12538
rect 5090 12486 5092 12538
rect 4846 12484 4852 12486
rect 4908 12484 4932 12486
rect 4988 12484 5012 12486
rect 5068 12484 5092 12486
rect 5148 12484 5154 12486
rect 4846 12464 5154 12484
rect 7443 12540 7751 12560
rect 7443 12538 7449 12540
rect 7505 12538 7529 12540
rect 7585 12538 7609 12540
rect 7665 12538 7689 12540
rect 7745 12538 7751 12540
rect 7505 12486 7507 12538
rect 7687 12486 7689 12538
rect 7443 12484 7449 12486
rect 7505 12484 7529 12486
rect 7585 12484 7609 12486
rect 7665 12484 7689 12486
rect 7745 12484 7751 12486
rect 7443 12464 7751 12484
rect 8128 12481 8156 12582
rect 8114 12472 8170 12481
rect 8114 12407 8170 12416
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 3547 11996 3855 12016
rect 3547 11994 3553 11996
rect 3609 11994 3633 11996
rect 3689 11994 3713 11996
rect 3769 11994 3793 11996
rect 3849 11994 3855 11996
rect 3609 11942 3611 11994
rect 3791 11942 3793 11994
rect 3547 11940 3553 11942
rect 3609 11940 3633 11942
rect 3689 11940 3713 11942
rect 3769 11940 3793 11942
rect 3849 11940 3855 11942
rect 3547 11920 3855 11940
rect 6144 11996 6452 12016
rect 6144 11994 6150 11996
rect 6206 11994 6230 11996
rect 6286 11994 6310 11996
rect 6366 11994 6390 11996
rect 6446 11994 6452 11996
rect 6206 11942 6208 11994
rect 6388 11942 6390 11994
rect 6144 11940 6150 11942
rect 6206 11940 6230 11942
rect 6286 11940 6310 11942
rect 6366 11940 6390 11942
rect 6446 11940 6452 11942
rect 6144 11920 6452 11940
rect 8128 11937 8156 12174
rect 8114 11928 8170 11937
rect 8114 11863 8170 11872
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 2248 11452 2556 11472
rect 2248 11450 2254 11452
rect 2310 11450 2334 11452
rect 2390 11450 2414 11452
rect 2470 11450 2494 11452
rect 2550 11450 2556 11452
rect 2310 11398 2312 11450
rect 2492 11398 2494 11450
rect 2248 11396 2254 11398
rect 2310 11396 2334 11398
rect 2390 11396 2414 11398
rect 2470 11396 2494 11398
rect 2550 11396 2556 11398
rect 2248 11376 2556 11396
rect 4846 11452 5154 11472
rect 4846 11450 4852 11452
rect 4908 11450 4932 11452
rect 4988 11450 5012 11452
rect 5068 11450 5092 11452
rect 5148 11450 5154 11452
rect 4908 11398 4910 11450
rect 5090 11398 5092 11450
rect 4846 11396 4852 11398
rect 4908 11396 4932 11398
rect 4988 11396 5012 11398
rect 5068 11396 5092 11398
rect 5148 11396 5154 11398
rect 4846 11376 5154 11396
rect 7443 11452 7751 11472
rect 7443 11450 7449 11452
rect 7505 11450 7529 11452
rect 7585 11450 7609 11452
rect 7665 11450 7689 11452
rect 7745 11450 7751 11452
rect 7505 11398 7507 11450
rect 7687 11398 7689 11450
rect 7443 11396 7449 11398
rect 7505 11396 7529 11398
rect 7585 11396 7609 11398
rect 7665 11396 7689 11398
rect 7745 11396 7751 11398
rect 7443 11376 7751 11396
rect 8128 11393 8156 11494
rect 8114 11384 8170 11393
rect 8114 11319 8170 11328
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 3547 10908 3855 10928
rect 3547 10906 3553 10908
rect 3609 10906 3633 10908
rect 3689 10906 3713 10908
rect 3769 10906 3793 10908
rect 3849 10906 3855 10908
rect 3609 10854 3611 10906
rect 3791 10854 3793 10906
rect 3547 10852 3553 10854
rect 3609 10852 3633 10854
rect 3689 10852 3713 10854
rect 3769 10852 3793 10854
rect 3849 10852 3855 10854
rect 3547 10832 3855 10852
rect 6144 10908 6452 10928
rect 6144 10906 6150 10908
rect 6206 10906 6230 10908
rect 6286 10906 6310 10908
rect 6366 10906 6390 10908
rect 6446 10906 6452 10908
rect 6206 10854 6208 10906
rect 6388 10854 6390 10906
rect 6144 10852 6150 10854
rect 6206 10852 6230 10854
rect 6286 10852 6310 10854
rect 6366 10852 6390 10854
rect 6446 10852 6452 10854
rect 6144 10832 6452 10852
rect 8128 10849 8156 11086
rect 8114 10840 8170 10849
rect 8114 10775 8170 10784
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 2248 10364 2556 10384
rect 2248 10362 2254 10364
rect 2310 10362 2334 10364
rect 2390 10362 2414 10364
rect 2470 10362 2494 10364
rect 2550 10362 2556 10364
rect 2310 10310 2312 10362
rect 2492 10310 2494 10362
rect 2248 10308 2254 10310
rect 2310 10308 2334 10310
rect 2390 10308 2414 10310
rect 2470 10308 2494 10310
rect 2550 10308 2556 10310
rect 2248 10288 2556 10308
rect 4846 10364 5154 10384
rect 4846 10362 4852 10364
rect 4908 10362 4932 10364
rect 4988 10362 5012 10364
rect 5068 10362 5092 10364
rect 5148 10362 5154 10364
rect 4908 10310 4910 10362
rect 5090 10310 5092 10362
rect 4846 10308 4852 10310
rect 4908 10308 4932 10310
rect 4988 10308 5012 10310
rect 5068 10308 5092 10310
rect 5148 10308 5154 10310
rect 4846 10288 5154 10308
rect 7443 10364 7751 10384
rect 7443 10362 7449 10364
rect 7505 10362 7529 10364
rect 7585 10362 7609 10364
rect 7665 10362 7689 10364
rect 7745 10362 7751 10364
rect 7505 10310 7507 10362
rect 7687 10310 7689 10362
rect 7443 10308 7449 10310
rect 7505 10308 7529 10310
rect 7585 10308 7609 10310
rect 7665 10308 7689 10310
rect 7745 10308 7751 10310
rect 7443 10288 7751 10308
rect 8128 10305 8156 10406
rect 8114 10296 8170 10305
rect 8114 10231 8170 10240
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 3547 9820 3855 9840
rect 3547 9818 3553 9820
rect 3609 9818 3633 9820
rect 3689 9818 3713 9820
rect 3769 9818 3793 9820
rect 3849 9818 3855 9820
rect 3609 9766 3611 9818
rect 3791 9766 3793 9818
rect 3547 9764 3553 9766
rect 3609 9764 3633 9766
rect 3689 9764 3713 9766
rect 3769 9764 3793 9766
rect 3849 9764 3855 9766
rect 3547 9744 3855 9764
rect 6144 9820 6452 9840
rect 6144 9818 6150 9820
rect 6206 9818 6230 9820
rect 6286 9818 6310 9820
rect 6366 9818 6390 9820
rect 6446 9818 6452 9820
rect 6206 9766 6208 9818
rect 6388 9766 6390 9818
rect 6144 9764 6150 9766
rect 6206 9764 6230 9766
rect 6286 9764 6310 9766
rect 6366 9764 6390 9766
rect 6446 9764 6452 9766
rect 6144 9744 6452 9764
rect 8128 9761 8156 9998
rect 8114 9752 8170 9761
rect 8114 9687 8170 9696
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 2248 9276 2556 9296
rect 2248 9274 2254 9276
rect 2310 9274 2334 9276
rect 2390 9274 2414 9276
rect 2470 9274 2494 9276
rect 2550 9274 2556 9276
rect 2310 9222 2312 9274
rect 2492 9222 2494 9274
rect 2248 9220 2254 9222
rect 2310 9220 2334 9222
rect 2390 9220 2414 9222
rect 2470 9220 2494 9222
rect 2550 9220 2556 9222
rect 2248 9200 2556 9220
rect 4846 9276 5154 9296
rect 4846 9274 4852 9276
rect 4908 9274 4932 9276
rect 4988 9274 5012 9276
rect 5068 9274 5092 9276
rect 5148 9274 5154 9276
rect 4908 9222 4910 9274
rect 5090 9222 5092 9274
rect 4846 9220 4852 9222
rect 4908 9220 4932 9222
rect 4988 9220 5012 9222
rect 5068 9220 5092 9222
rect 5148 9220 5154 9222
rect 4846 9200 5154 9220
rect 7443 9276 7751 9296
rect 7443 9274 7449 9276
rect 7505 9274 7529 9276
rect 7585 9274 7609 9276
rect 7665 9274 7689 9276
rect 7745 9274 7751 9276
rect 7505 9222 7507 9274
rect 7687 9222 7689 9274
rect 7443 9220 7449 9222
rect 7505 9220 7529 9222
rect 7585 9220 7609 9222
rect 7665 9220 7689 9222
rect 7745 9220 7751 9222
rect 7443 9200 7751 9220
rect 8128 9217 8156 9318
rect 8114 9208 8170 9217
rect 8114 9143 8170 9152
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 3547 8732 3855 8752
rect 3547 8730 3553 8732
rect 3609 8730 3633 8732
rect 3689 8730 3713 8732
rect 3769 8730 3793 8732
rect 3849 8730 3855 8732
rect 3609 8678 3611 8730
rect 3791 8678 3793 8730
rect 3547 8676 3553 8678
rect 3609 8676 3633 8678
rect 3689 8676 3713 8678
rect 3769 8676 3793 8678
rect 3849 8676 3855 8678
rect 3547 8656 3855 8676
rect 6144 8732 6452 8752
rect 6144 8730 6150 8732
rect 6206 8730 6230 8732
rect 6286 8730 6310 8732
rect 6366 8730 6390 8732
rect 6446 8730 6452 8732
rect 6206 8678 6208 8730
rect 6388 8678 6390 8730
rect 6144 8676 6150 8678
rect 6206 8676 6230 8678
rect 6286 8676 6310 8678
rect 6366 8676 6390 8678
rect 6446 8676 6452 8678
rect 6144 8656 6452 8676
rect 8128 8673 8156 8910
rect 8114 8664 8170 8673
rect 8114 8599 8170 8608
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 2248 8188 2556 8208
rect 2248 8186 2254 8188
rect 2310 8186 2334 8188
rect 2390 8186 2414 8188
rect 2470 8186 2494 8188
rect 2550 8186 2556 8188
rect 2310 8134 2312 8186
rect 2492 8134 2494 8186
rect 2248 8132 2254 8134
rect 2310 8132 2334 8134
rect 2390 8132 2414 8134
rect 2470 8132 2494 8134
rect 2550 8132 2556 8134
rect 2248 8112 2556 8132
rect 4846 8188 5154 8208
rect 4846 8186 4852 8188
rect 4908 8186 4932 8188
rect 4988 8186 5012 8188
rect 5068 8186 5092 8188
rect 5148 8186 5154 8188
rect 4908 8134 4910 8186
rect 5090 8134 5092 8186
rect 4846 8132 4852 8134
rect 4908 8132 4932 8134
rect 4988 8132 5012 8134
rect 5068 8132 5092 8134
rect 5148 8132 5154 8134
rect 4846 8112 5154 8132
rect 7443 8188 7751 8208
rect 7443 8186 7449 8188
rect 7505 8186 7529 8188
rect 7585 8186 7609 8188
rect 7665 8186 7689 8188
rect 7745 8186 7751 8188
rect 7505 8134 7507 8186
rect 7687 8134 7689 8186
rect 7443 8132 7449 8134
rect 7505 8132 7529 8134
rect 7585 8132 7609 8134
rect 7665 8132 7689 8134
rect 7745 8132 7751 8134
rect 7443 8112 7751 8132
rect 8128 8129 8156 8298
rect 8114 8120 8170 8129
rect 8114 8055 8170 8064
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 3547 7644 3855 7664
rect 3547 7642 3553 7644
rect 3609 7642 3633 7644
rect 3689 7642 3713 7644
rect 3769 7642 3793 7644
rect 3849 7642 3855 7644
rect 3609 7590 3611 7642
rect 3791 7590 3793 7642
rect 3547 7588 3553 7590
rect 3609 7588 3633 7590
rect 3689 7588 3713 7590
rect 3769 7588 3793 7590
rect 3849 7588 3855 7590
rect 3547 7568 3855 7588
rect 6144 7644 6452 7664
rect 6144 7642 6150 7644
rect 6206 7642 6230 7644
rect 6286 7642 6310 7644
rect 6366 7642 6390 7644
rect 6446 7642 6452 7644
rect 6206 7590 6208 7642
rect 6388 7590 6390 7642
rect 6144 7588 6150 7590
rect 6206 7588 6230 7590
rect 6286 7588 6310 7590
rect 6366 7588 6390 7590
rect 6446 7588 6452 7590
rect 6144 7568 6452 7588
rect 8128 7585 8156 7822
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 2248 7100 2556 7120
rect 2248 7098 2254 7100
rect 2310 7098 2334 7100
rect 2390 7098 2414 7100
rect 2470 7098 2494 7100
rect 2550 7098 2556 7100
rect 2310 7046 2312 7098
rect 2492 7046 2494 7098
rect 2248 7044 2254 7046
rect 2310 7044 2334 7046
rect 2390 7044 2414 7046
rect 2470 7044 2494 7046
rect 2550 7044 2556 7046
rect 2248 7024 2556 7044
rect 4846 7100 5154 7120
rect 4846 7098 4852 7100
rect 4908 7098 4932 7100
rect 4988 7098 5012 7100
rect 5068 7098 5092 7100
rect 5148 7098 5154 7100
rect 4908 7046 4910 7098
rect 5090 7046 5092 7098
rect 4846 7044 4852 7046
rect 4908 7044 4932 7046
rect 4988 7044 5012 7046
rect 5068 7044 5092 7046
rect 5148 7044 5154 7046
rect 4846 7024 5154 7044
rect 7443 7100 7751 7120
rect 7443 7098 7449 7100
rect 7505 7098 7529 7100
rect 7585 7098 7609 7100
rect 7665 7098 7689 7100
rect 7745 7098 7751 7100
rect 7505 7046 7507 7098
rect 7687 7046 7689 7098
rect 7443 7044 7449 7046
rect 7505 7044 7529 7046
rect 7585 7044 7609 7046
rect 7665 7044 7689 7046
rect 7745 7044 7751 7046
rect 7443 7024 7751 7044
rect 8128 7041 8156 7142
rect 8114 7032 8170 7041
rect 8114 6967 8170 6976
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 3547 6556 3855 6576
rect 3547 6554 3553 6556
rect 3609 6554 3633 6556
rect 3689 6554 3713 6556
rect 3769 6554 3793 6556
rect 3849 6554 3855 6556
rect 3609 6502 3611 6554
rect 3791 6502 3793 6554
rect 3547 6500 3553 6502
rect 3609 6500 3633 6502
rect 3689 6500 3713 6502
rect 3769 6500 3793 6502
rect 3849 6500 3855 6502
rect 3547 6480 3855 6500
rect 6144 6556 6452 6576
rect 6144 6554 6150 6556
rect 6206 6554 6230 6556
rect 6286 6554 6310 6556
rect 6366 6554 6390 6556
rect 6446 6554 6452 6556
rect 6206 6502 6208 6554
rect 6388 6502 6390 6554
rect 6144 6500 6150 6502
rect 6206 6500 6230 6502
rect 6286 6500 6310 6502
rect 6366 6500 6390 6502
rect 6446 6500 6452 6502
rect 6144 6480 6452 6500
rect 8128 6497 8156 6734
rect 8114 6488 8170 6497
rect 8114 6423 8170 6432
rect 8116 6112 8168 6118
rect 8114 6080 8116 6089
rect 8168 6080 8170 6089
rect 2248 6012 2556 6032
rect 2248 6010 2254 6012
rect 2310 6010 2334 6012
rect 2390 6010 2414 6012
rect 2470 6010 2494 6012
rect 2550 6010 2556 6012
rect 2310 5958 2312 6010
rect 2492 5958 2494 6010
rect 2248 5956 2254 5958
rect 2310 5956 2334 5958
rect 2390 5956 2414 5958
rect 2470 5956 2494 5958
rect 2550 5956 2556 5958
rect 2248 5936 2556 5956
rect 4846 6012 5154 6032
rect 4846 6010 4852 6012
rect 4908 6010 4932 6012
rect 4988 6010 5012 6012
rect 5068 6010 5092 6012
rect 5148 6010 5154 6012
rect 4908 5958 4910 6010
rect 5090 5958 5092 6010
rect 4846 5956 4852 5958
rect 4908 5956 4932 5958
rect 4988 5956 5012 5958
rect 5068 5956 5092 5958
rect 5148 5956 5154 5958
rect 4846 5936 5154 5956
rect 7443 6012 7751 6032
rect 8114 6015 8170 6024
rect 7443 6010 7449 6012
rect 7505 6010 7529 6012
rect 7585 6010 7609 6012
rect 7665 6010 7689 6012
rect 7745 6010 7751 6012
rect 7505 5958 7507 6010
rect 7687 5958 7689 6010
rect 7443 5956 7449 5958
rect 7505 5956 7529 5958
rect 7585 5956 7609 5958
rect 7665 5956 7689 5958
rect 7745 5956 7751 5958
rect 7443 5936 7751 5956
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5545 8156 5646
rect 8114 5536 8170 5545
rect 3547 5468 3855 5488
rect 3547 5466 3553 5468
rect 3609 5466 3633 5468
rect 3689 5466 3713 5468
rect 3769 5466 3793 5468
rect 3849 5466 3855 5468
rect 3609 5414 3611 5466
rect 3791 5414 3793 5466
rect 3547 5412 3553 5414
rect 3609 5412 3633 5414
rect 3689 5412 3713 5414
rect 3769 5412 3793 5414
rect 3849 5412 3855 5414
rect 3547 5392 3855 5412
rect 6144 5468 6452 5488
rect 8114 5471 8170 5480
rect 6144 5466 6150 5468
rect 6206 5466 6230 5468
rect 6286 5466 6310 5468
rect 6366 5466 6390 5468
rect 6446 5466 6452 5468
rect 6206 5414 6208 5466
rect 6388 5414 6390 5466
rect 6144 5412 6150 5414
rect 6206 5412 6230 5414
rect 6286 5412 6310 5414
rect 6366 5412 6390 5414
rect 6446 5412 6452 5414
rect 6144 5392 6452 5412
rect 8116 5024 8168 5030
rect 8114 4992 8116 5001
rect 8168 4992 8170 5001
rect 2248 4924 2556 4944
rect 2248 4922 2254 4924
rect 2310 4922 2334 4924
rect 2390 4922 2414 4924
rect 2470 4922 2494 4924
rect 2550 4922 2556 4924
rect 2310 4870 2312 4922
rect 2492 4870 2494 4922
rect 2248 4868 2254 4870
rect 2310 4868 2334 4870
rect 2390 4868 2414 4870
rect 2470 4868 2494 4870
rect 2550 4868 2556 4870
rect 2248 4848 2556 4868
rect 4846 4924 5154 4944
rect 4846 4922 4852 4924
rect 4908 4922 4932 4924
rect 4988 4922 5012 4924
rect 5068 4922 5092 4924
rect 5148 4922 5154 4924
rect 4908 4870 4910 4922
rect 5090 4870 5092 4922
rect 4846 4868 4852 4870
rect 4908 4868 4932 4870
rect 4988 4868 5012 4870
rect 5068 4868 5092 4870
rect 5148 4868 5154 4870
rect 4846 4848 5154 4868
rect 7443 4924 7751 4944
rect 8114 4927 8170 4936
rect 7443 4922 7449 4924
rect 7505 4922 7529 4924
rect 7585 4922 7609 4924
rect 7665 4922 7689 4924
rect 7745 4922 7751 4924
rect 7505 4870 7507 4922
rect 7687 4870 7689 4922
rect 7443 4868 7449 4870
rect 7505 4868 7529 4870
rect 7585 4868 7609 4870
rect 7665 4868 7689 4870
rect 7745 4868 7751 4870
rect 7443 4848 7751 4868
rect 8116 4480 8168 4486
rect 8114 4448 8116 4457
rect 8168 4448 8170 4457
rect 3547 4380 3855 4400
rect 3547 4378 3553 4380
rect 3609 4378 3633 4380
rect 3689 4378 3713 4380
rect 3769 4378 3793 4380
rect 3849 4378 3855 4380
rect 3609 4326 3611 4378
rect 3791 4326 3793 4378
rect 3547 4324 3553 4326
rect 3609 4324 3633 4326
rect 3689 4324 3713 4326
rect 3769 4324 3793 4326
rect 3849 4324 3855 4326
rect 3547 4304 3855 4324
rect 6144 4380 6452 4400
rect 8114 4383 8170 4392
rect 6144 4378 6150 4380
rect 6206 4378 6230 4380
rect 6286 4378 6310 4380
rect 6366 4378 6390 4380
rect 6446 4378 6452 4380
rect 6206 4326 6208 4378
rect 6388 4326 6390 4378
rect 6144 4324 6150 4326
rect 6206 4324 6230 4326
rect 6286 4324 6310 4326
rect 6366 4324 6390 4326
rect 6446 4324 6452 4326
rect 6144 4304 6452 4324
rect 7840 3936 7892 3942
rect 7838 3904 7840 3913
rect 8116 3936 8168 3942
rect 7892 3904 7894 3913
rect 2248 3836 2556 3856
rect 2248 3834 2254 3836
rect 2310 3834 2334 3836
rect 2390 3834 2414 3836
rect 2470 3834 2494 3836
rect 2550 3834 2556 3836
rect 2310 3782 2312 3834
rect 2492 3782 2494 3834
rect 2248 3780 2254 3782
rect 2310 3780 2334 3782
rect 2390 3780 2414 3782
rect 2470 3780 2494 3782
rect 2550 3780 2556 3782
rect 2248 3760 2556 3780
rect 4846 3836 5154 3856
rect 4846 3834 4852 3836
rect 4908 3834 4932 3836
rect 4988 3834 5012 3836
rect 5068 3834 5092 3836
rect 5148 3834 5154 3836
rect 4908 3782 4910 3834
rect 5090 3782 5092 3834
rect 4846 3780 4852 3782
rect 4908 3780 4932 3782
rect 4988 3780 5012 3782
rect 5068 3780 5092 3782
rect 5148 3780 5154 3782
rect 4846 3760 5154 3780
rect 7443 3836 7751 3856
rect 8116 3878 8168 3884
rect 7838 3839 7894 3848
rect 7443 3834 7449 3836
rect 7505 3834 7529 3836
rect 7585 3834 7609 3836
rect 7665 3834 7689 3836
rect 7745 3834 7751 3836
rect 7505 3782 7507 3834
rect 7687 3782 7689 3834
rect 7443 3780 7449 3782
rect 7505 3780 7529 3782
rect 7585 3780 7609 3782
rect 7665 3780 7689 3782
rect 7745 3780 7751 3782
rect 7443 3760 7751 3780
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3369 7512 3470
rect 7470 3360 7526 3369
rect 3547 3292 3855 3312
rect 3547 3290 3553 3292
rect 3609 3290 3633 3292
rect 3689 3290 3713 3292
rect 3769 3290 3793 3292
rect 3849 3290 3855 3292
rect 3609 3238 3611 3290
rect 3791 3238 3793 3290
rect 3547 3236 3553 3238
rect 3609 3236 3633 3238
rect 3689 3236 3713 3238
rect 3769 3236 3793 3238
rect 3849 3236 3855 3238
rect 3547 3216 3855 3236
rect 6144 3292 6452 3312
rect 7470 3295 7526 3304
rect 6144 3290 6150 3292
rect 6206 3290 6230 3292
rect 6286 3290 6310 3292
rect 6366 3290 6390 3292
rect 6446 3290 6452 3292
rect 6206 3238 6208 3290
rect 6388 3238 6390 3290
rect 6144 3236 6150 3238
rect 6206 3236 6230 3238
rect 6286 3236 6310 3238
rect 6366 3236 6390 3238
rect 6446 3236 6452 3238
rect 6144 3216 6452 3236
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 8024 2848 8076 2854
rect 8128 2825 8156 3878
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8024 2790 8076 2796
rect 8114 2816 8170 2825
rect 2248 2748 2556 2768
rect 2248 2746 2254 2748
rect 2310 2746 2334 2748
rect 2390 2746 2414 2748
rect 2470 2746 2494 2748
rect 2550 2746 2556 2748
rect 2310 2694 2312 2746
rect 2492 2694 2494 2746
rect 2248 2692 2254 2694
rect 2310 2692 2334 2694
rect 2390 2692 2414 2694
rect 2470 2692 2494 2694
rect 2550 2692 2556 2694
rect 2248 2672 2556 2692
rect 4846 2748 5154 2768
rect 4846 2746 4852 2748
rect 4908 2746 4932 2748
rect 4988 2746 5012 2748
rect 5068 2746 5092 2748
rect 5148 2746 5154 2748
rect 4908 2694 4910 2746
rect 5090 2694 5092 2746
rect 4846 2692 4852 2694
rect 4908 2692 4932 2694
rect 4988 2692 5012 2694
rect 5068 2692 5092 2694
rect 5148 2692 5154 2694
rect 4846 2672 5154 2692
rect 7443 2748 7751 2768
rect 7443 2746 7449 2748
rect 7505 2746 7529 2748
rect 7585 2746 7609 2748
rect 7665 2746 7689 2748
rect 7745 2746 7751 2748
rect 7505 2694 7507 2746
rect 7687 2694 7689 2746
rect 7443 2692 7449 2694
rect 7505 2692 7529 2694
rect 7585 2692 7609 2694
rect 7665 2692 7689 2694
rect 7745 2692 7751 2694
rect 7443 2672 7751 2692
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 3547 2204 3855 2224
rect 3547 2202 3553 2204
rect 3609 2202 3633 2204
rect 3689 2202 3713 2204
rect 3769 2202 3793 2204
rect 3849 2202 3855 2204
rect 3609 2150 3611 2202
rect 3791 2150 3793 2202
rect 3547 2148 3553 2150
rect 3609 2148 3633 2150
rect 3689 2148 3713 2150
rect 3769 2148 3793 2150
rect 3849 2148 3855 2150
rect 3547 2128 3855 2148
rect 6144 2204 6452 2224
rect 6144 2202 6150 2204
rect 6206 2202 6230 2204
rect 6286 2202 6310 2204
rect 6366 2202 6390 2204
rect 6446 2202 6452 2204
rect 6206 2150 6208 2202
rect 6388 2150 6390 2202
rect 6144 2148 6150 2150
rect 6206 2148 6230 2150
rect 6286 2148 6310 2150
rect 6366 2148 6390 2150
rect 6446 2148 6452 2150
rect 6144 2128 6452 2148
rect 7484 1193 7512 2382
rect 7852 2281 7880 2790
rect 7838 2272 7894 2281
rect 7838 2207 7894 2216
rect 7470 1184 7526 1193
rect 7470 1119 7526 1128
rect 4986 0 5042 800
rect 8036 649 8064 2790
rect 8114 2751 8170 2760
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8022 640 8078 649
rect 8022 575 8078 584
rect 8128 241 8156 2382
rect 8220 1737 8248 3470
rect 8206 1728 8262 1737
rect 8206 1663 8262 1672
rect 8114 232 8170 241
rect 8114 167 8170 176
<< via2 >>
rect 6642 24656 6698 24712
rect 2254 22330 2310 22332
rect 2334 22330 2390 22332
rect 2414 22330 2470 22332
rect 2494 22330 2550 22332
rect 2254 22278 2300 22330
rect 2300 22278 2310 22330
rect 2334 22278 2364 22330
rect 2364 22278 2376 22330
rect 2376 22278 2390 22330
rect 2414 22278 2428 22330
rect 2428 22278 2440 22330
rect 2440 22278 2470 22330
rect 2494 22278 2504 22330
rect 2504 22278 2550 22330
rect 2254 22276 2310 22278
rect 2334 22276 2390 22278
rect 2414 22276 2470 22278
rect 2494 22276 2550 22278
rect 4852 22330 4908 22332
rect 4932 22330 4988 22332
rect 5012 22330 5068 22332
rect 5092 22330 5148 22332
rect 4852 22278 4898 22330
rect 4898 22278 4908 22330
rect 4932 22278 4962 22330
rect 4962 22278 4974 22330
rect 4974 22278 4988 22330
rect 5012 22278 5026 22330
rect 5026 22278 5038 22330
rect 5038 22278 5068 22330
rect 5092 22278 5102 22330
rect 5102 22278 5148 22330
rect 4852 22276 4908 22278
rect 4932 22276 4988 22278
rect 5012 22276 5068 22278
rect 5092 22276 5148 22278
rect 3553 21786 3609 21788
rect 3633 21786 3689 21788
rect 3713 21786 3769 21788
rect 3793 21786 3849 21788
rect 3553 21734 3599 21786
rect 3599 21734 3609 21786
rect 3633 21734 3663 21786
rect 3663 21734 3675 21786
rect 3675 21734 3689 21786
rect 3713 21734 3727 21786
rect 3727 21734 3739 21786
rect 3739 21734 3769 21786
rect 3793 21734 3803 21786
rect 3803 21734 3849 21786
rect 3553 21732 3609 21734
rect 3633 21732 3689 21734
rect 3713 21732 3769 21734
rect 3793 21732 3849 21734
rect 6150 21786 6206 21788
rect 6230 21786 6286 21788
rect 6310 21786 6366 21788
rect 6390 21786 6446 21788
rect 6150 21734 6196 21786
rect 6196 21734 6206 21786
rect 6230 21734 6260 21786
rect 6260 21734 6272 21786
rect 6272 21734 6286 21786
rect 6310 21734 6324 21786
rect 6324 21734 6336 21786
rect 6336 21734 6366 21786
rect 6390 21734 6400 21786
rect 6400 21734 6446 21786
rect 6150 21732 6206 21734
rect 6230 21732 6286 21734
rect 6310 21732 6366 21734
rect 6390 21732 6446 21734
rect 7838 24112 7894 24168
rect 6734 23568 6790 23624
rect 6826 23024 6882 23080
rect 7449 22330 7505 22332
rect 7529 22330 7585 22332
rect 7609 22330 7665 22332
rect 7689 22330 7745 22332
rect 7449 22278 7495 22330
rect 7495 22278 7505 22330
rect 7529 22278 7559 22330
rect 7559 22278 7571 22330
rect 7571 22278 7585 22330
rect 7609 22278 7623 22330
rect 7623 22278 7635 22330
rect 7635 22278 7665 22330
rect 7689 22278 7699 22330
rect 7699 22278 7745 22330
rect 7449 22276 7505 22278
rect 7529 22276 7585 22278
rect 7609 22276 7665 22278
rect 7689 22276 7745 22278
rect 7470 21412 7526 21448
rect 7470 21392 7472 21412
rect 7472 21392 7524 21412
rect 7524 21392 7526 21412
rect 2254 21242 2310 21244
rect 2334 21242 2390 21244
rect 2414 21242 2470 21244
rect 2494 21242 2550 21244
rect 2254 21190 2300 21242
rect 2300 21190 2310 21242
rect 2334 21190 2364 21242
rect 2364 21190 2376 21242
rect 2376 21190 2390 21242
rect 2414 21190 2428 21242
rect 2428 21190 2440 21242
rect 2440 21190 2470 21242
rect 2494 21190 2504 21242
rect 2504 21190 2550 21242
rect 2254 21188 2310 21190
rect 2334 21188 2390 21190
rect 2414 21188 2470 21190
rect 2494 21188 2550 21190
rect 4852 21242 4908 21244
rect 4932 21242 4988 21244
rect 5012 21242 5068 21244
rect 5092 21242 5148 21244
rect 4852 21190 4898 21242
rect 4898 21190 4908 21242
rect 4932 21190 4962 21242
rect 4962 21190 4974 21242
rect 4974 21190 4988 21242
rect 5012 21190 5026 21242
rect 5026 21190 5038 21242
rect 5038 21190 5068 21242
rect 5092 21190 5102 21242
rect 5102 21190 5148 21242
rect 4852 21188 4908 21190
rect 4932 21188 4988 21190
rect 5012 21188 5068 21190
rect 5092 21188 5148 21190
rect 7449 21242 7505 21244
rect 7529 21242 7585 21244
rect 7609 21242 7665 21244
rect 7689 21242 7745 21244
rect 7449 21190 7495 21242
rect 7495 21190 7505 21242
rect 7529 21190 7559 21242
rect 7559 21190 7571 21242
rect 7571 21190 7585 21242
rect 7609 21190 7623 21242
rect 7623 21190 7635 21242
rect 7635 21190 7665 21242
rect 7689 21190 7699 21242
rect 7699 21190 7745 21242
rect 7449 21188 7505 21190
rect 7529 21188 7585 21190
rect 7609 21188 7665 21190
rect 7689 21188 7745 21190
rect 8206 22480 8262 22536
rect 8114 21956 8170 21992
rect 8114 21936 8116 21956
rect 8116 21936 8168 21956
rect 8168 21936 8170 21956
rect 8114 20884 8116 20904
rect 8116 20884 8168 20904
rect 8168 20884 8170 20904
rect 8114 20848 8170 20884
rect 3553 20698 3609 20700
rect 3633 20698 3689 20700
rect 3713 20698 3769 20700
rect 3793 20698 3849 20700
rect 3553 20646 3599 20698
rect 3599 20646 3609 20698
rect 3633 20646 3663 20698
rect 3663 20646 3675 20698
rect 3675 20646 3689 20698
rect 3713 20646 3727 20698
rect 3727 20646 3739 20698
rect 3739 20646 3769 20698
rect 3793 20646 3803 20698
rect 3803 20646 3849 20698
rect 3553 20644 3609 20646
rect 3633 20644 3689 20646
rect 3713 20644 3769 20646
rect 3793 20644 3849 20646
rect 6150 20698 6206 20700
rect 6230 20698 6286 20700
rect 6310 20698 6366 20700
rect 6390 20698 6446 20700
rect 6150 20646 6196 20698
rect 6196 20646 6206 20698
rect 6230 20646 6260 20698
rect 6260 20646 6272 20698
rect 6272 20646 6286 20698
rect 6310 20646 6324 20698
rect 6324 20646 6336 20698
rect 6336 20646 6366 20698
rect 6390 20646 6400 20698
rect 6400 20646 6446 20698
rect 6150 20644 6206 20646
rect 6230 20644 6286 20646
rect 6310 20644 6366 20646
rect 6390 20644 6446 20646
rect 8114 20340 8116 20360
rect 8116 20340 8168 20360
rect 8168 20340 8170 20360
rect 8114 20304 8170 20340
rect 2254 20154 2310 20156
rect 2334 20154 2390 20156
rect 2414 20154 2470 20156
rect 2494 20154 2550 20156
rect 2254 20102 2300 20154
rect 2300 20102 2310 20154
rect 2334 20102 2364 20154
rect 2364 20102 2376 20154
rect 2376 20102 2390 20154
rect 2414 20102 2428 20154
rect 2428 20102 2440 20154
rect 2440 20102 2470 20154
rect 2494 20102 2504 20154
rect 2504 20102 2550 20154
rect 2254 20100 2310 20102
rect 2334 20100 2390 20102
rect 2414 20100 2470 20102
rect 2494 20100 2550 20102
rect 4852 20154 4908 20156
rect 4932 20154 4988 20156
rect 5012 20154 5068 20156
rect 5092 20154 5148 20156
rect 4852 20102 4898 20154
rect 4898 20102 4908 20154
rect 4932 20102 4962 20154
rect 4962 20102 4974 20154
rect 4974 20102 4988 20154
rect 5012 20102 5026 20154
rect 5026 20102 5038 20154
rect 5038 20102 5068 20154
rect 5092 20102 5102 20154
rect 5102 20102 5148 20154
rect 4852 20100 4908 20102
rect 4932 20100 4988 20102
rect 5012 20100 5068 20102
rect 5092 20100 5148 20102
rect 7449 20154 7505 20156
rect 7529 20154 7585 20156
rect 7609 20154 7665 20156
rect 7689 20154 7745 20156
rect 7449 20102 7495 20154
rect 7495 20102 7505 20154
rect 7529 20102 7559 20154
rect 7559 20102 7571 20154
rect 7571 20102 7585 20154
rect 7609 20102 7623 20154
rect 7623 20102 7635 20154
rect 7635 20102 7665 20154
rect 7689 20102 7699 20154
rect 7699 20102 7745 20154
rect 7449 20100 7505 20102
rect 7529 20100 7585 20102
rect 7609 20100 7665 20102
rect 7689 20100 7745 20102
rect 8114 19780 8170 19816
rect 8114 19760 8116 19780
rect 8116 19760 8168 19780
rect 8168 19760 8170 19780
rect 3553 19610 3609 19612
rect 3633 19610 3689 19612
rect 3713 19610 3769 19612
rect 3793 19610 3849 19612
rect 3553 19558 3599 19610
rect 3599 19558 3609 19610
rect 3633 19558 3663 19610
rect 3663 19558 3675 19610
rect 3675 19558 3689 19610
rect 3713 19558 3727 19610
rect 3727 19558 3739 19610
rect 3739 19558 3769 19610
rect 3793 19558 3803 19610
rect 3803 19558 3849 19610
rect 3553 19556 3609 19558
rect 3633 19556 3689 19558
rect 3713 19556 3769 19558
rect 3793 19556 3849 19558
rect 6150 19610 6206 19612
rect 6230 19610 6286 19612
rect 6310 19610 6366 19612
rect 6390 19610 6446 19612
rect 6150 19558 6196 19610
rect 6196 19558 6206 19610
rect 6230 19558 6260 19610
rect 6260 19558 6272 19610
rect 6272 19558 6286 19610
rect 6310 19558 6324 19610
rect 6324 19558 6336 19610
rect 6336 19558 6366 19610
rect 6390 19558 6400 19610
rect 6400 19558 6446 19610
rect 6150 19556 6206 19558
rect 6230 19556 6286 19558
rect 6310 19556 6366 19558
rect 6390 19556 6446 19558
rect 7470 19236 7526 19272
rect 7470 19216 7472 19236
rect 7472 19216 7524 19236
rect 7524 19216 7526 19236
rect 2254 19066 2310 19068
rect 2334 19066 2390 19068
rect 2414 19066 2470 19068
rect 2494 19066 2550 19068
rect 2254 19014 2300 19066
rect 2300 19014 2310 19066
rect 2334 19014 2364 19066
rect 2364 19014 2376 19066
rect 2376 19014 2390 19066
rect 2414 19014 2428 19066
rect 2428 19014 2440 19066
rect 2440 19014 2470 19066
rect 2494 19014 2504 19066
rect 2504 19014 2550 19066
rect 2254 19012 2310 19014
rect 2334 19012 2390 19014
rect 2414 19012 2470 19014
rect 2494 19012 2550 19014
rect 4852 19066 4908 19068
rect 4932 19066 4988 19068
rect 5012 19066 5068 19068
rect 5092 19066 5148 19068
rect 4852 19014 4898 19066
rect 4898 19014 4908 19066
rect 4932 19014 4962 19066
rect 4962 19014 4974 19066
rect 4974 19014 4988 19066
rect 5012 19014 5026 19066
rect 5026 19014 5038 19066
rect 5038 19014 5068 19066
rect 5092 19014 5102 19066
rect 5102 19014 5148 19066
rect 4852 19012 4908 19014
rect 4932 19012 4988 19014
rect 5012 19012 5068 19014
rect 5092 19012 5148 19014
rect 7449 19066 7505 19068
rect 7529 19066 7585 19068
rect 7609 19066 7665 19068
rect 7689 19066 7745 19068
rect 7449 19014 7495 19066
rect 7495 19014 7505 19066
rect 7529 19014 7559 19066
rect 7559 19014 7571 19066
rect 7571 19014 7585 19066
rect 7609 19014 7623 19066
rect 7623 19014 7635 19066
rect 7635 19014 7665 19066
rect 7689 19014 7699 19066
rect 7699 19014 7745 19066
rect 7449 19012 7505 19014
rect 7529 19012 7585 19014
rect 7609 19012 7665 19014
rect 7689 19012 7745 19014
rect 8114 18808 8170 18864
rect 3553 18522 3609 18524
rect 3633 18522 3689 18524
rect 3713 18522 3769 18524
rect 3793 18522 3849 18524
rect 3553 18470 3599 18522
rect 3599 18470 3609 18522
rect 3633 18470 3663 18522
rect 3663 18470 3675 18522
rect 3675 18470 3689 18522
rect 3713 18470 3727 18522
rect 3727 18470 3739 18522
rect 3739 18470 3769 18522
rect 3793 18470 3803 18522
rect 3803 18470 3849 18522
rect 3553 18468 3609 18470
rect 3633 18468 3689 18470
rect 3713 18468 3769 18470
rect 3793 18468 3849 18470
rect 6150 18522 6206 18524
rect 6230 18522 6286 18524
rect 6310 18522 6366 18524
rect 6390 18522 6446 18524
rect 6150 18470 6196 18522
rect 6196 18470 6206 18522
rect 6230 18470 6260 18522
rect 6260 18470 6272 18522
rect 6272 18470 6286 18522
rect 6310 18470 6324 18522
rect 6324 18470 6336 18522
rect 6336 18470 6366 18522
rect 6390 18470 6400 18522
rect 6400 18470 6446 18522
rect 6150 18468 6206 18470
rect 6230 18468 6286 18470
rect 6310 18468 6366 18470
rect 6390 18468 6446 18470
rect 8114 18264 8170 18320
rect 2254 17978 2310 17980
rect 2334 17978 2390 17980
rect 2414 17978 2470 17980
rect 2494 17978 2550 17980
rect 2254 17926 2300 17978
rect 2300 17926 2310 17978
rect 2334 17926 2364 17978
rect 2364 17926 2376 17978
rect 2376 17926 2390 17978
rect 2414 17926 2428 17978
rect 2428 17926 2440 17978
rect 2440 17926 2470 17978
rect 2494 17926 2504 17978
rect 2504 17926 2550 17978
rect 2254 17924 2310 17926
rect 2334 17924 2390 17926
rect 2414 17924 2470 17926
rect 2494 17924 2550 17926
rect 4852 17978 4908 17980
rect 4932 17978 4988 17980
rect 5012 17978 5068 17980
rect 5092 17978 5148 17980
rect 4852 17926 4898 17978
rect 4898 17926 4908 17978
rect 4932 17926 4962 17978
rect 4962 17926 4974 17978
rect 4974 17926 4988 17978
rect 5012 17926 5026 17978
rect 5026 17926 5038 17978
rect 5038 17926 5068 17978
rect 5092 17926 5102 17978
rect 5102 17926 5148 17978
rect 4852 17924 4908 17926
rect 4932 17924 4988 17926
rect 5012 17924 5068 17926
rect 5092 17924 5148 17926
rect 7449 17978 7505 17980
rect 7529 17978 7585 17980
rect 7609 17978 7665 17980
rect 7689 17978 7745 17980
rect 7449 17926 7495 17978
rect 7495 17926 7505 17978
rect 7529 17926 7559 17978
rect 7559 17926 7571 17978
rect 7571 17926 7585 17978
rect 7609 17926 7623 17978
rect 7623 17926 7635 17978
rect 7635 17926 7665 17978
rect 7689 17926 7699 17978
rect 7699 17926 7745 17978
rect 7449 17924 7505 17926
rect 7529 17924 7585 17926
rect 7609 17924 7665 17926
rect 7689 17924 7745 17926
rect 8114 17720 8170 17776
rect 3553 17434 3609 17436
rect 3633 17434 3689 17436
rect 3713 17434 3769 17436
rect 3793 17434 3849 17436
rect 3553 17382 3599 17434
rect 3599 17382 3609 17434
rect 3633 17382 3663 17434
rect 3663 17382 3675 17434
rect 3675 17382 3689 17434
rect 3713 17382 3727 17434
rect 3727 17382 3739 17434
rect 3739 17382 3769 17434
rect 3793 17382 3803 17434
rect 3803 17382 3849 17434
rect 3553 17380 3609 17382
rect 3633 17380 3689 17382
rect 3713 17380 3769 17382
rect 3793 17380 3849 17382
rect 6150 17434 6206 17436
rect 6230 17434 6286 17436
rect 6310 17434 6366 17436
rect 6390 17434 6446 17436
rect 6150 17382 6196 17434
rect 6196 17382 6206 17434
rect 6230 17382 6260 17434
rect 6260 17382 6272 17434
rect 6272 17382 6286 17434
rect 6310 17382 6324 17434
rect 6324 17382 6336 17434
rect 6336 17382 6366 17434
rect 6390 17382 6400 17434
rect 6400 17382 6446 17434
rect 6150 17380 6206 17382
rect 6230 17380 6286 17382
rect 6310 17380 6366 17382
rect 6390 17380 6446 17382
rect 8114 17176 8170 17232
rect 2254 16890 2310 16892
rect 2334 16890 2390 16892
rect 2414 16890 2470 16892
rect 2494 16890 2550 16892
rect 2254 16838 2300 16890
rect 2300 16838 2310 16890
rect 2334 16838 2364 16890
rect 2364 16838 2376 16890
rect 2376 16838 2390 16890
rect 2414 16838 2428 16890
rect 2428 16838 2440 16890
rect 2440 16838 2470 16890
rect 2494 16838 2504 16890
rect 2504 16838 2550 16890
rect 2254 16836 2310 16838
rect 2334 16836 2390 16838
rect 2414 16836 2470 16838
rect 2494 16836 2550 16838
rect 4852 16890 4908 16892
rect 4932 16890 4988 16892
rect 5012 16890 5068 16892
rect 5092 16890 5148 16892
rect 4852 16838 4898 16890
rect 4898 16838 4908 16890
rect 4932 16838 4962 16890
rect 4962 16838 4974 16890
rect 4974 16838 4988 16890
rect 5012 16838 5026 16890
rect 5026 16838 5038 16890
rect 5038 16838 5068 16890
rect 5092 16838 5102 16890
rect 5102 16838 5148 16890
rect 4852 16836 4908 16838
rect 4932 16836 4988 16838
rect 5012 16836 5068 16838
rect 5092 16836 5148 16838
rect 7449 16890 7505 16892
rect 7529 16890 7585 16892
rect 7609 16890 7665 16892
rect 7689 16890 7745 16892
rect 7449 16838 7495 16890
rect 7495 16838 7505 16890
rect 7529 16838 7559 16890
rect 7559 16838 7571 16890
rect 7571 16838 7585 16890
rect 7609 16838 7623 16890
rect 7623 16838 7635 16890
rect 7635 16838 7665 16890
rect 7689 16838 7699 16890
rect 7699 16838 7745 16890
rect 7449 16836 7505 16838
rect 7529 16836 7585 16838
rect 7609 16836 7665 16838
rect 7689 16836 7745 16838
rect 8206 16632 8262 16688
rect 3553 16346 3609 16348
rect 3633 16346 3689 16348
rect 3713 16346 3769 16348
rect 3793 16346 3849 16348
rect 3553 16294 3599 16346
rect 3599 16294 3609 16346
rect 3633 16294 3663 16346
rect 3663 16294 3675 16346
rect 3675 16294 3689 16346
rect 3713 16294 3727 16346
rect 3727 16294 3739 16346
rect 3739 16294 3769 16346
rect 3793 16294 3803 16346
rect 3803 16294 3849 16346
rect 3553 16292 3609 16294
rect 3633 16292 3689 16294
rect 3713 16292 3769 16294
rect 3793 16292 3849 16294
rect 6150 16346 6206 16348
rect 6230 16346 6286 16348
rect 6310 16346 6366 16348
rect 6390 16346 6446 16348
rect 6150 16294 6196 16346
rect 6196 16294 6206 16346
rect 6230 16294 6260 16346
rect 6260 16294 6272 16346
rect 6272 16294 6286 16346
rect 6310 16294 6324 16346
rect 6324 16294 6336 16346
rect 6336 16294 6366 16346
rect 6390 16294 6400 16346
rect 6400 16294 6446 16346
rect 6150 16292 6206 16294
rect 6230 16292 6286 16294
rect 6310 16292 6366 16294
rect 6390 16292 6446 16294
rect 8114 16088 8170 16144
rect 2254 15802 2310 15804
rect 2334 15802 2390 15804
rect 2414 15802 2470 15804
rect 2494 15802 2550 15804
rect 2254 15750 2300 15802
rect 2300 15750 2310 15802
rect 2334 15750 2364 15802
rect 2364 15750 2376 15802
rect 2376 15750 2390 15802
rect 2414 15750 2428 15802
rect 2428 15750 2440 15802
rect 2440 15750 2470 15802
rect 2494 15750 2504 15802
rect 2504 15750 2550 15802
rect 2254 15748 2310 15750
rect 2334 15748 2390 15750
rect 2414 15748 2470 15750
rect 2494 15748 2550 15750
rect 4852 15802 4908 15804
rect 4932 15802 4988 15804
rect 5012 15802 5068 15804
rect 5092 15802 5148 15804
rect 4852 15750 4898 15802
rect 4898 15750 4908 15802
rect 4932 15750 4962 15802
rect 4962 15750 4974 15802
rect 4974 15750 4988 15802
rect 5012 15750 5026 15802
rect 5026 15750 5038 15802
rect 5038 15750 5068 15802
rect 5092 15750 5102 15802
rect 5102 15750 5148 15802
rect 4852 15748 4908 15750
rect 4932 15748 4988 15750
rect 5012 15748 5068 15750
rect 5092 15748 5148 15750
rect 7449 15802 7505 15804
rect 7529 15802 7585 15804
rect 7609 15802 7665 15804
rect 7689 15802 7745 15804
rect 7449 15750 7495 15802
rect 7495 15750 7505 15802
rect 7529 15750 7559 15802
rect 7559 15750 7571 15802
rect 7571 15750 7585 15802
rect 7609 15750 7623 15802
rect 7623 15750 7635 15802
rect 7635 15750 7665 15802
rect 7689 15750 7699 15802
rect 7699 15750 7745 15802
rect 7449 15748 7505 15750
rect 7529 15748 7585 15750
rect 7609 15748 7665 15750
rect 7689 15748 7745 15750
rect 8114 15544 8170 15600
rect 3553 15258 3609 15260
rect 3633 15258 3689 15260
rect 3713 15258 3769 15260
rect 3793 15258 3849 15260
rect 3553 15206 3599 15258
rect 3599 15206 3609 15258
rect 3633 15206 3663 15258
rect 3663 15206 3675 15258
rect 3675 15206 3689 15258
rect 3713 15206 3727 15258
rect 3727 15206 3739 15258
rect 3739 15206 3769 15258
rect 3793 15206 3803 15258
rect 3803 15206 3849 15258
rect 3553 15204 3609 15206
rect 3633 15204 3689 15206
rect 3713 15204 3769 15206
rect 3793 15204 3849 15206
rect 6150 15258 6206 15260
rect 6230 15258 6286 15260
rect 6310 15258 6366 15260
rect 6390 15258 6446 15260
rect 6150 15206 6196 15258
rect 6196 15206 6206 15258
rect 6230 15206 6260 15258
rect 6260 15206 6272 15258
rect 6272 15206 6286 15258
rect 6310 15206 6324 15258
rect 6324 15206 6336 15258
rect 6336 15206 6366 15258
rect 6390 15206 6400 15258
rect 6400 15206 6446 15258
rect 6150 15204 6206 15206
rect 6230 15204 6286 15206
rect 6310 15204 6366 15206
rect 6390 15204 6446 15206
rect 8114 15000 8170 15056
rect 2254 14714 2310 14716
rect 2334 14714 2390 14716
rect 2414 14714 2470 14716
rect 2494 14714 2550 14716
rect 2254 14662 2300 14714
rect 2300 14662 2310 14714
rect 2334 14662 2364 14714
rect 2364 14662 2376 14714
rect 2376 14662 2390 14714
rect 2414 14662 2428 14714
rect 2428 14662 2440 14714
rect 2440 14662 2470 14714
rect 2494 14662 2504 14714
rect 2504 14662 2550 14714
rect 2254 14660 2310 14662
rect 2334 14660 2390 14662
rect 2414 14660 2470 14662
rect 2494 14660 2550 14662
rect 4852 14714 4908 14716
rect 4932 14714 4988 14716
rect 5012 14714 5068 14716
rect 5092 14714 5148 14716
rect 4852 14662 4898 14714
rect 4898 14662 4908 14714
rect 4932 14662 4962 14714
rect 4962 14662 4974 14714
rect 4974 14662 4988 14714
rect 5012 14662 5026 14714
rect 5026 14662 5038 14714
rect 5038 14662 5068 14714
rect 5092 14662 5102 14714
rect 5102 14662 5148 14714
rect 4852 14660 4908 14662
rect 4932 14660 4988 14662
rect 5012 14660 5068 14662
rect 5092 14660 5148 14662
rect 7449 14714 7505 14716
rect 7529 14714 7585 14716
rect 7609 14714 7665 14716
rect 7689 14714 7745 14716
rect 7449 14662 7495 14714
rect 7495 14662 7505 14714
rect 7529 14662 7559 14714
rect 7559 14662 7571 14714
rect 7571 14662 7585 14714
rect 7609 14662 7623 14714
rect 7623 14662 7635 14714
rect 7635 14662 7665 14714
rect 7689 14662 7699 14714
rect 7699 14662 7745 14714
rect 7449 14660 7505 14662
rect 7529 14660 7585 14662
rect 7609 14660 7665 14662
rect 7689 14660 7745 14662
rect 8114 14456 8170 14512
rect 3553 14170 3609 14172
rect 3633 14170 3689 14172
rect 3713 14170 3769 14172
rect 3793 14170 3849 14172
rect 3553 14118 3599 14170
rect 3599 14118 3609 14170
rect 3633 14118 3663 14170
rect 3663 14118 3675 14170
rect 3675 14118 3689 14170
rect 3713 14118 3727 14170
rect 3727 14118 3739 14170
rect 3739 14118 3769 14170
rect 3793 14118 3803 14170
rect 3803 14118 3849 14170
rect 3553 14116 3609 14118
rect 3633 14116 3689 14118
rect 3713 14116 3769 14118
rect 3793 14116 3849 14118
rect 6150 14170 6206 14172
rect 6230 14170 6286 14172
rect 6310 14170 6366 14172
rect 6390 14170 6446 14172
rect 6150 14118 6196 14170
rect 6196 14118 6206 14170
rect 6230 14118 6260 14170
rect 6260 14118 6272 14170
rect 6272 14118 6286 14170
rect 6310 14118 6324 14170
rect 6324 14118 6336 14170
rect 6336 14118 6366 14170
rect 6390 14118 6400 14170
rect 6400 14118 6446 14170
rect 6150 14116 6206 14118
rect 6230 14116 6286 14118
rect 6310 14116 6366 14118
rect 6390 14116 6446 14118
rect 8114 13912 8170 13968
rect 2254 13626 2310 13628
rect 2334 13626 2390 13628
rect 2414 13626 2470 13628
rect 2494 13626 2550 13628
rect 2254 13574 2300 13626
rect 2300 13574 2310 13626
rect 2334 13574 2364 13626
rect 2364 13574 2376 13626
rect 2376 13574 2390 13626
rect 2414 13574 2428 13626
rect 2428 13574 2440 13626
rect 2440 13574 2470 13626
rect 2494 13574 2504 13626
rect 2504 13574 2550 13626
rect 2254 13572 2310 13574
rect 2334 13572 2390 13574
rect 2414 13572 2470 13574
rect 2494 13572 2550 13574
rect 4852 13626 4908 13628
rect 4932 13626 4988 13628
rect 5012 13626 5068 13628
rect 5092 13626 5148 13628
rect 4852 13574 4898 13626
rect 4898 13574 4908 13626
rect 4932 13574 4962 13626
rect 4962 13574 4974 13626
rect 4974 13574 4988 13626
rect 5012 13574 5026 13626
rect 5026 13574 5038 13626
rect 5038 13574 5068 13626
rect 5092 13574 5102 13626
rect 5102 13574 5148 13626
rect 4852 13572 4908 13574
rect 4932 13572 4988 13574
rect 5012 13572 5068 13574
rect 5092 13572 5148 13574
rect 7449 13626 7505 13628
rect 7529 13626 7585 13628
rect 7609 13626 7665 13628
rect 7689 13626 7745 13628
rect 7449 13574 7495 13626
rect 7495 13574 7505 13626
rect 7529 13574 7559 13626
rect 7559 13574 7571 13626
rect 7571 13574 7585 13626
rect 7609 13574 7623 13626
rect 7623 13574 7635 13626
rect 7635 13574 7665 13626
rect 7689 13574 7699 13626
rect 7699 13574 7745 13626
rect 7449 13572 7505 13574
rect 7529 13572 7585 13574
rect 7609 13572 7665 13574
rect 7689 13572 7745 13574
rect 8114 13368 8170 13424
rect 3553 13082 3609 13084
rect 3633 13082 3689 13084
rect 3713 13082 3769 13084
rect 3793 13082 3849 13084
rect 3553 13030 3599 13082
rect 3599 13030 3609 13082
rect 3633 13030 3663 13082
rect 3663 13030 3675 13082
rect 3675 13030 3689 13082
rect 3713 13030 3727 13082
rect 3727 13030 3739 13082
rect 3739 13030 3769 13082
rect 3793 13030 3803 13082
rect 3803 13030 3849 13082
rect 3553 13028 3609 13030
rect 3633 13028 3689 13030
rect 3713 13028 3769 13030
rect 3793 13028 3849 13030
rect 6150 13082 6206 13084
rect 6230 13082 6286 13084
rect 6310 13082 6366 13084
rect 6390 13082 6446 13084
rect 6150 13030 6196 13082
rect 6196 13030 6206 13082
rect 6230 13030 6260 13082
rect 6260 13030 6272 13082
rect 6272 13030 6286 13082
rect 6310 13030 6324 13082
rect 6324 13030 6336 13082
rect 6336 13030 6366 13082
rect 6390 13030 6400 13082
rect 6400 13030 6446 13082
rect 6150 13028 6206 13030
rect 6230 13028 6286 13030
rect 6310 13028 6366 13030
rect 6390 13028 6446 13030
rect 8114 12824 8170 12880
rect 2254 12538 2310 12540
rect 2334 12538 2390 12540
rect 2414 12538 2470 12540
rect 2494 12538 2550 12540
rect 2254 12486 2300 12538
rect 2300 12486 2310 12538
rect 2334 12486 2364 12538
rect 2364 12486 2376 12538
rect 2376 12486 2390 12538
rect 2414 12486 2428 12538
rect 2428 12486 2440 12538
rect 2440 12486 2470 12538
rect 2494 12486 2504 12538
rect 2504 12486 2550 12538
rect 2254 12484 2310 12486
rect 2334 12484 2390 12486
rect 2414 12484 2470 12486
rect 2494 12484 2550 12486
rect 4852 12538 4908 12540
rect 4932 12538 4988 12540
rect 5012 12538 5068 12540
rect 5092 12538 5148 12540
rect 4852 12486 4898 12538
rect 4898 12486 4908 12538
rect 4932 12486 4962 12538
rect 4962 12486 4974 12538
rect 4974 12486 4988 12538
rect 5012 12486 5026 12538
rect 5026 12486 5038 12538
rect 5038 12486 5068 12538
rect 5092 12486 5102 12538
rect 5102 12486 5148 12538
rect 4852 12484 4908 12486
rect 4932 12484 4988 12486
rect 5012 12484 5068 12486
rect 5092 12484 5148 12486
rect 7449 12538 7505 12540
rect 7529 12538 7585 12540
rect 7609 12538 7665 12540
rect 7689 12538 7745 12540
rect 7449 12486 7495 12538
rect 7495 12486 7505 12538
rect 7529 12486 7559 12538
rect 7559 12486 7571 12538
rect 7571 12486 7585 12538
rect 7609 12486 7623 12538
rect 7623 12486 7635 12538
rect 7635 12486 7665 12538
rect 7689 12486 7699 12538
rect 7699 12486 7745 12538
rect 7449 12484 7505 12486
rect 7529 12484 7585 12486
rect 7609 12484 7665 12486
rect 7689 12484 7745 12486
rect 8114 12416 8170 12472
rect 3553 11994 3609 11996
rect 3633 11994 3689 11996
rect 3713 11994 3769 11996
rect 3793 11994 3849 11996
rect 3553 11942 3599 11994
rect 3599 11942 3609 11994
rect 3633 11942 3663 11994
rect 3663 11942 3675 11994
rect 3675 11942 3689 11994
rect 3713 11942 3727 11994
rect 3727 11942 3739 11994
rect 3739 11942 3769 11994
rect 3793 11942 3803 11994
rect 3803 11942 3849 11994
rect 3553 11940 3609 11942
rect 3633 11940 3689 11942
rect 3713 11940 3769 11942
rect 3793 11940 3849 11942
rect 6150 11994 6206 11996
rect 6230 11994 6286 11996
rect 6310 11994 6366 11996
rect 6390 11994 6446 11996
rect 6150 11942 6196 11994
rect 6196 11942 6206 11994
rect 6230 11942 6260 11994
rect 6260 11942 6272 11994
rect 6272 11942 6286 11994
rect 6310 11942 6324 11994
rect 6324 11942 6336 11994
rect 6336 11942 6366 11994
rect 6390 11942 6400 11994
rect 6400 11942 6446 11994
rect 6150 11940 6206 11942
rect 6230 11940 6286 11942
rect 6310 11940 6366 11942
rect 6390 11940 6446 11942
rect 8114 11872 8170 11928
rect 2254 11450 2310 11452
rect 2334 11450 2390 11452
rect 2414 11450 2470 11452
rect 2494 11450 2550 11452
rect 2254 11398 2300 11450
rect 2300 11398 2310 11450
rect 2334 11398 2364 11450
rect 2364 11398 2376 11450
rect 2376 11398 2390 11450
rect 2414 11398 2428 11450
rect 2428 11398 2440 11450
rect 2440 11398 2470 11450
rect 2494 11398 2504 11450
rect 2504 11398 2550 11450
rect 2254 11396 2310 11398
rect 2334 11396 2390 11398
rect 2414 11396 2470 11398
rect 2494 11396 2550 11398
rect 4852 11450 4908 11452
rect 4932 11450 4988 11452
rect 5012 11450 5068 11452
rect 5092 11450 5148 11452
rect 4852 11398 4898 11450
rect 4898 11398 4908 11450
rect 4932 11398 4962 11450
rect 4962 11398 4974 11450
rect 4974 11398 4988 11450
rect 5012 11398 5026 11450
rect 5026 11398 5038 11450
rect 5038 11398 5068 11450
rect 5092 11398 5102 11450
rect 5102 11398 5148 11450
rect 4852 11396 4908 11398
rect 4932 11396 4988 11398
rect 5012 11396 5068 11398
rect 5092 11396 5148 11398
rect 7449 11450 7505 11452
rect 7529 11450 7585 11452
rect 7609 11450 7665 11452
rect 7689 11450 7745 11452
rect 7449 11398 7495 11450
rect 7495 11398 7505 11450
rect 7529 11398 7559 11450
rect 7559 11398 7571 11450
rect 7571 11398 7585 11450
rect 7609 11398 7623 11450
rect 7623 11398 7635 11450
rect 7635 11398 7665 11450
rect 7689 11398 7699 11450
rect 7699 11398 7745 11450
rect 7449 11396 7505 11398
rect 7529 11396 7585 11398
rect 7609 11396 7665 11398
rect 7689 11396 7745 11398
rect 8114 11328 8170 11384
rect 3553 10906 3609 10908
rect 3633 10906 3689 10908
rect 3713 10906 3769 10908
rect 3793 10906 3849 10908
rect 3553 10854 3599 10906
rect 3599 10854 3609 10906
rect 3633 10854 3663 10906
rect 3663 10854 3675 10906
rect 3675 10854 3689 10906
rect 3713 10854 3727 10906
rect 3727 10854 3739 10906
rect 3739 10854 3769 10906
rect 3793 10854 3803 10906
rect 3803 10854 3849 10906
rect 3553 10852 3609 10854
rect 3633 10852 3689 10854
rect 3713 10852 3769 10854
rect 3793 10852 3849 10854
rect 6150 10906 6206 10908
rect 6230 10906 6286 10908
rect 6310 10906 6366 10908
rect 6390 10906 6446 10908
rect 6150 10854 6196 10906
rect 6196 10854 6206 10906
rect 6230 10854 6260 10906
rect 6260 10854 6272 10906
rect 6272 10854 6286 10906
rect 6310 10854 6324 10906
rect 6324 10854 6336 10906
rect 6336 10854 6366 10906
rect 6390 10854 6400 10906
rect 6400 10854 6446 10906
rect 6150 10852 6206 10854
rect 6230 10852 6286 10854
rect 6310 10852 6366 10854
rect 6390 10852 6446 10854
rect 8114 10784 8170 10840
rect 2254 10362 2310 10364
rect 2334 10362 2390 10364
rect 2414 10362 2470 10364
rect 2494 10362 2550 10364
rect 2254 10310 2300 10362
rect 2300 10310 2310 10362
rect 2334 10310 2364 10362
rect 2364 10310 2376 10362
rect 2376 10310 2390 10362
rect 2414 10310 2428 10362
rect 2428 10310 2440 10362
rect 2440 10310 2470 10362
rect 2494 10310 2504 10362
rect 2504 10310 2550 10362
rect 2254 10308 2310 10310
rect 2334 10308 2390 10310
rect 2414 10308 2470 10310
rect 2494 10308 2550 10310
rect 4852 10362 4908 10364
rect 4932 10362 4988 10364
rect 5012 10362 5068 10364
rect 5092 10362 5148 10364
rect 4852 10310 4898 10362
rect 4898 10310 4908 10362
rect 4932 10310 4962 10362
rect 4962 10310 4974 10362
rect 4974 10310 4988 10362
rect 5012 10310 5026 10362
rect 5026 10310 5038 10362
rect 5038 10310 5068 10362
rect 5092 10310 5102 10362
rect 5102 10310 5148 10362
rect 4852 10308 4908 10310
rect 4932 10308 4988 10310
rect 5012 10308 5068 10310
rect 5092 10308 5148 10310
rect 7449 10362 7505 10364
rect 7529 10362 7585 10364
rect 7609 10362 7665 10364
rect 7689 10362 7745 10364
rect 7449 10310 7495 10362
rect 7495 10310 7505 10362
rect 7529 10310 7559 10362
rect 7559 10310 7571 10362
rect 7571 10310 7585 10362
rect 7609 10310 7623 10362
rect 7623 10310 7635 10362
rect 7635 10310 7665 10362
rect 7689 10310 7699 10362
rect 7699 10310 7745 10362
rect 7449 10308 7505 10310
rect 7529 10308 7585 10310
rect 7609 10308 7665 10310
rect 7689 10308 7745 10310
rect 8114 10240 8170 10296
rect 3553 9818 3609 9820
rect 3633 9818 3689 9820
rect 3713 9818 3769 9820
rect 3793 9818 3849 9820
rect 3553 9766 3599 9818
rect 3599 9766 3609 9818
rect 3633 9766 3663 9818
rect 3663 9766 3675 9818
rect 3675 9766 3689 9818
rect 3713 9766 3727 9818
rect 3727 9766 3739 9818
rect 3739 9766 3769 9818
rect 3793 9766 3803 9818
rect 3803 9766 3849 9818
rect 3553 9764 3609 9766
rect 3633 9764 3689 9766
rect 3713 9764 3769 9766
rect 3793 9764 3849 9766
rect 6150 9818 6206 9820
rect 6230 9818 6286 9820
rect 6310 9818 6366 9820
rect 6390 9818 6446 9820
rect 6150 9766 6196 9818
rect 6196 9766 6206 9818
rect 6230 9766 6260 9818
rect 6260 9766 6272 9818
rect 6272 9766 6286 9818
rect 6310 9766 6324 9818
rect 6324 9766 6336 9818
rect 6336 9766 6366 9818
rect 6390 9766 6400 9818
rect 6400 9766 6446 9818
rect 6150 9764 6206 9766
rect 6230 9764 6286 9766
rect 6310 9764 6366 9766
rect 6390 9764 6446 9766
rect 8114 9696 8170 9752
rect 2254 9274 2310 9276
rect 2334 9274 2390 9276
rect 2414 9274 2470 9276
rect 2494 9274 2550 9276
rect 2254 9222 2300 9274
rect 2300 9222 2310 9274
rect 2334 9222 2364 9274
rect 2364 9222 2376 9274
rect 2376 9222 2390 9274
rect 2414 9222 2428 9274
rect 2428 9222 2440 9274
rect 2440 9222 2470 9274
rect 2494 9222 2504 9274
rect 2504 9222 2550 9274
rect 2254 9220 2310 9222
rect 2334 9220 2390 9222
rect 2414 9220 2470 9222
rect 2494 9220 2550 9222
rect 4852 9274 4908 9276
rect 4932 9274 4988 9276
rect 5012 9274 5068 9276
rect 5092 9274 5148 9276
rect 4852 9222 4898 9274
rect 4898 9222 4908 9274
rect 4932 9222 4962 9274
rect 4962 9222 4974 9274
rect 4974 9222 4988 9274
rect 5012 9222 5026 9274
rect 5026 9222 5038 9274
rect 5038 9222 5068 9274
rect 5092 9222 5102 9274
rect 5102 9222 5148 9274
rect 4852 9220 4908 9222
rect 4932 9220 4988 9222
rect 5012 9220 5068 9222
rect 5092 9220 5148 9222
rect 7449 9274 7505 9276
rect 7529 9274 7585 9276
rect 7609 9274 7665 9276
rect 7689 9274 7745 9276
rect 7449 9222 7495 9274
rect 7495 9222 7505 9274
rect 7529 9222 7559 9274
rect 7559 9222 7571 9274
rect 7571 9222 7585 9274
rect 7609 9222 7623 9274
rect 7623 9222 7635 9274
rect 7635 9222 7665 9274
rect 7689 9222 7699 9274
rect 7699 9222 7745 9274
rect 7449 9220 7505 9222
rect 7529 9220 7585 9222
rect 7609 9220 7665 9222
rect 7689 9220 7745 9222
rect 8114 9152 8170 9208
rect 3553 8730 3609 8732
rect 3633 8730 3689 8732
rect 3713 8730 3769 8732
rect 3793 8730 3849 8732
rect 3553 8678 3599 8730
rect 3599 8678 3609 8730
rect 3633 8678 3663 8730
rect 3663 8678 3675 8730
rect 3675 8678 3689 8730
rect 3713 8678 3727 8730
rect 3727 8678 3739 8730
rect 3739 8678 3769 8730
rect 3793 8678 3803 8730
rect 3803 8678 3849 8730
rect 3553 8676 3609 8678
rect 3633 8676 3689 8678
rect 3713 8676 3769 8678
rect 3793 8676 3849 8678
rect 6150 8730 6206 8732
rect 6230 8730 6286 8732
rect 6310 8730 6366 8732
rect 6390 8730 6446 8732
rect 6150 8678 6196 8730
rect 6196 8678 6206 8730
rect 6230 8678 6260 8730
rect 6260 8678 6272 8730
rect 6272 8678 6286 8730
rect 6310 8678 6324 8730
rect 6324 8678 6336 8730
rect 6336 8678 6366 8730
rect 6390 8678 6400 8730
rect 6400 8678 6446 8730
rect 6150 8676 6206 8678
rect 6230 8676 6286 8678
rect 6310 8676 6366 8678
rect 6390 8676 6446 8678
rect 8114 8608 8170 8664
rect 2254 8186 2310 8188
rect 2334 8186 2390 8188
rect 2414 8186 2470 8188
rect 2494 8186 2550 8188
rect 2254 8134 2300 8186
rect 2300 8134 2310 8186
rect 2334 8134 2364 8186
rect 2364 8134 2376 8186
rect 2376 8134 2390 8186
rect 2414 8134 2428 8186
rect 2428 8134 2440 8186
rect 2440 8134 2470 8186
rect 2494 8134 2504 8186
rect 2504 8134 2550 8186
rect 2254 8132 2310 8134
rect 2334 8132 2390 8134
rect 2414 8132 2470 8134
rect 2494 8132 2550 8134
rect 4852 8186 4908 8188
rect 4932 8186 4988 8188
rect 5012 8186 5068 8188
rect 5092 8186 5148 8188
rect 4852 8134 4898 8186
rect 4898 8134 4908 8186
rect 4932 8134 4962 8186
rect 4962 8134 4974 8186
rect 4974 8134 4988 8186
rect 5012 8134 5026 8186
rect 5026 8134 5038 8186
rect 5038 8134 5068 8186
rect 5092 8134 5102 8186
rect 5102 8134 5148 8186
rect 4852 8132 4908 8134
rect 4932 8132 4988 8134
rect 5012 8132 5068 8134
rect 5092 8132 5148 8134
rect 7449 8186 7505 8188
rect 7529 8186 7585 8188
rect 7609 8186 7665 8188
rect 7689 8186 7745 8188
rect 7449 8134 7495 8186
rect 7495 8134 7505 8186
rect 7529 8134 7559 8186
rect 7559 8134 7571 8186
rect 7571 8134 7585 8186
rect 7609 8134 7623 8186
rect 7623 8134 7635 8186
rect 7635 8134 7665 8186
rect 7689 8134 7699 8186
rect 7699 8134 7745 8186
rect 7449 8132 7505 8134
rect 7529 8132 7585 8134
rect 7609 8132 7665 8134
rect 7689 8132 7745 8134
rect 8114 8064 8170 8120
rect 3553 7642 3609 7644
rect 3633 7642 3689 7644
rect 3713 7642 3769 7644
rect 3793 7642 3849 7644
rect 3553 7590 3599 7642
rect 3599 7590 3609 7642
rect 3633 7590 3663 7642
rect 3663 7590 3675 7642
rect 3675 7590 3689 7642
rect 3713 7590 3727 7642
rect 3727 7590 3739 7642
rect 3739 7590 3769 7642
rect 3793 7590 3803 7642
rect 3803 7590 3849 7642
rect 3553 7588 3609 7590
rect 3633 7588 3689 7590
rect 3713 7588 3769 7590
rect 3793 7588 3849 7590
rect 6150 7642 6206 7644
rect 6230 7642 6286 7644
rect 6310 7642 6366 7644
rect 6390 7642 6446 7644
rect 6150 7590 6196 7642
rect 6196 7590 6206 7642
rect 6230 7590 6260 7642
rect 6260 7590 6272 7642
rect 6272 7590 6286 7642
rect 6310 7590 6324 7642
rect 6324 7590 6336 7642
rect 6336 7590 6366 7642
rect 6390 7590 6400 7642
rect 6400 7590 6446 7642
rect 6150 7588 6206 7590
rect 6230 7588 6286 7590
rect 6310 7588 6366 7590
rect 6390 7588 6446 7590
rect 8114 7520 8170 7576
rect 2254 7098 2310 7100
rect 2334 7098 2390 7100
rect 2414 7098 2470 7100
rect 2494 7098 2550 7100
rect 2254 7046 2300 7098
rect 2300 7046 2310 7098
rect 2334 7046 2364 7098
rect 2364 7046 2376 7098
rect 2376 7046 2390 7098
rect 2414 7046 2428 7098
rect 2428 7046 2440 7098
rect 2440 7046 2470 7098
rect 2494 7046 2504 7098
rect 2504 7046 2550 7098
rect 2254 7044 2310 7046
rect 2334 7044 2390 7046
rect 2414 7044 2470 7046
rect 2494 7044 2550 7046
rect 4852 7098 4908 7100
rect 4932 7098 4988 7100
rect 5012 7098 5068 7100
rect 5092 7098 5148 7100
rect 4852 7046 4898 7098
rect 4898 7046 4908 7098
rect 4932 7046 4962 7098
rect 4962 7046 4974 7098
rect 4974 7046 4988 7098
rect 5012 7046 5026 7098
rect 5026 7046 5038 7098
rect 5038 7046 5068 7098
rect 5092 7046 5102 7098
rect 5102 7046 5148 7098
rect 4852 7044 4908 7046
rect 4932 7044 4988 7046
rect 5012 7044 5068 7046
rect 5092 7044 5148 7046
rect 7449 7098 7505 7100
rect 7529 7098 7585 7100
rect 7609 7098 7665 7100
rect 7689 7098 7745 7100
rect 7449 7046 7495 7098
rect 7495 7046 7505 7098
rect 7529 7046 7559 7098
rect 7559 7046 7571 7098
rect 7571 7046 7585 7098
rect 7609 7046 7623 7098
rect 7623 7046 7635 7098
rect 7635 7046 7665 7098
rect 7689 7046 7699 7098
rect 7699 7046 7745 7098
rect 7449 7044 7505 7046
rect 7529 7044 7585 7046
rect 7609 7044 7665 7046
rect 7689 7044 7745 7046
rect 8114 6976 8170 7032
rect 3553 6554 3609 6556
rect 3633 6554 3689 6556
rect 3713 6554 3769 6556
rect 3793 6554 3849 6556
rect 3553 6502 3599 6554
rect 3599 6502 3609 6554
rect 3633 6502 3663 6554
rect 3663 6502 3675 6554
rect 3675 6502 3689 6554
rect 3713 6502 3727 6554
rect 3727 6502 3739 6554
rect 3739 6502 3769 6554
rect 3793 6502 3803 6554
rect 3803 6502 3849 6554
rect 3553 6500 3609 6502
rect 3633 6500 3689 6502
rect 3713 6500 3769 6502
rect 3793 6500 3849 6502
rect 6150 6554 6206 6556
rect 6230 6554 6286 6556
rect 6310 6554 6366 6556
rect 6390 6554 6446 6556
rect 6150 6502 6196 6554
rect 6196 6502 6206 6554
rect 6230 6502 6260 6554
rect 6260 6502 6272 6554
rect 6272 6502 6286 6554
rect 6310 6502 6324 6554
rect 6324 6502 6336 6554
rect 6336 6502 6366 6554
rect 6390 6502 6400 6554
rect 6400 6502 6446 6554
rect 6150 6500 6206 6502
rect 6230 6500 6286 6502
rect 6310 6500 6366 6502
rect 6390 6500 6446 6502
rect 8114 6432 8170 6488
rect 8114 6060 8116 6080
rect 8116 6060 8168 6080
rect 8168 6060 8170 6080
rect 2254 6010 2310 6012
rect 2334 6010 2390 6012
rect 2414 6010 2470 6012
rect 2494 6010 2550 6012
rect 2254 5958 2300 6010
rect 2300 5958 2310 6010
rect 2334 5958 2364 6010
rect 2364 5958 2376 6010
rect 2376 5958 2390 6010
rect 2414 5958 2428 6010
rect 2428 5958 2440 6010
rect 2440 5958 2470 6010
rect 2494 5958 2504 6010
rect 2504 5958 2550 6010
rect 2254 5956 2310 5958
rect 2334 5956 2390 5958
rect 2414 5956 2470 5958
rect 2494 5956 2550 5958
rect 4852 6010 4908 6012
rect 4932 6010 4988 6012
rect 5012 6010 5068 6012
rect 5092 6010 5148 6012
rect 4852 5958 4898 6010
rect 4898 5958 4908 6010
rect 4932 5958 4962 6010
rect 4962 5958 4974 6010
rect 4974 5958 4988 6010
rect 5012 5958 5026 6010
rect 5026 5958 5038 6010
rect 5038 5958 5068 6010
rect 5092 5958 5102 6010
rect 5102 5958 5148 6010
rect 4852 5956 4908 5958
rect 4932 5956 4988 5958
rect 5012 5956 5068 5958
rect 5092 5956 5148 5958
rect 8114 6024 8170 6060
rect 7449 6010 7505 6012
rect 7529 6010 7585 6012
rect 7609 6010 7665 6012
rect 7689 6010 7745 6012
rect 7449 5958 7495 6010
rect 7495 5958 7505 6010
rect 7529 5958 7559 6010
rect 7559 5958 7571 6010
rect 7571 5958 7585 6010
rect 7609 5958 7623 6010
rect 7623 5958 7635 6010
rect 7635 5958 7665 6010
rect 7689 5958 7699 6010
rect 7699 5958 7745 6010
rect 7449 5956 7505 5958
rect 7529 5956 7585 5958
rect 7609 5956 7665 5958
rect 7689 5956 7745 5958
rect 3553 5466 3609 5468
rect 3633 5466 3689 5468
rect 3713 5466 3769 5468
rect 3793 5466 3849 5468
rect 3553 5414 3599 5466
rect 3599 5414 3609 5466
rect 3633 5414 3663 5466
rect 3663 5414 3675 5466
rect 3675 5414 3689 5466
rect 3713 5414 3727 5466
rect 3727 5414 3739 5466
rect 3739 5414 3769 5466
rect 3793 5414 3803 5466
rect 3803 5414 3849 5466
rect 3553 5412 3609 5414
rect 3633 5412 3689 5414
rect 3713 5412 3769 5414
rect 3793 5412 3849 5414
rect 8114 5480 8170 5536
rect 6150 5466 6206 5468
rect 6230 5466 6286 5468
rect 6310 5466 6366 5468
rect 6390 5466 6446 5468
rect 6150 5414 6196 5466
rect 6196 5414 6206 5466
rect 6230 5414 6260 5466
rect 6260 5414 6272 5466
rect 6272 5414 6286 5466
rect 6310 5414 6324 5466
rect 6324 5414 6336 5466
rect 6336 5414 6366 5466
rect 6390 5414 6400 5466
rect 6400 5414 6446 5466
rect 6150 5412 6206 5414
rect 6230 5412 6286 5414
rect 6310 5412 6366 5414
rect 6390 5412 6446 5414
rect 8114 4972 8116 4992
rect 8116 4972 8168 4992
rect 8168 4972 8170 4992
rect 2254 4922 2310 4924
rect 2334 4922 2390 4924
rect 2414 4922 2470 4924
rect 2494 4922 2550 4924
rect 2254 4870 2300 4922
rect 2300 4870 2310 4922
rect 2334 4870 2364 4922
rect 2364 4870 2376 4922
rect 2376 4870 2390 4922
rect 2414 4870 2428 4922
rect 2428 4870 2440 4922
rect 2440 4870 2470 4922
rect 2494 4870 2504 4922
rect 2504 4870 2550 4922
rect 2254 4868 2310 4870
rect 2334 4868 2390 4870
rect 2414 4868 2470 4870
rect 2494 4868 2550 4870
rect 4852 4922 4908 4924
rect 4932 4922 4988 4924
rect 5012 4922 5068 4924
rect 5092 4922 5148 4924
rect 4852 4870 4898 4922
rect 4898 4870 4908 4922
rect 4932 4870 4962 4922
rect 4962 4870 4974 4922
rect 4974 4870 4988 4922
rect 5012 4870 5026 4922
rect 5026 4870 5038 4922
rect 5038 4870 5068 4922
rect 5092 4870 5102 4922
rect 5102 4870 5148 4922
rect 4852 4868 4908 4870
rect 4932 4868 4988 4870
rect 5012 4868 5068 4870
rect 5092 4868 5148 4870
rect 8114 4936 8170 4972
rect 7449 4922 7505 4924
rect 7529 4922 7585 4924
rect 7609 4922 7665 4924
rect 7689 4922 7745 4924
rect 7449 4870 7495 4922
rect 7495 4870 7505 4922
rect 7529 4870 7559 4922
rect 7559 4870 7571 4922
rect 7571 4870 7585 4922
rect 7609 4870 7623 4922
rect 7623 4870 7635 4922
rect 7635 4870 7665 4922
rect 7689 4870 7699 4922
rect 7699 4870 7745 4922
rect 7449 4868 7505 4870
rect 7529 4868 7585 4870
rect 7609 4868 7665 4870
rect 7689 4868 7745 4870
rect 8114 4428 8116 4448
rect 8116 4428 8168 4448
rect 8168 4428 8170 4448
rect 3553 4378 3609 4380
rect 3633 4378 3689 4380
rect 3713 4378 3769 4380
rect 3793 4378 3849 4380
rect 3553 4326 3599 4378
rect 3599 4326 3609 4378
rect 3633 4326 3663 4378
rect 3663 4326 3675 4378
rect 3675 4326 3689 4378
rect 3713 4326 3727 4378
rect 3727 4326 3739 4378
rect 3739 4326 3769 4378
rect 3793 4326 3803 4378
rect 3803 4326 3849 4378
rect 3553 4324 3609 4326
rect 3633 4324 3689 4326
rect 3713 4324 3769 4326
rect 3793 4324 3849 4326
rect 8114 4392 8170 4428
rect 6150 4378 6206 4380
rect 6230 4378 6286 4380
rect 6310 4378 6366 4380
rect 6390 4378 6446 4380
rect 6150 4326 6196 4378
rect 6196 4326 6206 4378
rect 6230 4326 6260 4378
rect 6260 4326 6272 4378
rect 6272 4326 6286 4378
rect 6310 4326 6324 4378
rect 6324 4326 6336 4378
rect 6336 4326 6366 4378
rect 6390 4326 6400 4378
rect 6400 4326 6446 4378
rect 6150 4324 6206 4326
rect 6230 4324 6286 4326
rect 6310 4324 6366 4326
rect 6390 4324 6446 4326
rect 7838 3884 7840 3904
rect 7840 3884 7892 3904
rect 7892 3884 7894 3904
rect 2254 3834 2310 3836
rect 2334 3834 2390 3836
rect 2414 3834 2470 3836
rect 2494 3834 2550 3836
rect 2254 3782 2300 3834
rect 2300 3782 2310 3834
rect 2334 3782 2364 3834
rect 2364 3782 2376 3834
rect 2376 3782 2390 3834
rect 2414 3782 2428 3834
rect 2428 3782 2440 3834
rect 2440 3782 2470 3834
rect 2494 3782 2504 3834
rect 2504 3782 2550 3834
rect 2254 3780 2310 3782
rect 2334 3780 2390 3782
rect 2414 3780 2470 3782
rect 2494 3780 2550 3782
rect 4852 3834 4908 3836
rect 4932 3834 4988 3836
rect 5012 3834 5068 3836
rect 5092 3834 5148 3836
rect 4852 3782 4898 3834
rect 4898 3782 4908 3834
rect 4932 3782 4962 3834
rect 4962 3782 4974 3834
rect 4974 3782 4988 3834
rect 5012 3782 5026 3834
rect 5026 3782 5038 3834
rect 5038 3782 5068 3834
rect 5092 3782 5102 3834
rect 5102 3782 5148 3834
rect 4852 3780 4908 3782
rect 4932 3780 4988 3782
rect 5012 3780 5068 3782
rect 5092 3780 5148 3782
rect 7838 3848 7894 3884
rect 7449 3834 7505 3836
rect 7529 3834 7585 3836
rect 7609 3834 7665 3836
rect 7689 3834 7745 3836
rect 7449 3782 7495 3834
rect 7495 3782 7505 3834
rect 7529 3782 7559 3834
rect 7559 3782 7571 3834
rect 7571 3782 7585 3834
rect 7609 3782 7623 3834
rect 7623 3782 7635 3834
rect 7635 3782 7665 3834
rect 7689 3782 7699 3834
rect 7699 3782 7745 3834
rect 7449 3780 7505 3782
rect 7529 3780 7585 3782
rect 7609 3780 7665 3782
rect 7689 3780 7745 3782
rect 3553 3290 3609 3292
rect 3633 3290 3689 3292
rect 3713 3290 3769 3292
rect 3793 3290 3849 3292
rect 3553 3238 3599 3290
rect 3599 3238 3609 3290
rect 3633 3238 3663 3290
rect 3663 3238 3675 3290
rect 3675 3238 3689 3290
rect 3713 3238 3727 3290
rect 3727 3238 3739 3290
rect 3739 3238 3769 3290
rect 3793 3238 3803 3290
rect 3803 3238 3849 3290
rect 3553 3236 3609 3238
rect 3633 3236 3689 3238
rect 3713 3236 3769 3238
rect 3793 3236 3849 3238
rect 7470 3304 7526 3360
rect 6150 3290 6206 3292
rect 6230 3290 6286 3292
rect 6310 3290 6366 3292
rect 6390 3290 6446 3292
rect 6150 3238 6196 3290
rect 6196 3238 6206 3290
rect 6230 3238 6260 3290
rect 6260 3238 6272 3290
rect 6272 3238 6286 3290
rect 6310 3238 6324 3290
rect 6324 3238 6336 3290
rect 6336 3238 6366 3290
rect 6390 3238 6400 3290
rect 6400 3238 6446 3290
rect 6150 3236 6206 3238
rect 6230 3236 6286 3238
rect 6310 3236 6366 3238
rect 6390 3236 6446 3238
rect 2254 2746 2310 2748
rect 2334 2746 2390 2748
rect 2414 2746 2470 2748
rect 2494 2746 2550 2748
rect 2254 2694 2300 2746
rect 2300 2694 2310 2746
rect 2334 2694 2364 2746
rect 2364 2694 2376 2746
rect 2376 2694 2390 2746
rect 2414 2694 2428 2746
rect 2428 2694 2440 2746
rect 2440 2694 2470 2746
rect 2494 2694 2504 2746
rect 2504 2694 2550 2746
rect 2254 2692 2310 2694
rect 2334 2692 2390 2694
rect 2414 2692 2470 2694
rect 2494 2692 2550 2694
rect 4852 2746 4908 2748
rect 4932 2746 4988 2748
rect 5012 2746 5068 2748
rect 5092 2746 5148 2748
rect 4852 2694 4898 2746
rect 4898 2694 4908 2746
rect 4932 2694 4962 2746
rect 4962 2694 4974 2746
rect 4974 2694 4988 2746
rect 5012 2694 5026 2746
rect 5026 2694 5038 2746
rect 5038 2694 5068 2746
rect 5092 2694 5102 2746
rect 5102 2694 5148 2746
rect 4852 2692 4908 2694
rect 4932 2692 4988 2694
rect 5012 2692 5068 2694
rect 5092 2692 5148 2694
rect 7449 2746 7505 2748
rect 7529 2746 7585 2748
rect 7609 2746 7665 2748
rect 7689 2746 7745 2748
rect 7449 2694 7495 2746
rect 7495 2694 7505 2746
rect 7529 2694 7559 2746
rect 7559 2694 7571 2746
rect 7571 2694 7585 2746
rect 7609 2694 7623 2746
rect 7623 2694 7635 2746
rect 7635 2694 7665 2746
rect 7689 2694 7699 2746
rect 7699 2694 7745 2746
rect 7449 2692 7505 2694
rect 7529 2692 7585 2694
rect 7609 2692 7665 2694
rect 7689 2692 7745 2694
rect 3553 2202 3609 2204
rect 3633 2202 3689 2204
rect 3713 2202 3769 2204
rect 3793 2202 3849 2204
rect 3553 2150 3599 2202
rect 3599 2150 3609 2202
rect 3633 2150 3663 2202
rect 3663 2150 3675 2202
rect 3675 2150 3689 2202
rect 3713 2150 3727 2202
rect 3727 2150 3739 2202
rect 3739 2150 3769 2202
rect 3793 2150 3803 2202
rect 3803 2150 3849 2202
rect 3553 2148 3609 2150
rect 3633 2148 3689 2150
rect 3713 2148 3769 2150
rect 3793 2148 3849 2150
rect 6150 2202 6206 2204
rect 6230 2202 6286 2204
rect 6310 2202 6366 2204
rect 6390 2202 6446 2204
rect 6150 2150 6196 2202
rect 6196 2150 6206 2202
rect 6230 2150 6260 2202
rect 6260 2150 6272 2202
rect 6272 2150 6286 2202
rect 6310 2150 6324 2202
rect 6324 2150 6336 2202
rect 6336 2150 6366 2202
rect 6390 2150 6400 2202
rect 6400 2150 6446 2202
rect 6150 2148 6206 2150
rect 6230 2148 6286 2150
rect 6310 2148 6366 2150
rect 6390 2148 6446 2150
rect 7838 2216 7894 2272
rect 7470 1128 7526 1184
rect 8114 2760 8170 2816
rect 8022 584 8078 640
rect 8206 1672 8262 1728
rect 8114 176 8170 232
<< metal3 >>
rect 6637 24714 6703 24717
rect 9200 24714 10000 24744
rect 6637 24712 10000 24714
rect 6637 24656 6642 24712
rect 6698 24656 10000 24712
rect 6637 24654 10000 24656
rect 6637 24651 6703 24654
rect 9200 24624 10000 24654
rect 7833 24170 7899 24173
rect 9200 24170 10000 24200
rect 7833 24168 10000 24170
rect 7833 24112 7838 24168
rect 7894 24112 10000 24168
rect 7833 24110 10000 24112
rect 7833 24107 7899 24110
rect 9200 24080 10000 24110
rect 6729 23626 6795 23629
rect 9200 23626 10000 23656
rect 6729 23624 10000 23626
rect 6729 23568 6734 23624
rect 6790 23568 10000 23624
rect 6729 23566 10000 23568
rect 6729 23563 6795 23566
rect 9200 23536 10000 23566
rect 6821 23082 6887 23085
rect 9200 23082 10000 23112
rect 6821 23080 10000 23082
rect 6821 23024 6826 23080
rect 6882 23024 10000 23080
rect 6821 23022 10000 23024
rect 6821 23019 6887 23022
rect 9200 22992 10000 23022
rect 8201 22538 8267 22541
rect 9200 22538 10000 22568
rect 8201 22536 10000 22538
rect 8201 22480 8206 22536
rect 8262 22480 10000 22536
rect 8201 22478 10000 22480
rect 8201 22475 8267 22478
rect 9200 22448 10000 22478
rect 2242 22336 2562 22337
rect 2242 22272 2250 22336
rect 2314 22272 2330 22336
rect 2394 22272 2410 22336
rect 2474 22272 2490 22336
rect 2554 22272 2562 22336
rect 2242 22271 2562 22272
rect 4840 22336 5160 22337
rect 4840 22272 4848 22336
rect 4912 22272 4928 22336
rect 4992 22272 5008 22336
rect 5072 22272 5088 22336
rect 5152 22272 5160 22336
rect 4840 22271 5160 22272
rect 7437 22336 7757 22337
rect 7437 22272 7445 22336
rect 7509 22272 7525 22336
rect 7589 22272 7605 22336
rect 7669 22272 7685 22336
rect 7749 22272 7757 22336
rect 7437 22271 7757 22272
rect 8109 21994 8175 21997
rect 9200 21994 10000 22024
rect 8109 21992 10000 21994
rect 8109 21936 8114 21992
rect 8170 21936 10000 21992
rect 8109 21934 10000 21936
rect 8109 21931 8175 21934
rect 9200 21904 10000 21934
rect 3541 21792 3861 21793
rect 3541 21728 3549 21792
rect 3613 21728 3629 21792
rect 3693 21728 3709 21792
rect 3773 21728 3789 21792
rect 3853 21728 3861 21792
rect 3541 21727 3861 21728
rect 6138 21792 6458 21793
rect 6138 21728 6146 21792
rect 6210 21728 6226 21792
rect 6290 21728 6306 21792
rect 6370 21728 6386 21792
rect 6450 21728 6458 21792
rect 6138 21727 6458 21728
rect 7465 21450 7531 21453
rect 9200 21450 10000 21480
rect 7465 21448 10000 21450
rect 7465 21392 7470 21448
rect 7526 21392 10000 21448
rect 7465 21390 10000 21392
rect 7465 21387 7531 21390
rect 9200 21360 10000 21390
rect 2242 21248 2562 21249
rect 2242 21184 2250 21248
rect 2314 21184 2330 21248
rect 2394 21184 2410 21248
rect 2474 21184 2490 21248
rect 2554 21184 2562 21248
rect 2242 21183 2562 21184
rect 4840 21248 5160 21249
rect 4840 21184 4848 21248
rect 4912 21184 4928 21248
rect 4992 21184 5008 21248
rect 5072 21184 5088 21248
rect 5152 21184 5160 21248
rect 4840 21183 5160 21184
rect 7437 21248 7757 21249
rect 7437 21184 7445 21248
rect 7509 21184 7525 21248
rect 7589 21184 7605 21248
rect 7669 21184 7685 21248
rect 7749 21184 7757 21248
rect 7437 21183 7757 21184
rect 8109 20906 8175 20909
rect 9200 20906 10000 20936
rect 8109 20904 10000 20906
rect 8109 20848 8114 20904
rect 8170 20848 10000 20904
rect 8109 20846 10000 20848
rect 8109 20843 8175 20846
rect 9200 20816 10000 20846
rect 3541 20704 3861 20705
rect 3541 20640 3549 20704
rect 3613 20640 3629 20704
rect 3693 20640 3709 20704
rect 3773 20640 3789 20704
rect 3853 20640 3861 20704
rect 3541 20639 3861 20640
rect 6138 20704 6458 20705
rect 6138 20640 6146 20704
rect 6210 20640 6226 20704
rect 6290 20640 6306 20704
rect 6370 20640 6386 20704
rect 6450 20640 6458 20704
rect 6138 20639 6458 20640
rect 8109 20362 8175 20365
rect 9200 20362 10000 20392
rect 8109 20360 10000 20362
rect 8109 20304 8114 20360
rect 8170 20304 10000 20360
rect 8109 20302 10000 20304
rect 8109 20299 8175 20302
rect 9200 20272 10000 20302
rect 2242 20160 2562 20161
rect 2242 20096 2250 20160
rect 2314 20096 2330 20160
rect 2394 20096 2410 20160
rect 2474 20096 2490 20160
rect 2554 20096 2562 20160
rect 2242 20095 2562 20096
rect 4840 20160 5160 20161
rect 4840 20096 4848 20160
rect 4912 20096 4928 20160
rect 4992 20096 5008 20160
rect 5072 20096 5088 20160
rect 5152 20096 5160 20160
rect 4840 20095 5160 20096
rect 7437 20160 7757 20161
rect 7437 20096 7445 20160
rect 7509 20096 7525 20160
rect 7589 20096 7605 20160
rect 7669 20096 7685 20160
rect 7749 20096 7757 20160
rect 7437 20095 7757 20096
rect 8109 19818 8175 19821
rect 9200 19818 10000 19848
rect 8109 19816 10000 19818
rect 8109 19760 8114 19816
rect 8170 19760 10000 19816
rect 8109 19758 10000 19760
rect 8109 19755 8175 19758
rect 9200 19728 10000 19758
rect 3541 19616 3861 19617
rect 3541 19552 3549 19616
rect 3613 19552 3629 19616
rect 3693 19552 3709 19616
rect 3773 19552 3789 19616
rect 3853 19552 3861 19616
rect 3541 19551 3861 19552
rect 6138 19616 6458 19617
rect 6138 19552 6146 19616
rect 6210 19552 6226 19616
rect 6290 19552 6306 19616
rect 6370 19552 6386 19616
rect 6450 19552 6458 19616
rect 6138 19551 6458 19552
rect 7465 19274 7531 19277
rect 9200 19274 10000 19304
rect 7465 19272 10000 19274
rect 7465 19216 7470 19272
rect 7526 19216 10000 19272
rect 7465 19214 10000 19216
rect 7465 19211 7531 19214
rect 9200 19184 10000 19214
rect 2242 19072 2562 19073
rect 2242 19008 2250 19072
rect 2314 19008 2330 19072
rect 2394 19008 2410 19072
rect 2474 19008 2490 19072
rect 2554 19008 2562 19072
rect 2242 19007 2562 19008
rect 4840 19072 5160 19073
rect 4840 19008 4848 19072
rect 4912 19008 4928 19072
rect 4992 19008 5008 19072
rect 5072 19008 5088 19072
rect 5152 19008 5160 19072
rect 4840 19007 5160 19008
rect 7437 19072 7757 19073
rect 7437 19008 7445 19072
rect 7509 19008 7525 19072
rect 7589 19008 7605 19072
rect 7669 19008 7685 19072
rect 7749 19008 7757 19072
rect 7437 19007 7757 19008
rect 8109 18866 8175 18869
rect 9200 18866 10000 18896
rect 8109 18864 10000 18866
rect 8109 18808 8114 18864
rect 8170 18808 10000 18864
rect 8109 18806 10000 18808
rect 8109 18803 8175 18806
rect 9200 18776 10000 18806
rect 3541 18528 3861 18529
rect 3541 18464 3549 18528
rect 3613 18464 3629 18528
rect 3693 18464 3709 18528
rect 3773 18464 3789 18528
rect 3853 18464 3861 18528
rect 3541 18463 3861 18464
rect 6138 18528 6458 18529
rect 6138 18464 6146 18528
rect 6210 18464 6226 18528
rect 6290 18464 6306 18528
rect 6370 18464 6386 18528
rect 6450 18464 6458 18528
rect 6138 18463 6458 18464
rect 8109 18322 8175 18325
rect 9200 18322 10000 18352
rect 8109 18320 10000 18322
rect 8109 18264 8114 18320
rect 8170 18264 10000 18320
rect 8109 18262 10000 18264
rect 8109 18259 8175 18262
rect 9200 18232 10000 18262
rect 2242 17984 2562 17985
rect 2242 17920 2250 17984
rect 2314 17920 2330 17984
rect 2394 17920 2410 17984
rect 2474 17920 2490 17984
rect 2554 17920 2562 17984
rect 2242 17919 2562 17920
rect 4840 17984 5160 17985
rect 4840 17920 4848 17984
rect 4912 17920 4928 17984
rect 4992 17920 5008 17984
rect 5072 17920 5088 17984
rect 5152 17920 5160 17984
rect 4840 17919 5160 17920
rect 7437 17984 7757 17985
rect 7437 17920 7445 17984
rect 7509 17920 7525 17984
rect 7589 17920 7605 17984
rect 7669 17920 7685 17984
rect 7749 17920 7757 17984
rect 7437 17919 7757 17920
rect 8109 17778 8175 17781
rect 9200 17778 10000 17808
rect 8109 17776 10000 17778
rect 8109 17720 8114 17776
rect 8170 17720 10000 17776
rect 8109 17718 10000 17720
rect 8109 17715 8175 17718
rect 9200 17688 10000 17718
rect 3541 17440 3861 17441
rect 3541 17376 3549 17440
rect 3613 17376 3629 17440
rect 3693 17376 3709 17440
rect 3773 17376 3789 17440
rect 3853 17376 3861 17440
rect 3541 17375 3861 17376
rect 6138 17440 6458 17441
rect 6138 17376 6146 17440
rect 6210 17376 6226 17440
rect 6290 17376 6306 17440
rect 6370 17376 6386 17440
rect 6450 17376 6458 17440
rect 6138 17375 6458 17376
rect 8109 17234 8175 17237
rect 9200 17234 10000 17264
rect 8109 17232 10000 17234
rect 8109 17176 8114 17232
rect 8170 17176 10000 17232
rect 8109 17174 10000 17176
rect 8109 17171 8175 17174
rect 9200 17144 10000 17174
rect 2242 16896 2562 16897
rect 2242 16832 2250 16896
rect 2314 16832 2330 16896
rect 2394 16832 2410 16896
rect 2474 16832 2490 16896
rect 2554 16832 2562 16896
rect 2242 16831 2562 16832
rect 4840 16896 5160 16897
rect 4840 16832 4848 16896
rect 4912 16832 4928 16896
rect 4992 16832 5008 16896
rect 5072 16832 5088 16896
rect 5152 16832 5160 16896
rect 4840 16831 5160 16832
rect 7437 16896 7757 16897
rect 7437 16832 7445 16896
rect 7509 16832 7525 16896
rect 7589 16832 7605 16896
rect 7669 16832 7685 16896
rect 7749 16832 7757 16896
rect 7437 16831 7757 16832
rect 8201 16690 8267 16693
rect 9200 16690 10000 16720
rect 8201 16688 10000 16690
rect 8201 16632 8206 16688
rect 8262 16632 10000 16688
rect 8201 16630 10000 16632
rect 8201 16627 8267 16630
rect 9200 16600 10000 16630
rect 3541 16352 3861 16353
rect 3541 16288 3549 16352
rect 3613 16288 3629 16352
rect 3693 16288 3709 16352
rect 3773 16288 3789 16352
rect 3853 16288 3861 16352
rect 3541 16287 3861 16288
rect 6138 16352 6458 16353
rect 6138 16288 6146 16352
rect 6210 16288 6226 16352
rect 6290 16288 6306 16352
rect 6370 16288 6386 16352
rect 6450 16288 6458 16352
rect 6138 16287 6458 16288
rect 8109 16146 8175 16149
rect 9200 16146 10000 16176
rect 8109 16144 10000 16146
rect 8109 16088 8114 16144
rect 8170 16088 10000 16144
rect 8109 16086 10000 16088
rect 8109 16083 8175 16086
rect 9200 16056 10000 16086
rect 2242 15808 2562 15809
rect 2242 15744 2250 15808
rect 2314 15744 2330 15808
rect 2394 15744 2410 15808
rect 2474 15744 2490 15808
rect 2554 15744 2562 15808
rect 2242 15743 2562 15744
rect 4840 15808 5160 15809
rect 4840 15744 4848 15808
rect 4912 15744 4928 15808
rect 4992 15744 5008 15808
rect 5072 15744 5088 15808
rect 5152 15744 5160 15808
rect 4840 15743 5160 15744
rect 7437 15808 7757 15809
rect 7437 15744 7445 15808
rect 7509 15744 7525 15808
rect 7589 15744 7605 15808
rect 7669 15744 7685 15808
rect 7749 15744 7757 15808
rect 7437 15743 7757 15744
rect 8109 15602 8175 15605
rect 9200 15602 10000 15632
rect 8109 15600 10000 15602
rect 8109 15544 8114 15600
rect 8170 15544 10000 15600
rect 8109 15542 10000 15544
rect 8109 15539 8175 15542
rect 9200 15512 10000 15542
rect 3541 15264 3861 15265
rect 3541 15200 3549 15264
rect 3613 15200 3629 15264
rect 3693 15200 3709 15264
rect 3773 15200 3789 15264
rect 3853 15200 3861 15264
rect 3541 15199 3861 15200
rect 6138 15264 6458 15265
rect 6138 15200 6146 15264
rect 6210 15200 6226 15264
rect 6290 15200 6306 15264
rect 6370 15200 6386 15264
rect 6450 15200 6458 15264
rect 6138 15199 6458 15200
rect 8109 15058 8175 15061
rect 9200 15058 10000 15088
rect 8109 15056 10000 15058
rect 8109 15000 8114 15056
rect 8170 15000 10000 15056
rect 8109 14998 10000 15000
rect 8109 14995 8175 14998
rect 9200 14968 10000 14998
rect 2242 14720 2562 14721
rect 2242 14656 2250 14720
rect 2314 14656 2330 14720
rect 2394 14656 2410 14720
rect 2474 14656 2490 14720
rect 2554 14656 2562 14720
rect 2242 14655 2562 14656
rect 4840 14720 5160 14721
rect 4840 14656 4848 14720
rect 4912 14656 4928 14720
rect 4992 14656 5008 14720
rect 5072 14656 5088 14720
rect 5152 14656 5160 14720
rect 4840 14655 5160 14656
rect 7437 14720 7757 14721
rect 7437 14656 7445 14720
rect 7509 14656 7525 14720
rect 7589 14656 7605 14720
rect 7669 14656 7685 14720
rect 7749 14656 7757 14720
rect 7437 14655 7757 14656
rect 8109 14514 8175 14517
rect 9200 14514 10000 14544
rect 8109 14512 10000 14514
rect 8109 14456 8114 14512
rect 8170 14456 10000 14512
rect 8109 14454 10000 14456
rect 8109 14451 8175 14454
rect 9200 14424 10000 14454
rect 3541 14176 3861 14177
rect 3541 14112 3549 14176
rect 3613 14112 3629 14176
rect 3693 14112 3709 14176
rect 3773 14112 3789 14176
rect 3853 14112 3861 14176
rect 3541 14111 3861 14112
rect 6138 14176 6458 14177
rect 6138 14112 6146 14176
rect 6210 14112 6226 14176
rect 6290 14112 6306 14176
rect 6370 14112 6386 14176
rect 6450 14112 6458 14176
rect 6138 14111 6458 14112
rect 8109 13970 8175 13973
rect 9200 13970 10000 14000
rect 8109 13968 10000 13970
rect 8109 13912 8114 13968
rect 8170 13912 10000 13968
rect 8109 13910 10000 13912
rect 8109 13907 8175 13910
rect 9200 13880 10000 13910
rect 2242 13632 2562 13633
rect 2242 13568 2250 13632
rect 2314 13568 2330 13632
rect 2394 13568 2410 13632
rect 2474 13568 2490 13632
rect 2554 13568 2562 13632
rect 2242 13567 2562 13568
rect 4840 13632 5160 13633
rect 4840 13568 4848 13632
rect 4912 13568 4928 13632
rect 4992 13568 5008 13632
rect 5072 13568 5088 13632
rect 5152 13568 5160 13632
rect 4840 13567 5160 13568
rect 7437 13632 7757 13633
rect 7437 13568 7445 13632
rect 7509 13568 7525 13632
rect 7589 13568 7605 13632
rect 7669 13568 7685 13632
rect 7749 13568 7757 13632
rect 7437 13567 7757 13568
rect 8109 13426 8175 13429
rect 9200 13426 10000 13456
rect 8109 13424 10000 13426
rect 8109 13368 8114 13424
rect 8170 13368 10000 13424
rect 8109 13366 10000 13368
rect 8109 13363 8175 13366
rect 9200 13336 10000 13366
rect 3541 13088 3861 13089
rect 3541 13024 3549 13088
rect 3613 13024 3629 13088
rect 3693 13024 3709 13088
rect 3773 13024 3789 13088
rect 3853 13024 3861 13088
rect 3541 13023 3861 13024
rect 6138 13088 6458 13089
rect 6138 13024 6146 13088
rect 6210 13024 6226 13088
rect 6290 13024 6306 13088
rect 6370 13024 6386 13088
rect 6450 13024 6458 13088
rect 6138 13023 6458 13024
rect 8109 12882 8175 12885
rect 9200 12882 10000 12912
rect 8109 12880 10000 12882
rect 8109 12824 8114 12880
rect 8170 12824 10000 12880
rect 8109 12822 10000 12824
rect 8109 12819 8175 12822
rect 9200 12792 10000 12822
rect 2242 12544 2562 12545
rect 2242 12480 2250 12544
rect 2314 12480 2330 12544
rect 2394 12480 2410 12544
rect 2474 12480 2490 12544
rect 2554 12480 2562 12544
rect 2242 12479 2562 12480
rect 4840 12544 5160 12545
rect 4840 12480 4848 12544
rect 4912 12480 4928 12544
rect 4992 12480 5008 12544
rect 5072 12480 5088 12544
rect 5152 12480 5160 12544
rect 4840 12479 5160 12480
rect 7437 12544 7757 12545
rect 7437 12480 7445 12544
rect 7509 12480 7525 12544
rect 7589 12480 7605 12544
rect 7669 12480 7685 12544
rect 7749 12480 7757 12544
rect 7437 12479 7757 12480
rect 8109 12474 8175 12477
rect 9200 12474 10000 12504
rect 8109 12472 10000 12474
rect 8109 12416 8114 12472
rect 8170 12416 10000 12472
rect 8109 12414 10000 12416
rect 8109 12411 8175 12414
rect 9200 12384 10000 12414
rect 3541 12000 3861 12001
rect 3541 11936 3549 12000
rect 3613 11936 3629 12000
rect 3693 11936 3709 12000
rect 3773 11936 3789 12000
rect 3853 11936 3861 12000
rect 3541 11935 3861 11936
rect 6138 12000 6458 12001
rect 6138 11936 6146 12000
rect 6210 11936 6226 12000
rect 6290 11936 6306 12000
rect 6370 11936 6386 12000
rect 6450 11936 6458 12000
rect 6138 11935 6458 11936
rect 8109 11930 8175 11933
rect 9200 11930 10000 11960
rect 8109 11928 10000 11930
rect 8109 11872 8114 11928
rect 8170 11872 10000 11928
rect 8109 11870 10000 11872
rect 8109 11867 8175 11870
rect 9200 11840 10000 11870
rect 2242 11456 2562 11457
rect 2242 11392 2250 11456
rect 2314 11392 2330 11456
rect 2394 11392 2410 11456
rect 2474 11392 2490 11456
rect 2554 11392 2562 11456
rect 2242 11391 2562 11392
rect 4840 11456 5160 11457
rect 4840 11392 4848 11456
rect 4912 11392 4928 11456
rect 4992 11392 5008 11456
rect 5072 11392 5088 11456
rect 5152 11392 5160 11456
rect 4840 11391 5160 11392
rect 7437 11456 7757 11457
rect 7437 11392 7445 11456
rect 7509 11392 7525 11456
rect 7589 11392 7605 11456
rect 7669 11392 7685 11456
rect 7749 11392 7757 11456
rect 7437 11391 7757 11392
rect 8109 11386 8175 11389
rect 9200 11386 10000 11416
rect 8109 11384 10000 11386
rect 8109 11328 8114 11384
rect 8170 11328 10000 11384
rect 8109 11326 10000 11328
rect 8109 11323 8175 11326
rect 9200 11296 10000 11326
rect 3541 10912 3861 10913
rect 3541 10848 3549 10912
rect 3613 10848 3629 10912
rect 3693 10848 3709 10912
rect 3773 10848 3789 10912
rect 3853 10848 3861 10912
rect 3541 10847 3861 10848
rect 6138 10912 6458 10913
rect 6138 10848 6146 10912
rect 6210 10848 6226 10912
rect 6290 10848 6306 10912
rect 6370 10848 6386 10912
rect 6450 10848 6458 10912
rect 6138 10847 6458 10848
rect 8109 10842 8175 10845
rect 9200 10842 10000 10872
rect 8109 10840 10000 10842
rect 8109 10784 8114 10840
rect 8170 10784 10000 10840
rect 8109 10782 10000 10784
rect 8109 10779 8175 10782
rect 9200 10752 10000 10782
rect 2242 10368 2562 10369
rect 2242 10304 2250 10368
rect 2314 10304 2330 10368
rect 2394 10304 2410 10368
rect 2474 10304 2490 10368
rect 2554 10304 2562 10368
rect 2242 10303 2562 10304
rect 4840 10368 5160 10369
rect 4840 10304 4848 10368
rect 4912 10304 4928 10368
rect 4992 10304 5008 10368
rect 5072 10304 5088 10368
rect 5152 10304 5160 10368
rect 4840 10303 5160 10304
rect 7437 10368 7757 10369
rect 7437 10304 7445 10368
rect 7509 10304 7525 10368
rect 7589 10304 7605 10368
rect 7669 10304 7685 10368
rect 7749 10304 7757 10368
rect 7437 10303 7757 10304
rect 8109 10298 8175 10301
rect 9200 10298 10000 10328
rect 8109 10296 10000 10298
rect 8109 10240 8114 10296
rect 8170 10240 10000 10296
rect 8109 10238 10000 10240
rect 8109 10235 8175 10238
rect 9200 10208 10000 10238
rect 3541 9824 3861 9825
rect 3541 9760 3549 9824
rect 3613 9760 3629 9824
rect 3693 9760 3709 9824
rect 3773 9760 3789 9824
rect 3853 9760 3861 9824
rect 3541 9759 3861 9760
rect 6138 9824 6458 9825
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 6138 9759 6458 9760
rect 8109 9754 8175 9757
rect 9200 9754 10000 9784
rect 8109 9752 10000 9754
rect 8109 9696 8114 9752
rect 8170 9696 10000 9752
rect 8109 9694 10000 9696
rect 8109 9691 8175 9694
rect 9200 9664 10000 9694
rect 2242 9280 2562 9281
rect 2242 9216 2250 9280
rect 2314 9216 2330 9280
rect 2394 9216 2410 9280
rect 2474 9216 2490 9280
rect 2554 9216 2562 9280
rect 2242 9215 2562 9216
rect 4840 9280 5160 9281
rect 4840 9216 4848 9280
rect 4912 9216 4928 9280
rect 4992 9216 5008 9280
rect 5072 9216 5088 9280
rect 5152 9216 5160 9280
rect 4840 9215 5160 9216
rect 7437 9280 7757 9281
rect 7437 9216 7445 9280
rect 7509 9216 7525 9280
rect 7589 9216 7605 9280
rect 7669 9216 7685 9280
rect 7749 9216 7757 9280
rect 7437 9215 7757 9216
rect 8109 9210 8175 9213
rect 9200 9210 10000 9240
rect 8109 9208 10000 9210
rect 8109 9152 8114 9208
rect 8170 9152 10000 9208
rect 8109 9150 10000 9152
rect 8109 9147 8175 9150
rect 9200 9120 10000 9150
rect 3541 8736 3861 8737
rect 3541 8672 3549 8736
rect 3613 8672 3629 8736
rect 3693 8672 3709 8736
rect 3773 8672 3789 8736
rect 3853 8672 3861 8736
rect 3541 8671 3861 8672
rect 6138 8736 6458 8737
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 6138 8671 6458 8672
rect 8109 8666 8175 8669
rect 9200 8666 10000 8696
rect 8109 8664 10000 8666
rect 8109 8608 8114 8664
rect 8170 8608 10000 8664
rect 8109 8606 10000 8608
rect 8109 8603 8175 8606
rect 9200 8576 10000 8606
rect 2242 8192 2562 8193
rect 2242 8128 2250 8192
rect 2314 8128 2330 8192
rect 2394 8128 2410 8192
rect 2474 8128 2490 8192
rect 2554 8128 2562 8192
rect 2242 8127 2562 8128
rect 4840 8192 5160 8193
rect 4840 8128 4848 8192
rect 4912 8128 4928 8192
rect 4992 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5160 8192
rect 4840 8127 5160 8128
rect 7437 8192 7757 8193
rect 7437 8128 7445 8192
rect 7509 8128 7525 8192
rect 7589 8128 7605 8192
rect 7669 8128 7685 8192
rect 7749 8128 7757 8192
rect 7437 8127 7757 8128
rect 8109 8122 8175 8125
rect 9200 8122 10000 8152
rect 8109 8120 10000 8122
rect 8109 8064 8114 8120
rect 8170 8064 10000 8120
rect 8109 8062 10000 8064
rect 8109 8059 8175 8062
rect 9200 8032 10000 8062
rect 3541 7648 3861 7649
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 7583 3861 7584
rect 6138 7648 6458 7649
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 7583 6458 7584
rect 8109 7578 8175 7581
rect 9200 7578 10000 7608
rect 8109 7576 10000 7578
rect 8109 7520 8114 7576
rect 8170 7520 10000 7576
rect 8109 7518 10000 7520
rect 8109 7515 8175 7518
rect 9200 7488 10000 7518
rect 2242 7104 2562 7105
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2562 7104
rect 2242 7039 2562 7040
rect 4840 7104 5160 7105
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 7039 5160 7040
rect 7437 7104 7757 7105
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 7039 7757 7040
rect 8109 7034 8175 7037
rect 9200 7034 10000 7064
rect 8109 7032 10000 7034
rect 8109 6976 8114 7032
rect 8170 6976 10000 7032
rect 8109 6974 10000 6976
rect 8109 6971 8175 6974
rect 9200 6944 10000 6974
rect 3541 6560 3861 6561
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 6495 3861 6496
rect 6138 6560 6458 6561
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 6138 6495 6458 6496
rect 8109 6490 8175 6493
rect 9200 6490 10000 6520
rect 8109 6488 10000 6490
rect 8109 6432 8114 6488
rect 8170 6432 10000 6488
rect 8109 6430 10000 6432
rect 8109 6427 8175 6430
rect 9200 6400 10000 6430
rect 8109 6082 8175 6085
rect 9200 6082 10000 6112
rect 8109 6080 10000 6082
rect 8109 6024 8114 6080
rect 8170 6024 10000 6080
rect 8109 6022 10000 6024
rect 8109 6019 8175 6022
rect 2242 6016 2562 6017
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2562 6016
rect 2242 5951 2562 5952
rect 4840 6016 5160 6017
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 5951 5160 5952
rect 7437 6016 7757 6017
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 9200 5992 10000 6022
rect 7437 5951 7757 5952
rect 8109 5538 8175 5541
rect 9200 5538 10000 5568
rect 8109 5536 10000 5538
rect 8109 5480 8114 5536
rect 8170 5480 10000 5536
rect 8109 5478 10000 5480
rect 8109 5475 8175 5478
rect 3541 5472 3861 5473
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 5407 3861 5408
rect 6138 5472 6458 5473
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 9200 5448 10000 5478
rect 6138 5407 6458 5408
rect 8109 4994 8175 4997
rect 9200 4994 10000 5024
rect 8109 4992 10000 4994
rect 8109 4936 8114 4992
rect 8170 4936 10000 4992
rect 8109 4934 10000 4936
rect 8109 4931 8175 4934
rect 2242 4928 2562 4929
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2562 4928
rect 2242 4863 2562 4864
rect 4840 4928 5160 4929
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 4863 5160 4864
rect 7437 4928 7757 4929
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 9200 4904 10000 4934
rect 7437 4863 7757 4864
rect 8109 4450 8175 4453
rect 9200 4450 10000 4480
rect 8109 4448 10000 4450
rect 8109 4392 8114 4448
rect 8170 4392 10000 4448
rect 8109 4390 10000 4392
rect 8109 4387 8175 4390
rect 3541 4384 3861 4385
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 4319 3861 4320
rect 6138 4384 6458 4385
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 9200 4360 10000 4390
rect 6138 4319 6458 4320
rect 7833 3906 7899 3909
rect 9200 3906 10000 3936
rect 7833 3904 10000 3906
rect 7833 3848 7838 3904
rect 7894 3848 10000 3904
rect 7833 3846 10000 3848
rect 7833 3843 7899 3846
rect 2242 3840 2562 3841
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2562 3840
rect 2242 3775 2562 3776
rect 4840 3840 5160 3841
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 3775 5160 3776
rect 7437 3840 7757 3841
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 9200 3816 10000 3846
rect 7437 3775 7757 3776
rect 7465 3362 7531 3365
rect 9200 3362 10000 3392
rect 7465 3360 10000 3362
rect 7465 3304 7470 3360
rect 7526 3304 10000 3360
rect 7465 3302 10000 3304
rect 7465 3299 7531 3302
rect 3541 3296 3861 3297
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 3231 3861 3232
rect 6138 3296 6458 3297
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 9200 3272 10000 3302
rect 6138 3231 6458 3232
rect 8109 2818 8175 2821
rect 9200 2818 10000 2848
rect 8109 2816 10000 2818
rect 8109 2760 8114 2816
rect 8170 2760 10000 2816
rect 8109 2758 10000 2760
rect 8109 2755 8175 2758
rect 2242 2752 2562 2753
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2562 2752
rect 2242 2687 2562 2688
rect 4840 2752 5160 2753
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2687 5160 2688
rect 7437 2752 7757 2753
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 9200 2728 10000 2758
rect 7437 2687 7757 2688
rect 7833 2274 7899 2277
rect 9200 2274 10000 2304
rect 7833 2272 10000 2274
rect 7833 2216 7838 2272
rect 7894 2216 10000 2272
rect 7833 2214 10000 2216
rect 7833 2211 7899 2214
rect 3541 2208 3861 2209
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2143 3861 2144
rect 6138 2208 6458 2209
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 9200 2184 10000 2214
rect 6138 2143 6458 2144
rect 8201 1730 8267 1733
rect 9200 1730 10000 1760
rect 8201 1728 10000 1730
rect 8201 1672 8206 1728
rect 8262 1672 10000 1728
rect 8201 1670 10000 1672
rect 8201 1667 8267 1670
rect 9200 1640 10000 1670
rect 7465 1186 7531 1189
rect 9200 1186 10000 1216
rect 7465 1184 10000 1186
rect 7465 1128 7470 1184
rect 7526 1128 10000 1184
rect 7465 1126 10000 1128
rect 7465 1123 7531 1126
rect 9200 1096 10000 1126
rect 8017 642 8083 645
rect 9200 642 10000 672
rect 8017 640 10000 642
rect 8017 584 8022 640
rect 8078 584 10000 640
rect 8017 582 10000 584
rect 8017 579 8083 582
rect 9200 552 10000 582
rect 8109 234 8175 237
rect 9200 234 10000 264
rect 8109 232 10000 234
rect 8109 176 8114 232
rect 8170 176 10000 232
rect 8109 174 10000 176
rect 8109 171 8175 174
rect 9200 144 10000 174
<< via3 >>
rect 2250 22332 2314 22336
rect 2250 22276 2254 22332
rect 2254 22276 2310 22332
rect 2310 22276 2314 22332
rect 2250 22272 2314 22276
rect 2330 22332 2394 22336
rect 2330 22276 2334 22332
rect 2334 22276 2390 22332
rect 2390 22276 2394 22332
rect 2330 22272 2394 22276
rect 2410 22332 2474 22336
rect 2410 22276 2414 22332
rect 2414 22276 2470 22332
rect 2470 22276 2474 22332
rect 2410 22272 2474 22276
rect 2490 22332 2554 22336
rect 2490 22276 2494 22332
rect 2494 22276 2550 22332
rect 2550 22276 2554 22332
rect 2490 22272 2554 22276
rect 4848 22332 4912 22336
rect 4848 22276 4852 22332
rect 4852 22276 4908 22332
rect 4908 22276 4912 22332
rect 4848 22272 4912 22276
rect 4928 22332 4992 22336
rect 4928 22276 4932 22332
rect 4932 22276 4988 22332
rect 4988 22276 4992 22332
rect 4928 22272 4992 22276
rect 5008 22332 5072 22336
rect 5008 22276 5012 22332
rect 5012 22276 5068 22332
rect 5068 22276 5072 22332
rect 5008 22272 5072 22276
rect 5088 22332 5152 22336
rect 5088 22276 5092 22332
rect 5092 22276 5148 22332
rect 5148 22276 5152 22332
rect 5088 22272 5152 22276
rect 7445 22332 7509 22336
rect 7445 22276 7449 22332
rect 7449 22276 7505 22332
rect 7505 22276 7509 22332
rect 7445 22272 7509 22276
rect 7525 22332 7589 22336
rect 7525 22276 7529 22332
rect 7529 22276 7585 22332
rect 7585 22276 7589 22332
rect 7525 22272 7589 22276
rect 7605 22332 7669 22336
rect 7605 22276 7609 22332
rect 7609 22276 7665 22332
rect 7665 22276 7669 22332
rect 7605 22272 7669 22276
rect 7685 22332 7749 22336
rect 7685 22276 7689 22332
rect 7689 22276 7745 22332
rect 7745 22276 7749 22332
rect 7685 22272 7749 22276
rect 3549 21788 3613 21792
rect 3549 21732 3553 21788
rect 3553 21732 3609 21788
rect 3609 21732 3613 21788
rect 3549 21728 3613 21732
rect 3629 21788 3693 21792
rect 3629 21732 3633 21788
rect 3633 21732 3689 21788
rect 3689 21732 3693 21788
rect 3629 21728 3693 21732
rect 3709 21788 3773 21792
rect 3709 21732 3713 21788
rect 3713 21732 3769 21788
rect 3769 21732 3773 21788
rect 3709 21728 3773 21732
rect 3789 21788 3853 21792
rect 3789 21732 3793 21788
rect 3793 21732 3849 21788
rect 3849 21732 3853 21788
rect 3789 21728 3853 21732
rect 6146 21788 6210 21792
rect 6146 21732 6150 21788
rect 6150 21732 6206 21788
rect 6206 21732 6210 21788
rect 6146 21728 6210 21732
rect 6226 21788 6290 21792
rect 6226 21732 6230 21788
rect 6230 21732 6286 21788
rect 6286 21732 6290 21788
rect 6226 21728 6290 21732
rect 6306 21788 6370 21792
rect 6306 21732 6310 21788
rect 6310 21732 6366 21788
rect 6366 21732 6370 21788
rect 6306 21728 6370 21732
rect 6386 21788 6450 21792
rect 6386 21732 6390 21788
rect 6390 21732 6446 21788
rect 6446 21732 6450 21788
rect 6386 21728 6450 21732
rect 2250 21244 2314 21248
rect 2250 21188 2254 21244
rect 2254 21188 2310 21244
rect 2310 21188 2314 21244
rect 2250 21184 2314 21188
rect 2330 21244 2394 21248
rect 2330 21188 2334 21244
rect 2334 21188 2390 21244
rect 2390 21188 2394 21244
rect 2330 21184 2394 21188
rect 2410 21244 2474 21248
rect 2410 21188 2414 21244
rect 2414 21188 2470 21244
rect 2470 21188 2474 21244
rect 2410 21184 2474 21188
rect 2490 21244 2554 21248
rect 2490 21188 2494 21244
rect 2494 21188 2550 21244
rect 2550 21188 2554 21244
rect 2490 21184 2554 21188
rect 4848 21244 4912 21248
rect 4848 21188 4852 21244
rect 4852 21188 4908 21244
rect 4908 21188 4912 21244
rect 4848 21184 4912 21188
rect 4928 21244 4992 21248
rect 4928 21188 4932 21244
rect 4932 21188 4988 21244
rect 4988 21188 4992 21244
rect 4928 21184 4992 21188
rect 5008 21244 5072 21248
rect 5008 21188 5012 21244
rect 5012 21188 5068 21244
rect 5068 21188 5072 21244
rect 5008 21184 5072 21188
rect 5088 21244 5152 21248
rect 5088 21188 5092 21244
rect 5092 21188 5148 21244
rect 5148 21188 5152 21244
rect 5088 21184 5152 21188
rect 7445 21244 7509 21248
rect 7445 21188 7449 21244
rect 7449 21188 7505 21244
rect 7505 21188 7509 21244
rect 7445 21184 7509 21188
rect 7525 21244 7589 21248
rect 7525 21188 7529 21244
rect 7529 21188 7585 21244
rect 7585 21188 7589 21244
rect 7525 21184 7589 21188
rect 7605 21244 7669 21248
rect 7605 21188 7609 21244
rect 7609 21188 7665 21244
rect 7665 21188 7669 21244
rect 7605 21184 7669 21188
rect 7685 21244 7749 21248
rect 7685 21188 7689 21244
rect 7689 21188 7745 21244
rect 7745 21188 7749 21244
rect 7685 21184 7749 21188
rect 3549 20700 3613 20704
rect 3549 20644 3553 20700
rect 3553 20644 3609 20700
rect 3609 20644 3613 20700
rect 3549 20640 3613 20644
rect 3629 20700 3693 20704
rect 3629 20644 3633 20700
rect 3633 20644 3689 20700
rect 3689 20644 3693 20700
rect 3629 20640 3693 20644
rect 3709 20700 3773 20704
rect 3709 20644 3713 20700
rect 3713 20644 3769 20700
rect 3769 20644 3773 20700
rect 3709 20640 3773 20644
rect 3789 20700 3853 20704
rect 3789 20644 3793 20700
rect 3793 20644 3849 20700
rect 3849 20644 3853 20700
rect 3789 20640 3853 20644
rect 6146 20700 6210 20704
rect 6146 20644 6150 20700
rect 6150 20644 6206 20700
rect 6206 20644 6210 20700
rect 6146 20640 6210 20644
rect 6226 20700 6290 20704
rect 6226 20644 6230 20700
rect 6230 20644 6286 20700
rect 6286 20644 6290 20700
rect 6226 20640 6290 20644
rect 6306 20700 6370 20704
rect 6306 20644 6310 20700
rect 6310 20644 6366 20700
rect 6366 20644 6370 20700
rect 6306 20640 6370 20644
rect 6386 20700 6450 20704
rect 6386 20644 6390 20700
rect 6390 20644 6446 20700
rect 6446 20644 6450 20700
rect 6386 20640 6450 20644
rect 2250 20156 2314 20160
rect 2250 20100 2254 20156
rect 2254 20100 2310 20156
rect 2310 20100 2314 20156
rect 2250 20096 2314 20100
rect 2330 20156 2394 20160
rect 2330 20100 2334 20156
rect 2334 20100 2390 20156
rect 2390 20100 2394 20156
rect 2330 20096 2394 20100
rect 2410 20156 2474 20160
rect 2410 20100 2414 20156
rect 2414 20100 2470 20156
rect 2470 20100 2474 20156
rect 2410 20096 2474 20100
rect 2490 20156 2554 20160
rect 2490 20100 2494 20156
rect 2494 20100 2550 20156
rect 2550 20100 2554 20156
rect 2490 20096 2554 20100
rect 4848 20156 4912 20160
rect 4848 20100 4852 20156
rect 4852 20100 4908 20156
rect 4908 20100 4912 20156
rect 4848 20096 4912 20100
rect 4928 20156 4992 20160
rect 4928 20100 4932 20156
rect 4932 20100 4988 20156
rect 4988 20100 4992 20156
rect 4928 20096 4992 20100
rect 5008 20156 5072 20160
rect 5008 20100 5012 20156
rect 5012 20100 5068 20156
rect 5068 20100 5072 20156
rect 5008 20096 5072 20100
rect 5088 20156 5152 20160
rect 5088 20100 5092 20156
rect 5092 20100 5148 20156
rect 5148 20100 5152 20156
rect 5088 20096 5152 20100
rect 7445 20156 7509 20160
rect 7445 20100 7449 20156
rect 7449 20100 7505 20156
rect 7505 20100 7509 20156
rect 7445 20096 7509 20100
rect 7525 20156 7589 20160
rect 7525 20100 7529 20156
rect 7529 20100 7585 20156
rect 7585 20100 7589 20156
rect 7525 20096 7589 20100
rect 7605 20156 7669 20160
rect 7605 20100 7609 20156
rect 7609 20100 7665 20156
rect 7665 20100 7669 20156
rect 7605 20096 7669 20100
rect 7685 20156 7749 20160
rect 7685 20100 7689 20156
rect 7689 20100 7745 20156
rect 7745 20100 7749 20156
rect 7685 20096 7749 20100
rect 3549 19612 3613 19616
rect 3549 19556 3553 19612
rect 3553 19556 3609 19612
rect 3609 19556 3613 19612
rect 3549 19552 3613 19556
rect 3629 19612 3693 19616
rect 3629 19556 3633 19612
rect 3633 19556 3689 19612
rect 3689 19556 3693 19612
rect 3629 19552 3693 19556
rect 3709 19612 3773 19616
rect 3709 19556 3713 19612
rect 3713 19556 3769 19612
rect 3769 19556 3773 19612
rect 3709 19552 3773 19556
rect 3789 19612 3853 19616
rect 3789 19556 3793 19612
rect 3793 19556 3849 19612
rect 3849 19556 3853 19612
rect 3789 19552 3853 19556
rect 6146 19612 6210 19616
rect 6146 19556 6150 19612
rect 6150 19556 6206 19612
rect 6206 19556 6210 19612
rect 6146 19552 6210 19556
rect 6226 19612 6290 19616
rect 6226 19556 6230 19612
rect 6230 19556 6286 19612
rect 6286 19556 6290 19612
rect 6226 19552 6290 19556
rect 6306 19612 6370 19616
rect 6306 19556 6310 19612
rect 6310 19556 6366 19612
rect 6366 19556 6370 19612
rect 6306 19552 6370 19556
rect 6386 19612 6450 19616
rect 6386 19556 6390 19612
rect 6390 19556 6446 19612
rect 6446 19556 6450 19612
rect 6386 19552 6450 19556
rect 2250 19068 2314 19072
rect 2250 19012 2254 19068
rect 2254 19012 2310 19068
rect 2310 19012 2314 19068
rect 2250 19008 2314 19012
rect 2330 19068 2394 19072
rect 2330 19012 2334 19068
rect 2334 19012 2390 19068
rect 2390 19012 2394 19068
rect 2330 19008 2394 19012
rect 2410 19068 2474 19072
rect 2410 19012 2414 19068
rect 2414 19012 2470 19068
rect 2470 19012 2474 19068
rect 2410 19008 2474 19012
rect 2490 19068 2554 19072
rect 2490 19012 2494 19068
rect 2494 19012 2550 19068
rect 2550 19012 2554 19068
rect 2490 19008 2554 19012
rect 4848 19068 4912 19072
rect 4848 19012 4852 19068
rect 4852 19012 4908 19068
rect 4908 19012 4912 19068
rect 4848 19008 4912 19012
rect 4928 19068 4992 19072
rect 4928 19012 4932 19068
rect 4932 19012 4988 19068
rect 4988 19012 4992 19068
rect 4928 19008 4992 19012
rect 5008 19068 5072 19072
rect 5008 19012 5012 19068
rect 5012 19012 5068 19068
rect 5068 19012 5072 19068
rect 5008 19008 5072 19012
rect 5088 19068 5152 19072
rect 5088 19012 5092 19068
rect 5092 19012 5148 19068
rect 5148 19012 5152 19068
rect 5088 19008 5152 19012
rect 7445 19068 7509 19072
rect 7445 19012 7449 19068
rect 7449 19012 7505 19068
rect 7505 19012 7509 19068
rect 7445 19008 7509 19012
rect 7525 19068 7589 19072
rect 7525 19012 7529 19068
rect 7529 19012 7585 19068
rect 7585 19012 7589 19068
rect 7525 19008 7589 19012
rect 7605 19068 7669 19072
rect 7605 19012 7609 19068
rect 7609 19012 7665 19068
rect 7665 19012 7669 19068
rect 7605 19008 7669 19012
rect 7685 19068 7749 19072
rect 7685 19012 7689 19068
rect 7689 19012 7745 19068
rect 7745 19012 7749 19068
rect 7685 19008 7749 19012
rect 3549 18524 3613 18528
rect 3549 18468 3553 18524
rect 3553 18468 3609 18524
rect 3609 18468 3613 18524
rect 3549 18464 3613 18468
rect 3629 18524 3693 18528
rect 3629 18468 3633 18524
rect 3633 18468 3689 18524
rect 3689 18468 3693 18524
rect 3629 18464 3693 18468
rect 3709 18524 3773 18528
rect 3709 18468 3713 18524
rect 3713 18468 3769 18524
rect 3769 18468 3773 18524
rect 3709 18464 3773 18468
rect 3789 18524 3853 18528
rect 3789 18468 3793 18524
rect 3793 18468 3849 18524
rect 3849 18468 3853 18524
rect 3789 18464 3853 18468
rect 6146 18524 6210 18528
rect 6146 18468 6150 18524
rect 6150 18468 6206 18524
rect 6206 18468 6210 18524
rect 6146 18464 6210 18468
rect 6226 18524 6290 18528
rect 6226 18468 6230 18524
rect 6230 18468 6286 18524
rect 6286 18468 6290 18524
rect 6226 18464 6290 18468
rect 6306 18524 6370 18528
rect 6306 18468 6310 18524
rect 6310 18468 6366 18524
rect 6366 18468 6370 18524
rect 6306 18464 6370 18468
rect 6386 18524 6450 18528
rect 6386 18468 6390 18524
rect 6390 18468 6446 18524
rect 6446 18468 6450 18524
rect 6386 18464 6450 18468
rect 2250 17980 2314 17984
rect 2250 17924 2254 17980
rect 2254 17924 2310 17980
rect 2310 17924 2314 17980
rect 2250 17920 2314 17924
rect 2330 17980 2394 17984
rect 2330 17924 2334 17980
rect 2334 17924 2390 17980
rect 2390 17924 2394 17980
rect 2330 17920 2394 17924
rect 2410 17980 2474 17984
rect 2410 17924 2414 17980
rect 2414 17924 2470 17980
rect 2470 17924 2474 17980
rect 2410 17920 2474 17924
rect 2490 17980 2554 17984
rect 2490 17924 2494 17980
rect 2494 17924 2550 17980
rect 2550 17924 2554 17980
rect 2490 17920 2554 17924
rect 4848 17980 4912 17984
rect 4848 17924 4852 17980
rect 4852 17924 4908 17980
rect 4908 17924 4912 17980
rect 4848 17920 4912 17924
rect 4928 17980 4992 17984
rect 4928 17924 4932 17980
rect 4932 17924 4988 17980
rect 4988 17924 4992 17980
rect 4928 17920 4992 17924
rect 5008 17980 5072 17984
rect 5008 17924 5012 17980
rect 5012 17924 5068 17980
rect 5068 17924 5072 17980
rect 5008 17920 5072 17924
rect 5088 17980 5152 17984
rect 5088 17924 5092 17980
rect 5092 17924 5148 17980
rect 5148 17924 5152 17980
rect 5088 17920 5152 17924
rect 7445 17980 7509 17984
rect 7445 17924 7449 17980
rect 7449 17924 7505 17980
rect 7505 17924 7509 17980
rect 7445 17920 7509 17924
rect 7525 17980 7589 17984
rect 7525 17924 7529 17980
rect 7529 17924 7585 17980
rect 7585 17924 7589 17980
rect 7525 17920 7589 17924
rect 7605 17980 7669 17984
rect 7605 17924 7609 17980
rect 7609 17924 7665 17980
rect 7665 17924 7669 17980
rect 7605 17920 7669 17924
rect 7685 17980 7749 17984
rect 7685 17924 7689 17980
rect 7689 17924 7745 17980
rect 7745 17924 7749 17980
rect 7685 17920 7749 17924
rect 3549 17436 3613 17440
rect 3549 17380 3553 17436
rect 3553 17380 3609 17436
rect 3609 17380 3613 17436
rect 3549 17376 3613 17380
rect 3629 17436 3693 17440
rect 3629 17380 3633 17436
rect 3633 17380 3689 17436
rect 3689 17380 3693 17436
rect 3629 17376 3693 17380
rect 3709 17436 3773 17440
rect 3709 17380 3713 17436
rect 3713 17380 3769 17436
rect 3769 17380 3773 17436
rect 3709 17376 3773 17380
rect 3789 17436 3853 17440
rect 3789 17380 3793 17436
rect 3793 17380 3849 17436
rect 3849 17380 3853 17436
rect 3789 17376 3853 17380
rect 6146 17436 6210 17440
rect 6146 17380 6150 17436
rect 6150 17380 6206 17436
rect 6206 17380 6210 17436
rect 6146 17376 6210 17380
rect 6226 17436 6290 17440
rect 6226 17380 6230 17436
rect 6230 17380 6286 17436
rect 6286 17380 6290 17436
rect 6226 17376 6290 17380
rect 6306 17436 6370 17440
rect 6306 17380 6310 17436
rect 6310 17380 6366 17436
rect 6366 17380 6370 17436
rect 6306 17376 6370 17380
rect 6386 17436 6450 17440
rect 6386 17380 6390 17436
rect 6390 17380 6446 17436
rect 6446 17380 6450 17436
rect 6386 17376 6450 17380
rect 2250 16892 2314 16896
rect 2250 16836 2254 16892
rect 2254 16836 2310 16892
rect 2310 16836 2314 16892
rect 2250 16832 2314 16836
rect 2330 16892 2394 16896
rect 2330 16836 2334 16892
rect 2334 16836 2390 16892
rect 2390 16836 2394 16892
rect 2330 16832 2394 16836
rect 2410 16892 2474 16896
rect 2410 16836 2414 16892
rect 2414 16836 2470 16892
rect 2470 16836 2474 16892
rect 2410 16832 2474 16836
rect 2490 16892 2554 16896
rect 2490 16836 2494 16892
rect 2494 16836 2550 16892
rect 2550 16836 2554 16892
rect 2490 16832 2554 16836
rect 4848 16892 4912 16896
rect 4848 16836 4852 16892
rect 4852 16836 4908 16892
rect 4908 16836 4912 16892
rect 4848 16832 4912 16836
rect 4928 16892 4992 16896
rect 4928 16836 4932 16892
rect 4932 16836 4988 16892
rect 4988 16836 4992 16892
rect 4928 16832 4992 16836
rect 5008 16892 5072 16896
rect 5008 16836 5012 16892
rect 5012 16836 5068 16892
rect 5068 16836 5072 16892
rect 5008 16832 5072 16836
rect 5088 16892 5152 16896
rect 5088 16836 5092 16892
rect 5092 16836 5148 16892
rect 5148 16836 5152 16892
rect 5088 16832 5152 16836
rect 7445 16892 7509 16896
rect 7445 16836 7449 16892
rect 7449 16836 7505 16892
rect 7505 16836 7509 16892
rect 7445 16832 7509 16836
rect 7525 16892 7589 16896
rect 7525 16836 7529 16892
rect 7529 16836 7585 16892
rect 7585 16836 7589 16892
rect 7525 16832 7589 16836
rect 7605 16892 7669 16896
rect 7605 16836 7609 16892
rect 7609 16836 7665 16892
rect 7665 16836 7669 16892
rect 7605 16832 7669 16836
rect 7685 16892 7749 16896
rect 7685 16836 7689 16892
rect 7689 16836 7745 16892
rect 7745 16836 7749 16892
rect 7685 16832 7749 16836
rect 3549 16348 3613 16352
rect 3549 16292 3553 16348
rect 3553 16292 3609 16348
rect 3609 16292 3613 16348
rect 3549 16288 3613 16292
rect 3629 16348 3693 16352
rect 3629 16292 3633 16348
rect 3633 16292 3689 16348
rect 3689 16292 3693 16348
rect 3629 16288 3693 16292
rect 3709 16348 3773 16352
rect 3709 16292 3713 16348
rect 3713 16292 3769 16348
rect 3769 16292 3773 16348
rect 3709 16288 3773 16292
rect 3789 16348 3853 16352
rect 3789 16292 3793 16348
rect 3793 16292 3849 16348
rect 3849 16292 3853 16348
rect 3789 16288 3853 16292
rect 6146 16348 6210 16352
rect 6146 16292 6150 16348
rect 6150 16292 6206 16348
rect 6206 16292 6210 16348
rect 6146 16288 6210 16292
rect 6226 16348 6290 16352
rect 6226 16292 6230 16348
rect 6230 16292 6286 16348
rect 6286 16292 6290 16348
rect 6226 16288 6290 16292
rect 6306 16348 6370 16352
rect 6306 16292 6310 16348
rect 6310 16292 6366 16348
rect 6366 16292 6370 16348
rect 6306 16288 6370 16292
rect 6386 16348 6450 16352
rect 6386 16292 6390 16348
rect 6390 16292 6446 16348
rect 6446 16292 6450 16348
rect 6386 16288 6450 16292
rect 2250 15804 2314 15808
rect 2250 15748 2254 15804
rect 2254 15748 2310 15804
rect 2310 15748 2314 15804
rect 2250 15744 2314 15748
rect 2330 15804 2394 15808
rect 2330 15748 2334 15804
rect 2334 15748 2390 15804
rect 2390 15748 2394 15804
rect 2330 15744 2394 15748
rect 2410 15804 2474 15808
rect 2410 15748 2414 15804
rect 2414 15748 2470 15804
rect 2470 15748 2474 15804
rect 2410 15744 2474 15748
rect 2490 15804 2554 15808
rect 2490 15748 2494 15804
rect 2494 15748 2550 15804
rect 2550 15748 2554 15804
rect 2490 15744 2554 15748
rect 4848 15804 4912 15808
rect 4848 15748 4852 15804
rect 4852 15748 4908 15804
rect 4908 15748 4912 15804
rect 4848 15744 4912 15748
rect 4928 15804 4992 15808
rect 4928 15748 4932 15804
rect 4932 15748 4988 15804
rect 4988 15748 4992 15804
rect 4928 15744 4992 15748
rect 5008 15804 5072 15808
rect 5008 15748 5012 15804
rect 5012 15748 5068 15804
rect 5068 15748 5072 15804
rect 5008 15744 5072 15748
rect 5088 15804 5152 15808
rect 5088 15748 5092 15804
rect 5092 15748 5148 15804
rect 5148 15748 5152 15804
rect 5088 15744 5152 15748
rect 7445 15804 7509 15808
rect 7445 15748 7449 15804
rect 7449 15748 7505 15804
rect 7505 15748 7509 15804
rect 7445 15744 7509 15748
rect 7525 15804 7589 15808
rect 7525 15748 7529 15804
rect 7529 15748 7585 15804
rect 7585 15748 7589 15804
rect 7525 15744 7589 15748
rect 7605 15804 7669 15808
rect 7605 15748 7609 15804
rect 7609 15748 7665 15804
rect 7665 15748 7669 15804
rect 7605 15744 7669 15748
rect 7685 15804 7749 15808
rect 7685 15748 7689 15804
rect 7689 15748 7745 15804
rect 7745 15748 7749 15804
rect 7685 15744 7749 15748
rect 3549 15260 3613 15264
rect 3549 15204 3553 15260
rect 3553 15204 3609 15260
rect 3609 15204 3613 15260
rect 3549 15200 3613 15204
rect 3629 15260 3693 15264
rect 3629 15204 3633 15260
rect 3633 15204 3689 15260
rect 3689 15204 3693 15260
rect 3629 15200 3693 15204
rect 3709 15260 3773 15264
rect 3709 15204 3713 15260
rect 3713 15204 3769 15260
rect 3769 15204 3773 15260
rect 3709 15200 3773 15204
rect 3789 15260 3853 15264
rect 3789 15204 3793 15260
rect 3793 15204 3849 15260
rect 3849 15204 3853 15260
rect 3789 15200 3853 15204
rect 6146 15260 6210 15264
rect 6146 15204 6150 15260
rect 6150 15204 6206 15260
rect 6206 15204 6210 15260
rect 6146 15200 6210 15204
rect 6226 15260 6290 15264
rect 6226 15204 6230 15260
rect 6230 15204 6286 15260
rect 6286 15204 6290 15260
rect 6226 15200 6290 15204
rect 6306 15260 6370 15264
rect 6306 15204 6310 15260
rect 6310 15204 6366 15260
rect 6366 15204 6370 15260
rect 6306 15200 6370 15204
rect 6386 15260 6450 15264
rect 6386 15204 6390 15260
rect 6390 15204 6446 15260
rect 6446 15204 6450 15260
rect 6386 15200 6450 15204
rect 2250 14716 2314 14720
rect 2250 14660 2254 14716
rect 2254 14660 2310 14716
rect 2310 14660 2314 14716
rect 2250 14656 2314 14660
rect 2330 14716 2394 14720
rect 2330 14660 2334 14716
rect 2334 14660 2390 14716
rect 2390 14660 2394 14716
rect 2330 14656 2394 14660
rect 2410 14716 2474 14720
rect 2410 14660 2414 14716
rect 2414 14660 2470 14716
rect 2470 14660 2474 14716
rect 2410 14656 2474 14660
rect 2490 14716 2554 14720
rect 2490 14660 2494 14716
rect 2494 14660 2550 14716
rect 2550 14660 2554 14716
rect 2490 14656 2554 14660
rect 4848 14716 4912 14720
rect 4848 14660 4852 14716
rect 4852 14660 4908 14716
rect 4908 14660 4912 14716
rect 4848 14656 4912 14660
rect 4928 14716 4992 14720
rect 4928 14660 4932 14716
rect 4932 14660 4988 14716
rect 4988 14660 4992 14716
rect 4928 14656 4992 14660
rect 5008 14716 5072 14720
rect 5008 14660 5012 14716
rect 5012 14660 5068 14716
rect 5068 14660 5072 14716
rect 5008 14656 5072 14660
rect 5088 14716 5152 14720
rect 5088 14660 5092 14716
rect 5092 14660 5148 14716
rect 5148 14660 5152 14716
rect 5088 14656 5152 14660
rect 7445 14716 7509 14720
rect 7445 14660 7449 14716
rect 7449 14660 7505 14716
rect 7505 14660 7509 14716
rect 7445 14656 7509 14660
rect 7525 14716 7589 14720
rect 7525 14660 7529 14716
rect 7529 14660 7585 14716
rect 7585 14660 7589 14716
rect 7525 14656 7589 14660
rect 7605 14716 7669 14720
rect 7605 14660 7609 14716
rect 7609 14660 7665 14716
rect 7665 14660 7669 14716
rect 7605 14656 7669 14660
rect 7685 14716 7749 14720
rect 7685 14660 7689 14716
rect 7689 14660 7745 14716
rect 7745 14660 7749 14716
rect 7685 14656 7749 14660
rect 3549 14172 3613 14176
rect 3549 14116 3553 14172
rect 3553 14116 3609 14172
rect 3609 14116 3613 14172
rect 3549 14112 3613 14116
rect 3629 14172 3693 14176
rect 3629 14116 3633 14172
rect 3633 14116 3689 14172
rect 3689 14116 3693 14172
rect 3629 14112 3693 14116
rect 3709 14172 3773 14176
rect 3709 14116 3713 14172
rect 3713 14116 3769 14172
rect 3769 14116 3773 14172
rect 3709 14112 3773 14116
rect 3789 14172 3853 14176
rect 3789 14116 3793 14172
rect 3793 14116 3849 14172
rect 3849 14116 3853 14172
rect 3789 14112 3853 14116
rect 6146 14172 6210 14176
rect 6146 14116 6150 14172
rect 6150 14116 6206 14172
rect 6206 14116 6210 14172
rect 6146 14112 6210 14116
rect 6226 14172 6290 14176
rect 6226 14116 6230 14172
rect 6230 14116 6286 14172
rect 6286 14116 6290 14172
rect 6226 14112 6290 14116
rect 6306 14172 6370 14176
rect 6306 14116 6310 14172
rect 6310 14116 6366 14172
rect 6366 14116 6370 14172
rect 6306 14112 6370 14116
rect 6386 14172 6450 14176
rect 6386 14116 6390 14172
rect 6390 14116 6446 14172
rect 6446 14116 6450 14172
rect 6386 14112 6450 14116
rect 2250 13628 2314 13632
rect 2250 13572 2254 13628
rect 2254 13572 2310 13628
rect 2310 13572 2314 13628
rect 2250 13568 2314 13572
rect 2330 13628 2394 13632
rect 2330 13572 2334 13628
rect 2334 13572 2390 13628
rect 2390 13572 2394 13628
rect 2330 13568 2394 13572
rect 2410 13628 2474 13632
rect 2410 13572 2414 13628
rect 2414 13572 2470 13628
rect 2470 13572 2474 13628
rect 2410 13568 2474 13572
rect 2490 13628 2554 13632
rect 2490 13572 2494 13628
rect 2494 13572 2550 13628
rect 2550 13572 2554 13628
rect 2490 13568 2554 13572
rect 4848 13628 4912 13632
rect 4848 13572 4852 13628
rect 4852 13572 4908 13628
rect 4908 13572 4912 13628
rect 4848 13568 4912 13572
rect 4928 13628 4992 13632
rect 4928 13572 4932 13628
rect 4932 13572 4988 13628
rect 4988 13572 4992 13628
rect 4928 13568 4992 13572
rect 5008 13628 5072 13632
rect 5008 13572 5012 13628
rect 5012 13572 5068 13628
rect 5068 13572 5072 13628
rect 5008 13568 5072 13572
rect 5088 13628 5152 13632
rect 5088 13572 5092 13628
rect 5092 13572 5148 13628
rect 5148 13572 5152 13628
rect 5088 13568 5152 13572
rect 7445 13628 7509 13632
rect 7445 13572 7449 13628
rect 7449 13572 7505 13628
rect 7505 13572 7509 13628
rect 7445 13568 7509 13572
rect 7525 13628 7589 13632
rect 7525 13572 7529 13628
rect 7529 13572 7585 13628
rect 7585 13572 7589 13628
rect 7525 13568 7589 13572
rect 7605 13628 7669 13632
rect 7605 13572 7609 13628
rect 7609 13572 7665 13628
rect 7665 13572 7669 13628
rect 7605 13568 7669 13572
rect 7685 13628 7749 13632
rect 7685 13572 7689 13628
rect 7689 13572 7745 13628
rect 7745 13572 7749 13628
rect 7685 13568 7749 13572
rect 3549 13084 3613 13088
rect 3549 13028 3553 13084
rect 3553 13028 3609 13084
rect 3609 13028 3613 13084
rect 3549 13024 3613 13028
rect 3629 13084 3693 13088
rect 3629 13028 3633 13084
rect 3633 13028 3689 13084
rect 3689 13028 3693 13084
rect 3629 13024 3693 13028
rect 3709 13084 3773 13088
rect 3709 13028 3713 13084
rect 3713 13028 3769 13084
rect 3769 13028 3773 13084
rect 3709 13024 3773 13028
rect 3789 13084 3853 13088
rect 3789 13028 3793 13084
rect 3793 13028 3849 13084
rect 3849 13028 3853 13084
rect 3789 13024 3853 13028
rect 6146 13084 6210 13088
rect 6146 13028 6150 13084
rect 6150 13028 6206 13084
rect 6206 13028 6210 13084
rect 6146 13024 6210 13028
rect 6226 13084 6290 13088
rect 6226 13028 6230 13084
rect 6230 13028 6286 13084
rect 6286 13028 6290 13084
rect 6226 13024 6290 13028
rect 6306 13084 6370 13088
rect 6306 13028 6310 13084
rect 6310 13028 6366 13084
rect 6366 13028 6370 13084
rect 6306 13024 6370 13028
rect 6386 13084 6450 13088
rect 6386 13028 6390 13084
rect 6390 13028 6446 13084
rect 6446 13028 6450 13084
rect 6386 13024 6450 13028
rect 2250 12540 2314 12544
rect 2250 12484 2254 12540
rect 2254 12484 2310 12540
rect 2310 12484 2314 12540
rect 2250 12480 2314 12484
rect 2330 12540 2394 12544
rect 2330 12484 2334 12540
rect 2334 12484 2390 12540
rect 2390 12484 2394 12540
rect 2330 12480 2394 12484
rect 2410 12540 2474 12544
rect 2410 12484 2414 12540
rect 2414 12484 2470 12540
rect 2470 12484 2474 12540
rect 2410 12480 2474 12484
rect 2490 12540 2554 12544
rect 2490 12484 2494 12540
rect 2494 12484 2550 12540
rect 2550 12484 2554 12540
rect 2490 12480 2554 12484
rect 4848 12540 4912 12544
rect 4848 12484 4852 12540
rect 4852 12484 4908 12540
rect 4908 12484 4912 12540
rect 4848 12480 4912 12484
rect 4928 12540 4992 12544
rect 4928 12484 4932 12540
rect 4932 12484 4988 12540
rect 4988 12484 4992 12540
rect 4928 12480 4992 12484
rect 5008 12540 5072 12544
rect 5008 12484 5012 12540
rect 5012 12484 5068 12540
rect 5068 12484 5072 12540
rect 5008 12480 5072 12484
rect 5088 12540 5152 12544
rect 5088 12484 5092 12540
rect 5092 12484 5148 12540
rect 5148 12484 5152 12540
rect 5088 12480 5152 12484
rect 7445 12540 7509 12544
rect 7445 12484 7449 12540
rect 7449 12484 7505 12540
rect 7505 12484 7509 12540
rect 7445 12480 7509 12484
rect 7525 12540 7589 12544
rect 7525 12484 7529 12540
rect 7529 12484 7585 12540
rect 7585 12484 7589 12540
rect 7525 12480 7589 12484
rect 7605 12540 7669 12544
rect 7605 12484 7609 12540
rect 7609 12484 7665 12540
rect 7665 12484 7669 12540
rect 7605 12480 7669 12484
rect 7685 12540 7749 12544
rect 7685 12484 7689 12540
rect 7689 12484 7745 12540
rect 7745 12484 7749 12540
rect 7685 12480 7749 12484
rect 3549 11996 3613 12000
rect 3549 11940 3553 11996
rect 3553 11940 3609 11996
rect 3609 11940 3613 11996
rect 3549 11936 3613 11940
rect 3629 11996 3693 12000
rect 3629 11940 3633 11996
rect 3633 11940 3689 11996
rect 3689 11940 3693 11996
rect 3629 11936 3693 11940
rect 3709 11996 3773 12000
rect 3709 11940 3713 11996
rect 3713 11940 3769 11996
rect 3769 11940 3773 11996
rect 3709 11936 3773 11940
rect 3789 11996 3853 12000
rect 3789 11940 3793 11996
rect 3793 11940 3849 11996
rect 3849 11940 3853 11996
rect 3789 11936 3853 11940
rect 6146 11996 6210 12000
rect 6146 11940 6150 11996
rect 6150 11940 6206 11996
rect 6206 11940 6210 11996
rect 6146 11936 6210 11940
rect 6226 11996 6290 12000
rect 6226 11940 6230 11996
rect 6230 11940 6286 11996
rect 6286 11940 6290 11996
rect 6226 11936 6290 11940
rect 6306 11996 6370 12000
rect 6306 11940 6310 11996
rect 6310 11940 6366 11996
rect 6366 11940 6370 11996
rect 6306 11936 6370 11940
rect 6386 11996 6450 12000
rect 6386 11940 6390 11996
rect 6390 11940 6446 11996
rect 6446 11940 6450 11996
rect 6386 11936 6450 11940
rect 2250 11452 2314 11456
rect 2250 11396 2254 11452
rect 2254 11396 2310 11452
rect 2310 11396 2314 11452
rect 2250 11392 2314 11396
rect 2330 11452 2394 11456
rect 2330 11396 2334 11452
rect 2334 11396 2390 11452
rect 2390 11396 2394 11452
rect 2330 11392 2394 11396
rect 2410 11452 2474 11456
rect 2410 11396 2414 11452
rect 2414 11396 2470 11452
rect 2470 11396 2474 11452
rect 2410 11392 2474 11396
rect 2490 11452 2554 11456
rect 2490 11396 2494 11452
rect 2494 11396 2550 11452
rect 2550 11396 2554 11452
rect 2490 11392 2554 11396
rect 4848 11452 4912 11456
rect 4848 11396 4852 11452
rect 4852 11396 4908 11452
rect 4908 11396 4912 11452
rect 4848 11392 4912 11396
rect 4928 11452 4992 11456
rect 4928 11396 4932 11452
rect 4932 11396 4988 11452
rect 4988 11396 4992 11452
rect 4928 11392 4992 11396
rect 5008 11452 5072 11456
rect 5008 11396 5012 11452
rect 5012 11396 5068 11452
rect 5068 11396 5072 11452
rect 5008 11392 5072 11396
rect 5088 11452 5152 11456
rect 5088 11396 5092 11452
rect 5092 11396 5148 11452
rect 5148 11396 5152 11452
rect 5088 11392 5152 11396
rect 7445 11452 7509 11456
rect 7445 11396 7449 11452
rect 7449 11396 7505 11452
rect 7505 11396 7509 11452
rect 7445 11392 7509 11396
rect 7525 11452 7589 11456
rect 7525 11396 7529 11452
rect 7529 11396 7585 11452
rect 7585 11396 7589 11452
rect 7525 11392 7589 11396
rect 7605 11452 7669 11456
rect 7605 11396 7609 11452
rect 7609 11396 7665 11452
rect 7665 11396 7669 11452
rect 7605 11392 7669 11396
rect 7685 11452 7749 11456
rect 7685 11396 7689 11452
rect 7689 11396 7745 11452
rect 7745 11396 7749 11452
rect 7685 11392 7749 11396
rect 3549 10908 3613 10912
rect 3549 10852 3553 10908
rect 3553 10852 3609 10908
rect 3609 10852 3613 10908
rect 3549 10848 3613 10852
rect 3629 10908 3693 10912
rect 3629 10852 3633 10908
rect 3633 10852 3689 10908
rect 3689 10852 3693 10908
rect 3629 10848 3693 10852
rect 3709 10908 3773 10912
rect 3709 10852 3713 10908
rect 3713 10852 3769 10908
rect 3769 10852 3773 10908
rect 3709 10848 3773 10852
rect 3789 10908 3853 10912
rect 3789 10852 3793 10908
rect 3793 10852 3849 10908
rect 3849 10852 3853 10908
rect 3789 10848 3853 10852
rect 6146 10908 6210 10912
rect 6146 10852 6150 10908
rect 6150 10852 6206 10908
rect 6206 10852 6210 10908
rect 6146 10848 6210 10852
rect 6226 10908 6290 10912
rect 6226 10852 6230 10908
rect 6230 10852 6286 10908
rect 6286 10852 6290 10908
rect 6226 10848 6290 10852
rect 6306 10908 6370 10912
rect 6306 10852 6310 10908
rect 6310 10852 6366 10908
rect 6366 10852 6370 10908
rect 6306 10848 6370 10852
rect 6386 10908 6450 10912
rect 6386 10852 6390 10908
rect 6390 10852 6446 10908
rect 6446 10852 6450 10908
rect 6386 10848 6450 10852
rect 2250 10364 2314 10368
rect 2250 10308 2254 10364
rect 2254 10308 2310 10364
rect 2310 10308 2314 10364
rect 2250 10304 2314 10308
rect 2330 10364 2394 10368
rect 2330 10308 2334 10364
rect 2334 10308 2390 10364
rect 2390 10308 2394 10364
rect 2330 10304 2394 10308
rect 2410 10364 2474 10368
rect 2410 10308 2414 10364
rect 2414 10308 2470 10364
rect 2470 10308 2474 10364
rect 2410 10304 2474 10308
rect 2490 10364 2554 10368
rect 2490 10308 2494 10364
rect 2494 10308 2550 10364
rect 2550 10308 2554 10364
rect 2490 10304 2554 10308
rect 4848 10364 4912 10368
rect 4848 10308 4852 10364
rect 4852 10308 4908 10364
rect 4908 10308 4912 10364
rect 4848 10304 4912 10308
rect 4928 10364 4992 10368
rect 4928 10308 4932 10364
rect 4932 10308 4988 10364
rect 4988 10308 4992 10364
rect 4928 10304 4992 10308
rect 5008 10364 5072 10368
rect 5008 10308 5012 10364
rect 5012 10308 5068 10364
rect 5068 10308 5072 10364
rect 5008 10304 5072 10308
rect 5088 10364 5152 10368
rect 5088 10308 5092 10364
rect 5092 10308 5148 10364
rect 5148 10308 5152 10364
rect 5088 10304 5152 10308
rect 7445 10364 7509 10368
rect 7445 10308 7449 10364
rect 7449 10308 7505 10364
rect 7505 10308 7509 10364
rect 7445 10304 7509 10308
rect 7525 10364 7589 10368
rect 7525 10308 7529 10364
rect 7529 10308 7585 10364
rect 7585 10308 7589 10364
rect 7525 10304 7589 10308
rect 7605 10364 7669 10368
rect 7605 10308 7609 10364
rect 7609 10308 7665 10364
rect 7665 10308 7669 10364
rect 7605 10304 7669 10308
rect 7685 10364 7749 10368
rect 7685 10308 7689 10364
rect 7689 10308 7745 10364
rect 7745 10308 7749 10364
rect 7685 10304 7749 10308
rect 3549 9820 3613 9824
rect 3549 9764 3553 9820
rect 3553 9764 3609 9820
rect 3609 9764 3613 9820
rect 3549 9760 3613 9764
rect 3629 9820 3693 9824
rect 3629 9764 3633 9820
rect 3633 9764 3689 9820
rect 3689 9764 3693 9820
rect 3629 9760 3693 9764
rect 3709 9820 3773 9824
rect 3709 9764 3713 9820
rect 3713 9764 3769 9820
rect 3769 9764 3773 9820
rect 3709 9760 3773 9764
rect 3789 9820 3853 9824
rect 3789 9764 3793 9820
rect 3793 9764 3849 9820
rect 3849 9764 3853 9820
rect 3789 9760 3853 9764
rect 6146 9820 6210 9824
rect 6146 9764 6150 9820
rect 6150 9764 6206 9820
rect 6206 9764 6210 9820
rect 6146 9760 6210 9764
rect 6226 9820 6290 9824
rect 6226 9764 6230 9820
rect 6230 9764 6286 9820
rect 6286 9764 6290 9820
rect 6226 9760 6290 9764
rect 6306 9820 6370 9824
rect 6306 9764 6310 9820
rect 6310 9764 6366 9820
rect 6366 9764 6370 9820
rect 6306 9760 6370 9764
rect 6386 9820 6450 9824
rect 6386 9764 6390 9820
rect 6390 9764 6446 9820
rect 6446 9764 6450 9820
rect 6386 9760 6450 9764
rect 2250 9276 2314 9280
rect 2250 9220 2254 9276
rect 2254 9220 2310 9276
rect 2310 9220 2314 9276
rect 2250 9216 2314 9220
rect 2330 9276 2394 9280
rect 2330 9220 2334 9276
rect 2334 9220 2390 9276
rect 2390 9220 2394 9276
rect 2330 9216 2394 9220
rect 2410 9276 2474 9280
rect 2410 9220 2414 9276
rect 2414 9220 2470 9276
rect 2470 9220 2474 9276
rect 2410 9216 2474 9220
rect 2490 9276 2554 9280
rect 2490 9220 2494 9276
rect 2494 9220 2550 9276
rect 2550 9220 2554 9276
rect 2490 9216 2554 9220
rect 4848 9276 4912 9280
rect 4848 9220 4852 9276
rect 4852 9220 4908 9276
rect 4908 9220 4912 9276
rect 4848 9216 4912 9220
rect 4928 9276 4992 9280
rect 4928 9220 4932 9276
rect 4932 9220 4988 9276
rect 4988 9220 4992 9276
rect 4928 9216 4992 9220
rect 5008 9276 5072 9280
rect 5008 9220 5012 9276
rect 5012 9220 5068 9276
rect 5068 9220 5072 9276
rect 5008 9216 5072 9220
rect 5088 9276 5152 9280
rect 5088 9220 5092 9276
rect 5092 9220 5148 9276
rect 5148 9220 5152 9276
rect 5088 9216 5152 9220
rect 7445 9276 7509 9280
rect 7445 9220 7449 9276
rect 7449 9220 7505 9276
rect 7505 9220 7509 9276
rect 7445 9216 7509 9220
rect 7525 9276 7589 9280
rect 7525 9220 7529 9276
rect 7529 9220 7585 9276
rect 7585 9220 7589 9276
rect 7525 9216 7589 9220
rect 7605 9276 7669 9280
rect 7605 9220 7609 9276
rect 7609 9220 7665 9276
rect 7665 9220 7669 9276
rect 7605 9216 7669 9220
rect 7685 9276 7749 9280
rect 7685 9220 7689 9276
rect 7689 9220 7745 9276
rect 7745 9220 7749 9276
rect 7685 9216 7749 9220
rect 3549 8732 3613 8736
rect 3549 8676 3553 8732
rect 3553 8676 3609 8732
rect 3609 8676 3613 8732
rect 3549 8672 3613 8676
rect 3629 8732 3693 8736
rect 3629 8676 3633 8732
rect 3633 8676 3689 8732
rect 3689 8676 3693 8732
rect 3629 8672 3693 8676
rect 3709 8732 3773 8736
rect 3709 8676 3713 8732
rect 3713 8676 3769 8732
rect 3769 8676 3773 8732
rect 3709 8672 3773 8676
rect 3789 8732 3853 8736
rect 3789 8676 3793 8732
rect 3793 8676 3849 8732
rect 3849 8676 3853 8732
rect 3789 8672 3853 8676
rect 6146 8732 6210 8736
rect 6146 8676 6150 8732
rect 6150 8676 6206 8732
rect 6206 8676 6210 8732
rect 6146 8672 6210 8676
rect 6226 8732 6290 8736
rect 6226 8676 6230 8732
rect 6230 8676 6286 8732
rect 6286 8676 6290 8732
rect 6226 8672 6290 8676
rect 6306 8732 6370 8736
rect 6306 8676 6310 8732
rect 6310 8676 6366 8732
rect 6366 8676 6370 8732
rect 6306 8672 6370 8676
rect 6386 8732 6450 8736
rect 6386 8676 6390 8732
rect 6390 8676 6446 8732
rect 6446 8676 6450 8732
rect 6386 8672 6450 8676
rect 2250 8188 2314 8192
rect 2250 8132 2254 8188
rect 2254 8132 2310 8188
rect 2310 8132 2314 8188
rect 2250 8128 2314 8132
rect 2330 8188 2394 8192
rect 2330 8132 2334 8188
rect 2334 8132 2390 8188
rect 2390 8132 2394 8188
rect 2330 8128 2394 8132
rect 2410 8188 2474 8192
rect 2410 8132 2414 8188
rect 2414 8132 2470 8188
rect 2470 8132 2474 8188
rect 2410 8128 2474 8132
rect 2490 8188 2554 8192
rect 2490 8132 2494 8188
rect 2494 8132 2550 8188
rect 2550 8132 2554 8188
rect 2490 8128 2554 8132
rect 4848 8188 4912 8192
rect 4848 8132 4852 8188
rect 4852 8132 4908 8188
rect 4908 8132 4912 8188
rect 4848 8128 4912 8132
rect 4928 8188 4992 8192
rect 4928 8132 4932 8188
rect 4932 8132 4988 8188
rect 4988 8132 4992 8188
rect 4928 8128 4992 8132
rect 5008 8188 5072 8192
rect 5008 8132 5012 8188
rect 5012 8132 5068 8188
rect 5068 8132 5072 8188
rect 5008 8128 5072 8132
rect 5088 8188 5152 8192
rect 5088 8132 5092 8188
rect 5092 8132 5148 8188
rect 5148 8132 5152 8188
rect 5088 8128 5152 8132
rect 7445 8188 7509 8192
rect 7445 8132 7449 8188
rect 7449 8132 7505 8188
rect 7505 8132 7509 8188
rect 7445 8128 7509 8132
rect 7525 8188 7589 8192
rect 7525 8132 7529 8188
rect 7529 8132 7585 8188
rect 7585 8132 7589 8188
rect 7525 8128 7589 8132
rect 7605 8188 7669 8192
rect 7605 8132 7609 8188
rect 7609 8132 7665 8188
rect 7665 8132 7669 8188
rect 7605 8128 7669 8132
rect 7685 8188 7749 8192
rect 7685 8132 7689 8188
rect 7689 8132 7745 8188
rect 7745 8132 7749 8188
rect 7685 8128 7749 8132
rect 3549 7644 3613 7648
rect 3549 7588 3553 7644
rect 3553 7588 3609 7644
rect 3609 7588 3613 7644
rect 3549 7584 3613 7588
rect 3629 7644 3693 7648
rect 3629 7588 3633 7644
rect 3633 7588 3689 7644
rect 3689 7588 3693 7644
rect 3629 7584 3693 7588
rect 3709 7644 3773 7648
rect 3709 7588 3713 7644
rect 3713 7588 3769 7644
rect 3769 7588 3773 7644
rect 3709 7584 3773 7588
rect 3789 7644 3853 7648
rect 3789 7588 3793 7644
rect 3793 7588 3849 7644
rect 3849 7588 3853 7644
rect 3789 7584 3853 7588
rect 6146 7644 6210 7648
rect 6146 7588 6150 7644
rect 6150 7588 6206 7644
rect 6206 7588 6210 7644
rect 6146 7584 6210 7588
rect 6226 7644 6290 7648
rect 6226 7588 6230 7644
rect 6230 7588 6286 7644
rect 6286 7588 6290 7644
rect 6226 7584 6290 7588
rect 6306 7644 6370 7648
rect 6306 7588 6310 7644
rect 6310 7588 6366 7644
rect 6366 7588 6370 7644
rect 6306 7584 6370 7588
rect 6386 7644 6450 7648
rect 6386 7588 6390 7644
rect 6390 7588 6446 7644
rect 6446 7588 6450 7644
rect 6386 7584 6450 7588
rect 2250 7100 2314 7104
rect 2250 7044 2254 7100
rect 2254 7044 2310 7100
rect 2310 7044 2314 7100
rect 2250 7040 2314 7044
rect 2330 7100 2394 7104
rect 2330 7044 2334 7100
rect 2334 7044 2390 7100
rect 2390 7044 2394 7100
rect 2330 7040 2394 7044
rect 2410 7100 2474 7104
rect 2410 7044 2414 7100
rect 2414 7044 2470 7100
rect 2470 7044 2474 7100
rect 2410 7040 2474 7044
rect 2490 7100 2554 7104
rect 2490 7044 2494 7100
rect 2494 7044 2550 7100
rect 2550 7044 2554 7100
rect 2490 7040 2554 7044
rect 4848 7100 4912 7104
rect 4848 7044 4852 7100
rect 4852 7044 4908 7100
rect 4908 7044 4912 7100
rect 4848 7040 4912 7044
rect 4928 7100 4992 7104
rect 4928 7044 4932 7100
rect 4932 7044 4988 7100
rect 4988 7044 4992 7100
rect 4928 7040 4992 7044
rect 5008 7100 5072 7104
rect 5008 7044 5012 7100
rect 5012 7044 5068 7100
rect 5068 7044 5072 7100
rect 5008 7040 5072 7044
rect 5088 7100 5152 7104
rect 5088 7044 5092 7100
rect 5092 7044 5148 7100
rect 5148 7044 5152 7100
rect 5088 7040 5152 7044
rect 7445 7100 7509 7104
rect 7445 7044 7449 7100
rect 7449 7044 7505 7100
rect 7505 7044 7509 7100
rect 7445 7040 7509 7044
rect 7525 7100 7589 7104
rect 7525 7044 7529 7100
rect 7529 7044 7585 7100
rect 7585 7044 7589 7100
rect 7525 7040 7589 7044
rect 7605 7100 7669 7104
rect 7605 7044 7609 7100
rect 7609 7044 7665 7100
rect 7665 7044 7669 7100
rect 7605 7040 7669 7044
rect 7685 7100 7749 7104
rect 7685 7044 7689 7100
rect 7689 7044 7745 7100
rect 7745 7044 7749 7100
rect 7685 7040 7749 7044
rect 3549 6556 3613 6560
rect 3549 6500 3553 6556
rect 3553 6500 3609 6556
rect 3609 6500 3613 6556
rect 3549 6496 3613 6500
rect 3629 6556 3693 6560
rect 3629 6500 3633 6556
rect 3633 6500 3689 6556
rect 3689 6500 3693 6556
rect 3629 6496 3693 6500
rect 3709 6556 3773 6560
rect 3709 6500 3713 6556
rect 3713 6500 3769 6556
rect 3769 6500 3773 6556
rect 3709 6496 3773 6500
rect 3789 6556 3853 6560
rect 3789 6500 3793 6556
rect 3793 6500 3849 6556
rect 3849 6500 3853 6556
rect 3789 6496 3853 6500
rect 6146 6556 6210 6560
rect 6146 6500 6150 6556
rect 6150 6500 6206 6556
rect 6206 6500 6210 6556
rect 6146 6496 6210 6500
rect 6226 6556 6290 6560
rect 6226 6500 6230 6556
rect 6230 6500 6286 6556
rect 6286 6500 6290 6556
rect 6226 6496 6290 6500
rect 6306 6556 6370 6560
rect 6306 6500 6310 6556
rect 6310 6500 6366 6556
rect 6366 6500 6370 6556
rect 6306 6496 6370 6500
rect 6386 6556 6450 6560
rect 6386 6500 6390 6556
rect 6390 6500 6446 6556
rect 6446 6500 6450 6556
rect 6386 6496 6450 6500
rect 2250 6012 2314 6016
rect 2250 5956 2254 6012
rect 2254 5956 2310 6012
rect 2310 5956 2314 6012
rect 2250 5952 2314 5956
rect 2330 6012 2394 6016
rect 2330 5956 2334 6012
rect 2334 5956 2390 6012
rect 2390 5956 2394 6012
rect 2330 5952 2394 5956
rect 2410 6012 2474 6016
rect 2410 5956 2414 6012
rect 2414 5956 2470 6012
rect 2470 5956 2474 6012
rect 2410 5952 2474 5956
rect 2490 6012 2554 6016
rect 2490 5956 2494 6012
rect 2494 5956 2550 6012
rect 2550 5956 2554 6012
rect 2490 5952 2554 5956
rect 4848 6012 4912 6016
rect 4848 5956 4852 6012
rect 4852 5956 4908 6012
rect 4908 5956 4912 6012
rect 4848 5952 4912 5956
rect 4928 6012 4992 6016
rect 4928 5956 4932 6012
rect 4932 5956 4988 6012
rect 4988 5956 4992 6012
rect 4928 5952 4992 5956
rect 5008 6012 5072 6016
rect 5008 5956 5012 6012
rect 5012 5956 5068 6012
rect 5068 5956 5072 6012
rect 5008 5952 5072 5956
rect 5088 6012 5152 6016
rect 5088 5956 5092 6012
rect 5092 5956 5148 6012
rect 5148 5956 5152 6012
rect 5088 5952 5152 5956
rect 7445 6012 7509 6016
rect 7445 5956 7449 6012
rect 7449 5956 7505 6012
rect 7505 5956 7509 6012
rect 7445 5952 7509 5956
rect 7525 6012 7589 6016
rect 7525 5956 7529 6012
rect 7529 5956 7585 6012
rect 7585 5956 7589 6012
rect 7525 5952 7589 5956
rect 7605 6012 7669 6016
rect 7605 5956 7609 6012
rect 7609 5956 7665 6012
rect 7665 5956 7669 6012
rect 7605 5952 7669 5956
rect 7685 6012 7749 6016
rect 7685 5956 7689 6012
rect 7689 5956 7745 6012
rect 7745 5956 7749 6012
rect 7685 5952 7749 5956
rect 3549 5468 3613 5472
rect 3549 5412 3553 5468
rect 3553 5412 3609 5468
rect 3609 5412 3613 5468
rect 3549 5408 3613 5412
rect 3629 5468 3693 5472
rect 3629 5412 3633 5468
rect 3633 5412 3689 5468
rect 3689 5412 3693 5468
rect 3629 5408 3693 5412
rect 3709 5468 3773 5472
rect 3709 5412 3713 5468
rect 3713 5412 3769 5468
rect 3769 5412 3773 5468
rect 3709 5408 3773 5412
rect 3789 5468 3853 5472
rect 3789 5412 3793 5468
rect 3793 5412 3849 5468
rect 3849 5412 3853 5468
rect 3789 5408 3853 5412
rect 6146 5468 6210 5472
rect 6146 5412 6150 5468
rect 6150 5412 6206 5468
rect 6206 5412 6210 5468
rect 6146 5408 6210 5412
rect 6226 5468 6290 5472
rect 6226 5412 6230 5468
rect 6230 5412 6286 5468
rect 6286 5412 6290 5468
rect 6226 5408 6290 5412
rect 6306 5468 6370 5472
rect 6306 5412 6310 5468
rect 6310 5412 6366 5468
rect 6366 5412 6370 5468
rect 6306 5408 6370 5412
rect 6386 5468 6450 5472
rect 6386 5412 6390 5468
rect 6390 5412 6446 5468
rect 6446 5412 6450 5468
rect 6386 5408 6450 5412
rect 2250 4924 2314 4928
rect 2250 4868 2254 4924
rect 2254 4868 2310 4924
rect 2310 4868 2314 4924
rect 2250 4864 2314 4868
rect 2330 4924 2394 4928
rect 2330 4868 2334 4924
rect 2334 4868 2390 4924
rect 2390 4868 2394 4924
rect 2330 4864 2394 4868
rect 2410 4924 2474 4928
rect 2410 4868 2414 4924
rect 2414 4868 2470 4924
rect 2470 4868 2474 4924
rect 2410 4864 2474 4868
rect 2490 4924 2554 4928
rect 2490 4868 2494 4924
rect 2494 4868 2550 4924
rect 2550 4868 2554 4924
rect 2490 4864 2554 4868
rect 4848 4924 4912 4928
rect 4848 4868 4852 4924
rect 4852 4868 4908 4924
rect 4908 4868 4912 4924
rect 4848 4864 4912 4868
rect 4928 4924 4992 4928
rect 4928 4868 4932 4924
rect 4932 4868 4988 4924
rect 4988 4868 4992 4924
rect 4928 4864 4992 4868
rect 5008 4924 5072 4928
rect 5008 4868 5012 4924
rect 5012 4868 5068 4924
rect 5068 4868 5072 4924
rect 5008 4864 5072 4868
rect 5088 4924 5152 4928
rect 5088 4868 5092 4924
rect 5092 4868 5148 4924
rect 5148 4868 5152 4924
rect 5088 4864 5152 4868
rect 7445 4924 7509 4928
rect 7445 4868 7449 4924
rect 7449 4868 7505 4924
rect 7505 4868 7509 4924
rect 7445 4864 7509 4868
rect 7525 4924 7589 4928
rect 7525 4868 7529 4924
rect 7529 4868 7585 4924
rect 7585 4868 7589 4924
rect 7525 4864 7589 4868
rect 7605 4924 7669 4928
rect 7605 4868 7609 4924
rect 7609 4868 7665 4924
rect 7665 4868 7669 4924
rect 7605 4864 7669 4868
rect 7685 4924 7749 4928
rect 7685 4868 7689 4924
rect 7689 4868 7745 4924
rect 7745 4868 7749 4924
rect 7685 4864 7749 4868
rect 3549 4380 3613 4384
rect 3549 4324 3553 4380
rect 3553 4324 3609 4380
rect 3609 4324 3613 4380
rect 3549 4320 3613 4324
rect 3629 4380 3693 4384
rect 3629 4324 3633 4380
rect 3633 4324 3689 4380
rect 3689 4324 3693 4380
rect 3629 4320 3693 4324
rect 3709 4380 3773 4384
rect 3709 4324 3713 4380
rect 3713 4324 3769 4380
rect 3769 4324 3773 4380
rect 3709 4320 3773 4324
rect 3789 4380 3853 4384
rect 3789 4324 3793 4380
rect 3793 4324 3849 4380
rect 3849 4324 3853 4380
rect 3789 4320 3853 4324
rect 6146 4380 6210 4384
rect 6146 4324 6150 4380
rect 6150 4324 6206 4380
rect 6206 4324 6210 4380
rect 6146 4320 6210 4324
rect 6226 4380 6290 4384
rect 6226 4324 6230 4380
rect 6230 4324 6286 4380
rect 6286 4324 6290 4380
rect 6226 4320 6290 4324
rect 6306 4380 6370 4384
rect 6306 4324 6310 4380
rect 6310 4324 6366 4380
rect 6366 4324 6370 4380
rect 6306 4320 6370 4324
rect 6386 4380 6450 4384
rect 6386 4324 6390 4380
rect 6390 4324 6446 4380
rect 6446 4324 6450 4380
rect 6386 4320 6450 4324
rect 2250 3836 2314 3840
rect 2250 3780 2254 3836
rect 2254 3780 2310 3836
rect 2310 3780 2314 3836
rect 2250 3776 2314 3780
rect 2330 3836 2394 3840
rect 2330 3780 2334 3836
rect 2334 3780 2390 3836
rect 2390 3780 2394 3836
rect 2330 3776 2394 3780
rect 2410 3836 2474 3840
rect 2410 3780 2414 3836
rect 2414 3780 2470 3836
rect 2470 3780 2474 3836
rect 2410 3776 2474 3780
rect 2490 3836 2554 3840
rect 2490 3780 2494 3836
rect 2494 3780 2550 3836
rect 2550 3780 2554 3836
rect 2490 3776 2554 3780
rect 4848 3836 4912 3840
rect 4848 3780 4852 3836
rect 4852 3780 4908 3836
rect 4908 3780 4912 3836
rect 4848 3776 4912 3780
rect 4928 3836 4992 3840
rect 4928 3780 4932 3836
rect 4932 3780 4988 3836
rect 4988 3780 4992 3836
rect 4928 3776 4992 3780
rect 5008 3836 5072 3840
rect 5008 3780 5012 3836
rect 5012 3780 5068 3836
rect 5068 3780 5072 3836
rect 5008 3776 5072 3780
rect 5088 3836 5152 3840
rect 5088 3780 5092 3836
rect 5092 3780 5148 3836
rect 5148 3780 5152 3836
rect 5088 3776 5152 3780
rect 7445 3836 7509 3840
rect 7445 3780 7449 3836
rect 7449 3780 7505 3836
rect 7505 3780 7509 3836
rect 7445 3776 7509 3780
rect 7525 3836 7589 3840
rect 7525 3780 7529 3836
rect 7529 3780 7585 3836
rect 7585 3780 7589 3836
rect 7525 3776 7589 3780
rect 7605 3836 7669 3840
rect 7605 3780 7609 3836
rect 7609 3780 7665 3836
rect 7665 3780 7669 3836
rect 7605 3776 7669 3780
rect 7685 3836 7749 3840
rect 7685 3780 7689 3836
rect 7689 3780 7745 3836
rect 7745 3780 7749 3836
rect 7685 3776 7749 3780
rect 3549 3292 3613 3296
rect 3549 3236 3553 3292
rect 3553 3236 3609 3292
rect 3609 3236 3613 3292
rect 3549 3232 3613 3236
rect 3629 3292 3693 3296
rect 3629 3236 3633 3292
rect 3633 3236 3689 3292
rect 3689 3236 3693 3292
rect 3629 3232 3693 3236
rect 3709 3292 3773 3296
rect 3709 3236 3713 3292
rect 3713 3236 3769 3292
rect 3769 3236 3773 3292
rect 3709 3232 3773 3236
rect 3789 3292 3853 3296
rect 3789 3236 3793 3292
rect 3793 3236 3849 3292
rect 3849 3236 3853 3292
rect 3789 3232 3853 3236
rect 6146 3292 6210 3296
rect 6146 3236 6150 3292
rect 6150 3236 6206 3292
rect 6206 3236 6210 3292
rect 6146 3232 6210 3236
rect 6226 3292 6290 3296
rect 6226 3236 6230 3292
rect 6230 3236 6286 3292
rect 6286 3236 6290 3292
rect 6226 3232 6290 3236
rect 6306 3292 6370 3296
rect 6306 3236 6310 3292
rect 6310 3236 6366 3292
rect 6366 3236 6370 3292
rect 6306 3232 6370 3236
rect 6386 3292 6450 3296
rect 6386 3236 6390 3292
rect 6390 3236 6446 3292
rect 6446 3236 6450 3292
rect 6386 3232 6450 3236
rect 2250 2748 2314 2752
rect 2250 2692 2254 2748
rect 2254 2692 2310 2748
rect 2310 2692 2314 2748
rect 2250 2688 2314 2692
rect 2330 2748 2394 2752
rect 2330 2692 2334 2748
rect 2334 2692 2390 2748
rect 2390 2692 2394 2748
rect 2330 2688 2394 2692
rect 2410 2748 2474 2752
rect 2410 2692 2414 2748
rect 2414 2692 2470 2748
rect 2470 2692 2474 2748
rect 2410 2688 2474 2692
rect 2490 2748 2554 2752
rect 2490 2692 2494 2748
rect 2494 2692 2550 2748
rect 2550 2692 2554 2748
rect 2490 2688 2554 2692
rect 4848 2748 4912 2752
rect 4848 2692 4852 2748
rect 4852 2692 4908 2748
rect 4908 2692 4912 2748
rect 4848 2688 4912 2692
rect 4928 2748 4992 2752
rect 4928 2692 4932 2748
rect 4932 2692 4988 2748
rect 4988 2692 4992 2748
rect 4928 2688 4992 2692
rect 5008 2748 5072 2752
rect 5008 2692 5012 2748
rect 5012 2692 5068 2748
rect 5068 2692 5072 2748
rect 5008 2688 5072 2692
rect 5088 2748 5152 2752
rect 5088 2692 5092 2748
rect 5092 2692 5148 2748
rect 5148 2692 5152 2748
rect 5088 2688 5152 2692
rect 7445 2748 7509 2752
rect 7445 2692 7449 2748
rect 7449 2692 7505 2748
rect 7505 2692 7509 2748
rect 7445 2688 7509 2692
rect 7525 2748 7589 2752
rect 7525 2692 7529 2748
rect 7529 2692 7585 2748
rect 7585 2692 7589 2748
rect 7525 2688 7589 2692
rect 7605 2748 7669 2752
rect 7605 2692 7609 2748
rect 7609 2692 7665 2748
rect 7665 2692 7669 2748
rect 7605 2688 7669 2692
rect 7685 2748 7749 2752
rect 7685 2692 7689 2748
rect 7689 2692 7745 2748
rect 7745 2692 7749 2748
rect 7685 2688 7749 2692
rect 3549 2204 3613 2208
rect 3549 2148 3553 2204
rect 3553 2148 3609 2204
rect 3609 2148 3613 2204
rect 3549 2144 3613 2148
rect 3629 2204 3693 2208
rect 3629 2148 3633 2204
rect 3633 2148 3689 2204
rect 3689 2148 3693 2204
rect 3629 2144 3693 2148
rect 3709 2204 3773 2208
rect 3709 2148 3713 2204
rect 3713 2148 3769 2204
rect 3769 2148 3773 2204
rect 3709 2144 3773 2148
rect 3789 2204 3853 2208
rect 3789 2148 3793 2204
rect 3793 2148 3849 2204
rect 3849 2148 3853 2204
rect 3789 2144 3853 2148
rect 6146 2204 6210 2208
rect 6146 2148 6150 2204
rect 6150 2148 6206 2204
rect 6206 2148 6210 2204
rect 6146 2144 6210 2148
rect 6226 2204 6290 2208
rect 6226 2148 6230 2204
rect 6230 2148 6286 2204
rect 6286 2148 6290 2204
rect 6226 2144 6290 2148
rect 6306 2204 6370 2208
rect 6306 2148 6310 2204
rect 6310 2148 6366 2204
rect 6366 2148 6370 2204
rect 6306 2144 6370 2148
rect 6386 2204 6450 2208
rect 6386 2148 6390 2204
rect 6390 2148 6446 2204
rect 6446 2148 6450 2204
rect 6386 2144 6450 2148
<< metal4 >>
rect 2242 22336 2562 22352
rect 2242 22272 2250 22336
rect 2314 22272 2330 22336
rect 2394 22272 2410 22336
rect 2474 22272 2490 22336
rect 2554 22272 2562 22336
rect 2242 21248 2562 22272
rect 2242 21184 2250 21248
rect 2314 21184 2330 21248
rect 2394 21184 2410 21248
rect 2474 21184 2490 21248
rect 2554 21184 2562 21248
rect 2242 20160 2562 21184
rect 2242 20096 2250 20160
rect 2314 20096 2330 20160
rect 2394 20096 2410 20160
rect 2474 20096 2490 20160
rect 2554 20096 2562 20160
rect 2242 19072 2562 20096
rect 2242 19008 2250 19072
rect 2314 19008 2330 19072
rect 2394 19008 2410 19072
rect 2474 19008 2490 19072
rect 2554 19008 2562 19072
rect 2242 17984 2562 19008
rect 2242 17920 2250 17984
rect 2314 17920 2330 17984
rect 2394 17920 2410 17984
rect 2474 17920 2490 17984
rect 2554 17920 2562 17984
rect 2242 16896 2562 17920
rect 2242 16832 2250 16896
rect 2314 16832 2330 16896
rect 2394 16832 2410 16896
rect 2474 16832 2490 16896
rect 2554 16832 2562 16896
rect 2242 15808 2562 16832
rect 2242 15744 2250 15808
rect 2314 15744 2330 15808
rect 2394 15744 2410 15808
rect 2474 15744 2490 15808
rect 2554 15744 2562 15808
rect 2242 14720 2562 15744
rect 2242 14656 2250 14720
rect 2314 14656 2330 14720
rect 2394 14656 2410 14720
rect 2474 14656 2490 14720
rect 2554 14656 2562 14720
rect 2242 13632 2562 14656
rect 2242 13568 2250 13632
rect 2314 13568 2330 13632
rect 2394 13568 2410 13632
rect 2474 13568 2490 13632
rect 2554 13568 2562 13632
rect 2242 12544 2562 13568
rect 2242 12480 2250 12544
rect 2314 12480 2330 12544
rect 2394 12480 2410 12544
rect 2474 12480 2490 12544
rect 2554 12480 2562 12544
rect 2242 11456 2562 12480
rect 2242 11392 2250 11456
rect 2314 11392 2330 11456
rect 2394 11392 2410 11456
rect 2474 11392 2490 11456
rect 2554 11392 2562 11456
rect 2242 10368 2562 11392
rect 2242 10304 2250 10368
rect 2314 10304 2330 10368
rect 2394 10304 2410 10368
rect 2474 10304 2490 10368
rect 2554 10304 2562 10368
rect 2242 9280 2562 10304
rect 2242 9216 2250 9280
rect 2314 9216 2330 9280
rect 2394 9216 2410 9280
rect 2474 9216 2490 9280
rect 2554 9216 2562 9280
rect 2242 8192 2562 9216
rect 2242 8128 2250 8192
rect 2314 8128 2330 8192
rect 2394 8128 2410 8192
rect 2474 8128 2490 8192
rect 2554 8128 2562 8192
rect 2242 7104 2562 8128
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2562 7104
rect 2242 6016 2562 7040
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2562 6016
rect 2242 4928 2562 5952
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2562 4928
rect 2242 3840 2562 4864
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2562 3840
rect 2242 2752 2562 3776
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2562 2752
rect 2242 2128 2562 2688
rect 3541 21792 3862 22352
rect 3541 21728 3549 21792
rect 3613 21728 3629 21792
rect 3693 21728 3709 21792
rect 3773 21728 3789 21792
rect 3853 21728 3862 21792
rect 3541 20704 3862 21728
rect 3541 20640 3549 20704
rect 3613 20640 3629 20704
rect 3693 20640 3709 20704
rect 3773 20640 3789 20704
rect 3853 20640 3862 20704
rect 3541 19616 3862 20640
rect 3541 19552 3549 19616
rect 3613 19552 3629 19616
rect 3693 19552 3709 19616
rect 3773 19552 3789 19616
rect 3853 19552 3862 19616
rect 3541 18528 3862 19552
rect 3541 18464 3549 18528
rect 3613 18464 3629 18528
rect 3693 18464 3709 18528
rect 3773 18464 3789 18528
rect 3853 18464 3862 18528
rect 3541 17440 3862 18464
rect 3541 17376 3549 17440
rect 3613 17376 3629 17440
rect 3693 17376 3709 17440
rect 3773 17376 3789 17440
rect 3853 17376 3862 17440
rect 3541 16352 3862 17376
rect 3541 16288 3549 16352
rect 3613 16288 3629 16352
rect 3693 16288 3709 16352
rect 3773 16288 3789 16352
rect 3853 16288 3862 16352
rect 3541 15264 3862 16288
rect 3541 15200 3549 15264
rect 3613 15200 3629 15264
rect 3693 15200 3709 15264
rect 3773 15200 3789 15264
rect 3853 15200 3862 15264
rect 3541 14176 3862 15200
rect 3541 14112 3549 14176
rect 3613 14112 3629 14176
rect 3693 14112 3709 14176
rect 3773 14112 3789 14176
rect 3853 14112 3862 14176
rect 3541 13088 3862 14112
rect 3541 13024 3549 13088
rect 3613 13024 3629 13088
rect 3693 13024 3709 13088
rect 3773 13024 3789 13088
rect 3853 13024 3862 13088
rect 3541 12000 3862 13024
rect 3541 11936 3549 12000
rect 3613 11936 3629 12000
rect 3693 11936 3709 12000
rect 3773 11936 3789 12000
rect 3853 11936 3862 12000
rect 3541 10912 3862 11936
rect 3541 10848 3549 10912
rect 3613 10848 3629 10912
rect 3693 10848 3709 10912
rect 3773 10848 3789 10912
rect 3853 10848 3862 10912
rect 3541 9824 3862 10848
rect 3541 9760 3549 9824
rect 3613 9760 3629 9824
rect 3693 9760 3709 9824
rect 3773 9760 3789 9824
rect 3853 9760 3862 9824
rect 3541 8736 3862 9760
rect 3541 8672 3549 8736
rect 3613 8672 3629 8736
rect 3693 8672 3709 8736
rect 3773 8672 3789 8736
rect 3853 8672 3862 8736
rect 3541 7648 3862 8672
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3862 7648
rect 3541 6560 3862 7584
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3862 6560
rect 3541 5472 3862 6496
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3862 5472
rect 3541 4384 3862 5408
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3862 4384
rect 3541 3296 3862 4320
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3862 3296
rect 3541 2208 3862 3232
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3862 2208
rect 3541 2128 3862 2144
rect 4840 22336 5160 22352
rect 4840 22272 4848 22336
rect 4912 22272 4928 22336
rect 4992 22272 5008 22336
rect 5072 22272 5088 22336
rect 5152 22272 5160 22336
rect 4840 21248 5160 22272
rect 4840 21184 4848 21248
rect 4912 21184 4928 21248
rect 4992 21184 5008 21248
rect 5072 21184 5088 21248
rect 5152 21184 5160 21248
rect 4840 20160 5160 21184
rect 4840 20096 4848 20160
rect 4912 20096 4928 20160
rect 4992 20096 5008 20160
rect 5072 20096 5088 20160
rect 5152 20096 5160 20160
rect 4840 19072 5160 20096
rect 4840 19008 4848 19072
rect 4912 19008 4928 19072
rect 4992 19008 5008 19072
rect 5072 19008 5088 19072
rect 5152 19008 5160 19072
rect 4840 17984 5160 19008
rect 4840 17920 4848 17984
rect 4912 17920 4928 17984
rect 4992 17920 5008 17984
rect 5072 17920 5088 17984
rect 5152 17920 5160 17984
rect 4840 16896 5160 17920
rect 4840 16832 4848 16896
rect 4912 16832 4928 16896
rect 4992 16832 5008 16896
rect 5072 16832 5088 16896
rect 5152 16832 5160 16896
rect 4840 15808 5160 16832
rect 4840 15744 4848 15808
rect 4912 15744 4928 15808
rect 4992 15744 5008 15808
rect 5072 15744 5088 15808
rect 5152 15744 5160 15808
rect 4840 14720 5160 15744
rect 4840 14656 4848 14720
rect 4912 14656 4928 14720
rect 4992 14656 5008 14720
rect 5072 14656 5088 14720
rect 5152 14656 5160 14720
rect 4840 13632 5160 14656
rect 4840 13568 4848 13632
rect 4912 13568 4928 13632
rect 4992 13568 5008 13632
rect 5072 13568 5088 13632
rect 5152 13568 5160 13632
rect 4840 12544 5160 13568
rect 4840 12480 4848 12544
rect 4912 12480 4928 12544
rect 4992 12480 5008 12544
rect 5072 12480 5088 12544
rect 5152 12480 5160 12544
rect 4840 11456 5160 12480
rect 4840 11392 4848 11456
rect 4912 11392 4928 11456
rect 4992 11392 5008 11456
rect 5072 11392 5088 11456
rect 5152 11392 5160 11456
rect 4840 10368 5160 11392
rect 4840 10304 4848 10368
rect 4912 10304 4928 10368
rect 4992 10304 5008 10368
rect 5072 10304 5088 10368
rect 5152 10304 5160 10368
rect 4840 9280 5160 10304
rect 4840 9216 4848 9280
rect 4912 9216 4928 9280
rect 4992 9216 5008 9280
rect 5072 9216 5088 9280
rect 5152 9216 5160 9280
rect 4840 8192 5160 9216
rect 4840 8128 4848 8192
rect 4912 8128 4928 8192
rect 4992 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5160 8192
rect 4840 7104 5160 8128
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 6016 5160 7040
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 4928 5160 5952
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 3840 5160 4864
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 2752 5160 3776
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2128 5160 2688
rect 6138 21792 6459 22352
rect 6138 21728 6146 21792
rect 6210 21728 6226 21792
rect 6290 21728 6306 21792
rect 6370 21728 6386 21792
rect 6450 21728 6459 21792
rect 6138 20704 6459 21728
rect 6138 20640 6146 20704
rect 6210 20640 6226 20704
rect 6290 20640 6306 20704
rect 6370 20640 6386 20704
rect 6450 20640 6459 20704
rect 6138 19616 6459 20640
rect 6138 19552 6146 19616
rect 6210 19552 6226 19616
rect 6290 19552 6306 19616
rect 6370 19552 6386 19616
rect 6450 19552 6459 19616
rect 6138 18528 6459 19552
rect 6138 18464 6146 18528
rect 6210 18464 6226 18528
rect 6290 18464 6306 18528
rect 6370 18464 6386 18528
rect 6450 18464 6459 18528
rect 6138 17440 6459 18464
rect 6138 17376 6146 17440
rect 6210 17376 6226 17440
rect 6290 17376 6306 17440
rect 6370 17376 6386 17440
rect 6450 17376 6459 17440
rect 6138 16352 6459 17376
rect 6138 16288 6146 16352
rect 6210 16288 6226 16352
rect 6290 16288 6306 16352
rect 6370 16288 6386 16352
rect 6450 16288 6459 16352
rect 6138 15264 6459 16288
rect 6138 15200 6146 15264
rect 6210 15200 6226 15264
rect 6290 15200 6306 15264
rect 6370 15200 6386 15264
rect 6450 15200 6459 15264
rect 6138 14176 6459 15200
rect 6138 14112 6146 14176
rect 6210 14112 6226 14176
rect 6290 14112 6306 14176
rect 6370 14112 6386 14176
rect 6450 14112 6459 14176
rect 6138 13088 6459 14112
rect 6138 13024 6146 13088
rect 6210 13024 6226 13088
rect 6290 13024 6306 13088
rect 6370 13024 6386 13088
rect 6450 13024 6459 13088
rect 6138 12000 6459 13024
rect 6138 11936 6146 12000
rect 6210 11936 6226 12000
rect 6290 11936 6306 12000
rect 6370 11936 6386 12000
rect 6450 11936 6459 12000
rect 6138 10912 6459 11936
rect 6138 10848 6146 10912
rect 6210 10848 6226 10912
rect 6290 10848 6306 10912
rect 6370 10848 6386 10912
rect 6450 10848 6459 10912
rect 6138 9824 6459 10848
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6459 9824
rect 6138 8736 6459 9760
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6459 8736
rect 6138 7648 6459 8672
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6459 7648
rect 6138 6560 6459 7584
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6459 6560
rect 6138 5472 6459 6496
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6459 5472
rect 6138 4384 6459 5408
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6459 4384
rect 6138 3296 6459 4320
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6459 3296
rect 6138 2208 6459 3232
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6459 2208
rect 6138 2128 6459 2144
rect 7437 22336 7757 22352
rect 7437 22272 7445 22336
rect 7509 22272 7525 22336
rect 7589 22272 7605 22336
rect 7669 22272 7685 22336
rect 7749 22272 7757 22336
rect 7437 21248 7757 22272
rect 7437 21184 7445 21248
rect 7509 21184 7525 21248
rect 7589 21184 7605 21248
rect 7669 21184 7685 21248
rect 7749 21184 7757 21248
rect 7437 20160 7757 21184
rect 7437 20096 7445 20160
rect 7509 20096 7525 20160
rect 7589 20096 7605 20160
rect 7669 20096 7685 20160
rect 7749 20096 7757 20160
rect 7437 19072 7757 20096
rect 7437 19008 7445 19072
rect 7509 19008 7525 19072
rect 7589 19008 7605 19072
rect 7669 19008 7685 19072
rect 7749 19008 7757 19072
rect 7437 17984 7757 19008
rect 7437 17920 7445 17984
rect 7509 17920 7525 17984
rect 7589 17920 7605 17984
rect 7669 17920 7685 17984
rect 7749 17920 7757 17984
rect 7437 16896 7757 17920
rect 7437 16832 7445 16896
rect 7509 16832 7525 16896
rect 7589 16832 7605 16896
rect 7669 16832 7685 16896
rect 7749 16832 7757 16896
rect 7437 15808 7757 16832
rect 7437 15744 7445 15808
rect 7509 15744 7525 15808
rect 7589 15744 7605 15808
rect 7669 15744 7685 15808
rect 7749 15744 7757 15808
rect 7437 14720 7757 15744
rect 7437 14656 7445 14720
rect 7509 14656 7525 14720
rect 7589 14656 7605 14720
rect 7669 14656 7685 14720
rect 7749 14656 7757 14720
rect 7437 13632 7757 14656
rect 7437 13568 7445 13632
rect 7509 13568 7525 13632
rect 7589 13568 7605 13632
rect 7669 13568 7685 13632
rect 7749 13568 7757 13632
rect 7437 12544 7757 13568
rect 7437 12480 7445 12544
rect 7509 12480 7525 12544
rect 7589 12480 7605 12544
rect 7669 12480 7685 12544
rect 7749 12480 7757 12544
rect 7437 11456 7757 12480
rect 7437 11392 7445 11456
rect 7509 11392 7525 11456
rect 7589 11392 7605 11456
rect 7669 11392 7685 11456
rect 7749 11392 7757 11456
rect 7437 10368 7757 11392
rect 7437 10304 7445 10368
rect 7509 10304 7525 10368
rect 7589 10304 7605 10368
rect 7669 10304 7685 10368
rect 7749 10304 7757 10368
rect 7437 9280 7757 10304
rect 7437 9216 7445 9280
rect 7509 9216 7525 9280
rect 7589 9216 7605 9280
rect 7669 9216 7685 9280
rect 7749 9216 7757 9280
rect 7437 8192 7757 9216
rect 7437 8128 7445 8192
rect 7509 8128 7525 8192
rect 7589 8128 7605 8192
rect 7669 8128 7685 8192
rect 7749 8128 7757 8192
rect 7437 7104 7757 8128
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 6016 7757 7040
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 7437 4928 7757 5952
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 7437 3840 7757 4864
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 7437 2752 7757 3776
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 7437 2128 7757 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1644511149
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1644511149
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_77
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1644511149
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 1644511149
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_77
timestamp 1644511149
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_73
timestamp 1644511149
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp 1644511149
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1644511149
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_73
timestamp 1644511149
transform 1 0 7820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_73
timestamp 1644511149
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1644511149
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1644511149
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1644511149
transform 1 0 7820 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 1644511149
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_77
timestamp 1644511149
transform 1 0 8188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 1644511149
transform 1 0 7820 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 1644511149
transform 1 0 7820 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_73
timestamp 1644511149
transform 1 0 7820 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1644511149
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp 1644511149
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1644511149
transform 1 0 8188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp 1644511149
transform 1 0 7820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1644511149
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1644511149
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1644511149
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1644511149
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_73
timestamp 1644511149
transform 1 0 7820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1644511149
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1644511149
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_73
timestamp 1644511149
transform 1 0 7820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_77
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_73
timestamp 1644511149
transform 1 0 7820 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_73
timestamp 1644511149
transform 1 0 7820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_77
timestamp 1644511149
transform 1 0 8188 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_73
timestamp 1644511149
transform 1 0 7820 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_65
timestamp 1644511149
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_70
timestamp 1644511149
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_77
timestamp 1644511149
transform 1 0 8188 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_73
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_73
timestamp 1644511149
transform 1 0 7820 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_77
timestamp 1644511149
transform 1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1644511149
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_63
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_70
timestamp 1644511149
transform 1 0 7544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_77
timestamp 1644511149
transform 1 0 8188 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_57
timestamp 1644511149
transform 1 0 6348 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1644511149
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1644511149
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 8832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 8832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 8832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 8832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 8832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _00__38 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _01__39
timestamp 1644511149
transform -1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _02__40
timestamp 1644511149
transform -1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _03__41
timestamp 1644511149
transform -1 0 8188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _04__42
timestamp 1644511149
transform -1 0 8188 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _05__43
timestamp 1644511149
transform -1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _06__44
timestamp 1644511149
transform -1 0 8188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _07__45
timestamp 1644511149
transform -1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _08__46
timestamp 1644511149
transform -1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _09__47
timestamp 1644511149
transform -1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _10__1
timestamp 1644511149
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _11__2
timestamp 1644511149
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _12__3
timestamp 1644511149
transform 1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _13__4
timestamp 1644511149
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _14__5
timestamp 1644511149
transform 1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _15__6
timestamp 1644511149
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _16__7
timestamp 1644511149
transform 1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _17__8
timestamp 1644511149
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18__9
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19__10
timestamp 1644511149
transform 1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20__11
timestamp 1644511149
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21__12
timestamp 1644511149
transform 1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22__13
timestamp 1644511149
transform 1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23__14
timestamp 1644511149
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24__15
timestamp 1644511149
transform 1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25__16
timestamp 1644511149
transform 1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26__17
timestamp 1644511149
transform 1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27__18
timestamp 1644511149
transform 1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28__19
timestamp 1644511149
transform 1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29__20
timestamp 1644511149
transform 1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30__21
timestamp 1644511149
transform 1 0 7268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31__22
timestamp 1644511149
transform 1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32__23
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33__24
timestamp 1644511149
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _34__25
timestamp 1644511149
transform 1 0 6624 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _35__26
timestamp 1644511149
transform 1 0 7268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _36__27
timestamp 1644511149
transform 1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37__28
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38__29
timestamp 1644511149
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39__30
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40__31
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _41__32
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _42__33
timestamp 1644511149
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _43__34
timestamp 1644511149
transform 1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44__35
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45__36
timestamp 1644511149
transform 1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _46__37
timestamp 1644511149
transform 1 0 7912 0 1 5440
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4986 0 5042 800 6 clk
port 0 nsew signal input
rlabel metal3 s 9200 144 10000 264 6 core0Index[0]
port 1 nsew signal tristate
rlabel metal3 s 9200 552 10000 672 6 core0Index[1]
port 2 nsew signal tristate
rlabel metal3 s 9200 1096 10000 1216 6 core0Index[2]
port 3 nsew signal tristate
rlabel metal3 s 9200 1640 10000 1760 6 core0Index[3]
port 4 nsew signal tristate
rlabel metal3 s 9200 2184 10000 2304 6 core0Index[4]
port 5 nsew signal tristate
rlabel metal3 s 9200 2728 10000 2848 6 core0Index[5]
port 6 nsew signal tristate
rlabel metal3 s 9200 3272 10000 3392 6 core0Index[6]
port 7 nsew signal tristate
rlabel metal3 s 9200 3816 10000 3936 6 core0Index[7]
port 8 nsew signal tristate
rlabel metal3 s 9200 4360 10000 4480 6 core1Index[0]
port 9 nsew signal tristate
rlabel metal3 s 9200 4904 10000 5024 6 core1Index[1]
port 10 nsew signal tristate
rlabel metal3 s 9200 5448 10000 5568 6 core1Index[2]
port 11 nsew signal tristate
rlabel metal3 s 9200 5992 10000 6112 6 core1Index[3]
port 12 nsew signal tristate
rlabel metal3 s 9200 6400 10000 6520 6 core1Index[4]
port 13 nsew signal tristate
rlabel metal3 s 9200 6944 10000 7064 6 core1Index[5]
port 14 nsew signal tristate
rlabel metal3 s 9200 7488 10000 7608 6 core1Index[6]
port 15 nsew signal tristate
rlabel metal3 s 9200 8032 10000 8152 6 core1Index[7]
port 16 nsew signal tristate
rlabel metal3 s 9200 8576 10000 8696 6 manufacturerID[0]
port 17 nsew signal tristate
rlabel metal3 s 9200 13880 10000 14000 6 manufacturerID[10]
port 18 nsew signal tristate
rlabel metal3 s 9200 9120 10000 9240 6 manufacturerID[1]
port 19 nsew signal tristate
rlabel metal3 s 9200 9664 10000 9784 6 manufacturerID[2]
port 20 nsew signal tristate
rlabel metal3 s 9200 10208 10000 10328 6 manufacturerID[3]
port 21 nsew signal tristate
rlabel metal3 s 9200 10752 10000 10872 6 manufacturerID[4]
port 22 nsew signal tristate
rlabel metal3 s 9200 11296 10000 11416 6 manufacturerID[5]
port 23 nsew signal tristate
rlabel metal3 s 9200 11840 10000 11960 6 manufacturerID[6]
port 24 nsew signal tristate
rlabel metal3 s 9200 12384 10000 12504 6 manufacturerID[7]
port 25 nsew signal tristate
rlabel metal3 s 9200 12792 10000 12912 6 manufacturerID[8]
port 26 nsew signal tristate
rlabel metal3 s 9200 13336 10000 13456 6 manufacturerID[9]
port 27 nsew signal tristate
rlabel metal3 s 9200 14424 10000 14544 6 partID[0]
port 28 nsew signal tristate
rlabel metal3 s 9200 19728 10000 19848 6 partID[10]
port 29 nsew signal tristate
rlabel metal3 s 9200 20272 10000 20392 6 partID[11]
port 30 nsew signal tristate
rlabel metal3 s 9200 20816 10000 20936 6 partID[12]
port 31 nsew signal tristate
rlabel metal3 s 9200 21360 10000 21480 6 partID[13]
port 32 nsew signal tristate
rlabel metal3 s 9200 21904 10000 22024 6 partID[14]
port 33 nsew signal tristate
rlabel metal3 s 9200 22448 10000 22568 6 partID[15]
port 34 nsew signal tristate
rlabel metal3 s 9200 14968 10000 15088 6 partID[1]
port 35 nsew signal tristate
rlabel metal3 s 9200 15512 10000 15632 6 partID[2]
port 36 nsew signal tristate
rlabel metal3 s 9200 16056 10000 16176 6 partID[3]
port 37 nsew signal tristate
rlabel metal3 s 9200 16600 10000 16720 6 partID[4]
port 38 nsew signal tristate
rlabel metal3 s 9200 17144 10000 17264 6 partID[5]
port 39 nsew signal tristate
rlabel metal3 s 9200 17688 10000 17808 6 partID[6]
port 40 nsew signal tristate
rlabel metal3 s 9200 18232 10000 18352 6 partID[7]
port 41 nsew signal tristate
rlabel metal3 s 9200 18776 10000 18896 6 partID[8]
port 42 nsew signal tristate
rlabel metal3 s 9200 19184 10000 19304 6 partID[9]
port 43 nsew signal tristate
rlabel metal4 s 2242 2128 2562 22352 6 vccd1
port 44 nsew power input
rlabel metal4 s 4840 2128 5160 22352 6 vccd1
port 44 nsew power input
rlabel metal4 s 7437 2128 7757 22352 6 vccd1
port 44 nsew power input
rlabel metal3 s 9200 22992 10000 23112 6 versionID[0]
port 45 nsew signal tristate
rlabel metal3 s 9200 23536 10000 23656 6 versionID[1]
port 46 nsew signal tristate
rlabel metal3 s 9200 24080 10000 24200 6 versionID[2]
port 47 nsew signal tristate
rlabel metal3 s 9200 24624 10000 24744 6 versionID[3]
port 48 nsew signal tristate
rlabel metal4 s 3542 2128 3862 22352 6 vssd1
port 49 nsew ground input
rlabel metal4 s 6139 2128 6459 22352 6 vssd1
port 49 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 10000 25000
<< end >>
