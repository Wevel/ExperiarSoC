magic
tech sky130A
magscale 1 2
timestamp 1654449317
<< obsli1 >>
rect 1104 2159 98808 197489
<< obsm1 >>
rect 566 1300 99990 197520
<< metal2 >>
rect 1214 199200 1270 200000
rect 3698 199200 3754 200000
rect 6274 199200 6330 200000
rect 8850 199200 8906 200000
rect 11426 199200 11482 200000
rect 14002 199200 14058 200000
rect 16578 199200 16634 200000
rect 19154 199200 19210 200000
rect 21638 199200 21694 200000
rect 24214 199200 24270 200000
rect 26790 199200 26846 200000
rect 29366 199200 29422 200000
rect 31942 199200 31998 200000
rect 34518 199200 34574 200000
rect 37094 199200 37150 200000
rect 39670 199200 39726 200000
rect 42154 199200 42210 200000
rect 44730 199200 44786 200000
rect 47306 199200 47362 200000
rect 49882 199200 49938 200000
rect 52458 199200 52514 200000
rect 55034 199200 55090 200000
rect 57610 199200 57666 200000
rect 60186 199200 60242 200000
rect 62670 199200 62726 200000
rect 65246 199200 65302 200000
rect 67822 199200 67878 200000
rect 70398 199200 70454 200000
rect 72974 199200 73030 200000
rect 75550 199200 75606 200000
rect 78126 199200 78182 200000
rect 80702 199200 80758 200000
rect 83186 199200 83242 200000
rect 85762 199200 85818 200000
rect 88338 199200 88394 200000
rect 90914 199200 90970 200000
rect 93490 199200 93546 200000
rect 96066 199200 96122 200000
rect 98642 199200 98698 200000
rect 662 0 718 800
rect 2042 0 2098 800
rect 3422 0 3478 800
rect 4802 0 4858 800
rect 6274 0 6330 800
rect 7654 0 7710 800
rect 9034 0 9090 800
rect 10506 0 10562 800
rect 11886 0 11942 800
rect 13266 0 13322 800
rect 14738 0 14794 800
rect 16118 0 16174 800
rect 17498 0 17554 800
rect 18970 0 19026 800
rect 20350 0 20406 800
rect 21730 0 21786 800
rect 23110 0 23166 800
rect 24582 0 24638 800
rect 25962 0 26018 800
rect 27342 0 27398 800
rect 28814 0 28870 800
rect 30194 0 30250 800
rect 31574 0 31630 800
rect 33046 0 33102 800
rect 34426 0 34482 800
rect 35806 0 35862 800
rect 37278 0 37334 800
rect 38658 0 38714 800
rect 40038 0 40094 800
rect 41418 0 41474 800
rect 42890 0 42946 800
rect 44270 0 44326 800
rect 45650 0 45706 800
rect 47122 0 47178 800
rect 48502 0 48558 800
rect 49882 0 49938 800
rect 51354 0 51410 800
rect 52734 0 52790 800
rect 54114 0 54170 800
rect 55586 0 55642 800
rect 56966 0 57022 800
rect 58346 0 58402 800
rect 59818 0 59874 800
rect 61198 0 61254 800
rect 62578 0 62634 800
rect 63958 0 64014 800
rect 65430 0 65486 800
rect 66810 0 66866 800
rect 68190 0 68246 800
rect 69662 0 69718 800
rect 71042 0 71098 800
rect 72422 0 72478 800
rect 73894 0 73950 800
rect 75274 0 75330 800
rect 76654 0 76710 800
rect 78126 0 78182 800
rect 79506 0 79562 800
rect 80886 0 80942 800
rect 82266 0 82322 800
rect 83738 0 83794 800
rect 85118 0 85174 800
rect 86498 0 86554 800
rect 87970 0 88026 800
rect 89350 0 89406 800
rect 90730 0 90786 800
rect 92202 0 92258 800
rect 93582 0 93638 800
rect 94962 0 95018 800
rect 96434 0 96490 800
rect 97814 0 97870 800
rect 99194 0 99250 800
<< obsm2 >>
rect 572 199144 1158 199481
rect 1326 199144 3642 199481
rect 3810 199144 6218 199481
rect 6386 199144 8794 199481
rect 8962 199144 11370 199481
rect 11538 199144 13946 199481
rect 14114 199144 16522 199481
rect 16690 199144 19098 199481
rect 19266 199144 21582 199481
rect 21750 199144 24158 199481
rect 24326 199144 26734 199481
rect 26902 199144 29310 199481
rect 29478 199144 31886 199481
rect 32054 199144 34462 199481
rect 34630 199144 37038 199481
rect 37206 199144 39614 199481
rect 39782 199144 42098 199481
rect 42266 199144 44674 199481
rect 44842 199144 47250 199481
rect 47418 199144 49826 199481
rect 49994 199144 52402 199481
rect 52570 199144 54978 199481
rect 55146 199144 57554 199481
rect 57722 199144 60130 199481
rect 60298 199144 62614 199481
rect 62782 199144 65190 199481
rect 65358 199144 67766 199481
rect 67934 199144 70342 199481
rect 70510 199144 72918 199481
rect 73086 199144 75494 199481
rect 75662 199144 78070 199481
rect 78238 199144 80646 199481
rect 80814 199144 83130 199481
rect 83298 199144 85706 199481
rect 85874 199144 88282 199481
rect 88450 199144 90858 199481
rect 91026 199144 93434 199481
rect 93602 199144 96010 199481
rect 96178 199144 98586 199481
rect 98754 199144 99986 199481
rect 572 856 99986 199144
rect 572 439 606 856
rect 774 439 1986 856
rect 2154 439 3366 856
rect 3534 439 4746 856
rect 4914 439 6218 856
rect 6386 439 7598 856
rect 7766 439 8978 856
rect 9146 439 10450 856
rect 10618 439 11830 856
rect 11998 439 13210 856
rect 13378 439 14682 856
rect 14850 439 16062 856
rect 16230 439 17442 856
rect 17610 439 18914 856
rect 19082 439 20294 856
rect 20462 439 21674 856
rect 21842 439 23054 856
rect 23222 439 24526 856
rect 24694 439 25906 856
rect 26074 439 27286 856
rect 27454 439 28758 856
rect 28926 439 30138 856
rect 30306 439 31518 856
rect 31686 439 32990 856
rect 33158 439 34370 856
rect 34538 439 35750 856
rect 35918 439 37222 856
rect 37390 439 38602 856
rect 38770 439 39982 856
rect 40150 439 41362 856
rect 41530 439 42834 856
rect 43002 439 44214 856
rect 44382 439 45594 856
rect 45762 439 47066 856
rect 47234 439 48446 856
rect 48614 439 49826 856
rect 49994 439 51298 856
rect 51466 439 52678 856
rect 52846 439 54058 856
rect 54226 439 55530 856
rect 55698 439 56910 856
rect 57078 439 58290 856
rect 58458 439 59762 856
rect 59930 439 61142 856
rect 61310 439 62522 856
rect 62690 439 63902 856
rect 64070 439 65374 856
rect 65542 439 66754 856
rect 66922 439 68134 856
rect 68302 439 69606 856
rect 69774 439 70986 856
rect 71154 439 72366 856
rect 72534 439 73838 856
rect 74006 439 75218 856
rect 75386 439 76598 856
rect 76766 439 78070 856
rect 78238 439 79450 856
rect 79618 439 80830 856
rect 80998 439 82210 856
rect 82378 439 83682 856
rect 83850 439 85062 856
rect 85230 439 86442 856
rect 86610 439 87914 856
rect 88082 439 89294 856
rect 89462 439 90674 856
rect 90842 439 92146 856
rect 92314 439 93526 856
rect 93694 439 94906 856
rect 95074 439 96378 856
rect 96546 439 97758 856
rect 97926 439 99138 856
rect 99306 439 99986 856
<< metal3 >>
rect 0 199384 800 199504
rect 99200 199384 100000 199504
rect 0 198296 800 198416
rect 99200 198432 100000 198552
rect 0 197344 800 197464
rect 99200 197480 100000 197600
rect 0 196256 800 196376
rect 99200 196392 100000 196512
rect 99200 195440 100000 195560
rect 0 195168 800 195288
rect 99200 194488 100000 194608
rect 0 194216 800 194336
rect 99200 193536 100000 193656
rect 0 193128 800 193248
rect 99200 192448 100000 192568
rect 0 192176 800 192296
rect 99200 191496 100000 191616
rect 0 191088 800 191208
rect 99200 190544 100000 190664
rect 0 190000 800 190120
rect 99200 189456 100000 189576
rect 0 189048 800 189168
rect 99200 188504 100000 188624
rect 0 187960 800 188080
rect 99200 187552 100000 187672
rect 0 186872 800 186992
rect 99200 186600 100000 186720
rect 0 185920 800 186040
rect 99200 185512 100000 185632
rect 0 184832 800 184952
rect 99200 184560 100000 184680
rect 0 183880 800 184000
rect 99200 183608 100000 183728
rect 0 182792 800 182912
rect 99200 182520 100000 182640
rect 0 181704 800 181824
rect 99200 181568 100000 181688
rect 0 180752 800 180872
rect 99200 180616 100000 180736
rect 0 179664 800 179784
rect 99200 179664 100000 179784
rect 0 178576 800 178696
rect 99200 178576 100000 178696
rect 0 177624 800 177744
rect 99200 177624 100000 177744
rect 0 176536 800 176656
rect 99200 176672 100000 176792
rect 0 175584 800 175704
rect 99200 175584 100000 175704
rect 0 174496 800 174616
rect 99200 174632 100000 174752
rect 99200 173680 100000 173800
rect 0 173408 800 173528
rect 99200 172728 100000 172848
rect 0 172456 800 172576
rect 99200 171640 100000 171760
rect 0 171368 800 171488
rect 99200 170688 100000 170808
rect 0 170280 800 170400
rect 99200 169736 100000 169856
rect 0 169328 800 169448
rect 99200 168648 100000 168768
rect 0 168240 800 168360
rect 99200 167696 100000 167816
rect 0 167288 800 167408
rect 99200 166744 100000 166864
rect 0 166200 800 166320
rect 99200 165792 100000 165912
rect 0 165112 800 165232
rect 99200 164704 100000 164824
rect 0 164160 800 164280
rect 99200 163752 100000 163872
rect 0 163072 800 163192
rect 99200 162800 100000 162920
rect 0 161984 800 162104
rect 99200 161712 100000 161832
rect 0 161032 800 161152
rect 99200 160760 100000 160880
rect 0 159944 800 160064
rect 99200 159808 100000 159928
rect 0 158992 800 159112
rect 99200 158856 100000 158976
rect 0 157904 800 158024
rect 99200 157768 100000 157888
rect 0 156816 800 156936
rect 99200 156816 100000 156936
rect 0 155864 800 155984
rect 99200 155864 100000 155984
rect 0 154776 800 154896
rect 99200 154912 100000 155032
rect 0 153824 800 153944
rect 99200 153824 100000 153944
rect 0 152736 800 152856
rect 99200 152872 100000 152992
rect 99200 151920 100000 152040
rect 0 151648 800 151768
rect 0 150696 800 150816
rect 99200 150832 100000 150952
rect 99200 149880 100000 150000
rect 0 149608 800 149728
rect 99200 148928 100000 149048
rect 0 148520 800 148640
rect 99200 147976 100000 148096
rect 0 147568 800 147688
rect 99200 146888 100000 147008
rect 0 146480 800 146600
rect 99200 145936 100000 146056
rect 0 145528 800 145648
rect 99200 144984 100000 145104
rect 0 144440 800 144560
rect 99200 143896 100000 144016
rect 0 143352 800 143472
rect 99200 142944 100000 143064
rect 0 142400 800 142520
rect 99200 141992 100000 142112
rect 0 141312 800 141432
rect 99200 141040 100000 141160
rect 0 140224 800 140344
rect 99200 139952 100000 140072
rect 0 139272 800 139392
rect 99200 139000 100000 139120
rect 0 138184 800 138304
rect 99200 138048 100000 138168
rect 0 137232 800 137352
rect 99200 136960 100000 137080
rect 0 136144 800 136264
rect 99200 136008 100000 136128
rect 0 135056 800 135176
rect 99200 135056 100000 135176
rect 0 134104 800 134224
rect 99200 134104 100000 134224
rect 0 133016 800 133136
rect 99200 133016 100000 133136
rect 0 131928 800 132048
rect 99200 132064 100000 132184
rect 0 130976 800 131096
rect 99200 131112 100000 131232
rect 0 129888 800 130008
rect 99200 130024 100000 130144
rect 0 128936 800 129056
rect 99200 129072 100000 129192
rect 99200 128120 100000 128240
rect 0 127848 800 127968
rect 99200 127168 100000 127288
rect 0 126760 800 126880
rect 99200 126080 100000 126200
rect 0 125808 800 125928
rect 99200 125128 100000 125248
rect 0 124720 800 124840
rect 99200 124176 100000 124296
rect 0 123632 800 123752
rect 99200 123088 100000 123208
rect 0 122680 800 122800
rect 99200 122136 100000 122256
rect 0 121592 800 121712
rect 99200 121184 100000 121304
rect 0 120640 800 120760
rect 99200 120232 100000 120352
rect 0 119552 800 119672
rect 99200 119144 100000 119264
rect 0 118464 800 118584
rect 99200 118192 100000 118312
rect 0 117512 800 117632
rect 99200 117240 100000 117360
rect 0 116424 800 116544
rect 99200 116288 100000 116408
rect 0 115472 800 115592
rect 99200 115200 100000 115320
rect 0 114384 800 114504
rect 99200 114248 100000 114368
rect 0 113296 800 113416
rect 99200 113296 100000 113416
rect 0 112344 800 112464
rect 99200 112208 100000 112328
rect 0 111256 800 111376
rect 99200 111256 100000 111376
rect 0 110168 800 110288
rect 99200 110304 100000 110424
rect 0 109216 800 109336
rect 99200 109352 100000 109472
rect 0 108128 800 108248
rect 99200 108264 100000 108384
rect 0 107176 800 107296
rect 99200 107312 100000 107432
rect 99200 106360 100000 106480
rect 0 106088 800 106208
rect 99200 105272 100000 105392
rect 0 105000 800 105120
rect 99200 104320 100000 104440
rect 0 104048 800 104168
rect 99200 103368 100000 103488
rect 0 102960 800 103080
rect 99200 102416 100000 102536
rect 0 101872 800 101992
rect 99200 101328 100000 101448
rect 0 100920 800 101040
rect 99200 100376 100000 100496
rect 0 99832 800 99952
rect 99200 99424 100000 99544
rect 0 98880 800 99000
rect 99200 98336 100000 98456
rect 0 97792 800 97912
rect 99200 97384 100000 97504
rect 0 96704 800 96824
rect 99200 96432 100000 96552
rect 0 95752 800 95872
rect 99200 95480 100000 95600
rect 0 94664 800 94784
rect 99200 94392 100000 94512
rect 0 93576 800 93696
rect 99200 93440 100000 93560
rect 0 92624 800 92744
rect 99200 92488 100000 92608
rect 0 91536 800 91656
rect 99200 91400 100000 91520
rect 0 90584 800 90704
rect 99200 90448 100000 90568
rect 0 89496 800 89616
rect 99200 89496 100000 89616
rect 0 88408 800 88528
rect 99200 88544 100000 88664
rect 0 87456 800 87576
rect 99200 87456 100000 87576
rect 0 86368 800 86488
rect 99200 86504 100000 86624
rect 99200 85552 100000 85672
rect 0 85280 800 85400
rect 0 84328 800 84448
rect 99200 84464 100000 84584
rect 99200 83512 100000 83632
rect 0 83240 800 83360
rect 99200 82560 100000 82680
rect 0 82288 800 82408
rect 99200 81608 100000 81728
rect 0 81200 800 81320
rect 99200 80520 100000 80640
rect 0 80112 800 80232
rect 99200 79568 100000 79688
rect 0 79160 800 79280
rect 99200 78616 100000 78736
rect 0 78072 800 78192
rect 99200 77664 100000 77784
rect 0 77120 800 77240
rect 99200 76576 100000 76696
rect 0 76032 800 76152
rect 99200 75624 100000 75744
rect 0 74944 800 75064
rect 99200 74672 100000 74792
rect 0 73992 800 74112
rect 99200 73584 100000 73704
rect 0 72904 800 73024
rect 99200 72632 100000 72752
rect 0 71816 800 71936
rect 99200 71680 100000 71800
rect 0 70864 800 70984
rect 99200 70728 100000 70848
rect 0 69776 800 69896
rect 99200 69640 100000 69760
rect 0 68824 800 68944
rect 99200 68688 100000 68808
rect 0 67736 800 67856
rect 99200 67736 100000 67856
rect 0 66648 800 66768
rect 99200 66648 100000 66768
rect 0 65696 800 65816
rect 99200 65696 100000 65816
rect 0 64608 800 64728
rect 99200 64744 100000 64864
rect 99200 63792 100000 63912
rect 0 63520 800 63640
rect 0 62568 800 62688
rect 99200 62704 100000 62824
rect 99200 61752 100000 61872
rect 0 61480 800 61600
rect 99200 60800 100000 60920
rect 0 60528 800 60648
rect 99200 59712 100000 59832
rect 0 59440 800 59560
rect 99200 58760 100000 58880
rect 0 58352 800 58472
rect 99200 57808 100000 57928
rect 0 57400 800 57520
rect 99200 56856 100000 56976
rect 0 56312 800 56432
rect 99200 55768 100000 55888
rect 0 55224 800 55344
rect 99200 54816 100000 54936
rect 0 54272 800 54392
rect 99200 53864 100000 53984
rect 0 53184 800 53304
rect 99200 52776 100000 52896
rect 0 52232 800 52352
rect 99200 51824 100000 51944
rect 0 51144 800 51264
rect 99200 50872 100000 50992
rect 0 50056 800 50176
rect 99200 49920 100000 50040
rect 0 49104 800 49224
rect 99200 48832 100000 48952
rect 0 48016 800 48136
rect 99200 47880 100000 48000
rect 0 46928 800 47048
rect 99200 46928 100000 47048
rect 0 45976 800 46096
rect 99200 45840 100000 45960
rect 0 44888 800 45008
rect 99200 44888 100000 45008
rect 0 43936 800 44056
rect 99200 43936 100000 44056
rect 0 42848 800 42968
rect 99200 42984 100000 43104
rect 0 41760 800 41880
rect 99200 41896 100000 42016
rect 0 40808 800 40928
rect 99200 40944 100000 41064
rect 99200 39992 100000 40112
rect 0 39720 800 39840
rect 99200 39040 100000 39160
rect 0 38768 800 38888
rect 99200 37952 100000 38072
rect 0 37680 800 37800
rect 99200 37000 100000 37120
rect 0 36592 800 36712
rect 99200 36048 100000 36168
rect 0 35640 800 35760
rect 99200 34960 100000 35080
rect 0 34552 800 34672
rect 99200 34008 100000 34128
rect 0 33464 800 33584
rect 99200 33056 100000 33176
rect 0 32512 800 32632
rect 99200 32104 100000 32224
rect 0 31424 800 31544
rect 99200 31016 100000 31136
rect 0 30472 800 30592
rect 99200 30064 100000 30184
rect 0 29384 800 29504
rect 99200 29112 100000 29232
rect 0 28296 800 28416
rect 99200 28024 100000 28144
rect 0 27344 800 27464
rect 99200 27072 100000 27192
rect 0 26256 800 26376
rect 99200 26120 100000 26240
rect 0 25168 800 25288
rect 99200 25168 100000 25288
rect 0 24216 800 24336
rect 99200 24080 100000 24200
rect 0 23128 800 23248
rect 99200 23128 100000 23248
rect 0 22176 800 22296
rect 99200 22176 100000 22296
rect 0 21088 800 21208
rect 99200 21088 100000 21208
rect 0 20000 800 20120
rect 99200 20136 100000 20256
rect 0 19048 800 19168
rect 99200 19184 100000 19304
rect 99200 18232 100000 18352
rect 0 17960 800 18080
rect 99200 17144 100000 17264
rect 0 16872 800 16992
rect 99200 16192 100000 16312
rect 0 15920 800 16040
rect 99200 15240 100000 15360
rect 0 14832 800 14952
rect 99200 14152 100000 14272
rect 0 13880 800 14000
rect 99200 13200 100000 13320
rect 0 12792 800 12912
rect 99200 12248 100000 12368
rect 0 11704 800 11824
rect 99200 11296 100000 11416
rect 0 10752 800 10872
rect 99200 10208 100000 10328
rect 0 9664 800 9784
rect 99200 9256 100000 9376
rect 0 8576 800 8696
rect 99200 8304 100000 8424
rect 0 7624 800 7744
rect 99200 7216 100000 7336
rect 0 6536 800 6656
rect 99200 6264 100000 6384
rect 0 5584 800 5704
rect 99200 5312 100000 5432
rect 0 4496 800 4616
rect 99200 4360 100000 4480
rect 0 3408 800 3528
rect 99200 3272 100000 3392
rect 0 2456 800 2576
rect 99200 2320 100000 2440
rect 0 1368 800 1488
rect 99200 1368 100000 1488
rect 0 416 800 536
rect 99200 416 100000 536
<< obsm3 >>
rect 880 199304 99120 199477
rect 657 198632 99991 199304
rect 657 198496 99120 198632
rect 880 198352 99120 198496
rect 880 198216 99991 198352
rect 657 197680 99991 198216
rect 657 197544 99120 197680
rect 880 197400 99120 197544
rect 880 197264 99991 197400
rect 657 196592 99991 197264
rect 657 196456 99120 196592
rect 880 196312 99120 196456
rect 880 196176 99991 196312
rect 657 195640 99991 196176
rect 657 195368 99120 195640
rect 880 195360 99120 195368
rect 880 195088 99991 195360
rect 657 194688 99991 195088
rect 657 194416 99120 194688
rect 880 194408 99120 194416
rect 880 194136 99991 194408
rect 657 193736 99991 194136
rect 657 193456 99120 193736
rect 657 193328 99991 193456
rect 880 193048 99991 193328
rect 657 192648 99991 193048
rect 657 192376 99120 192648
rect 880 192368 99120 192376
rect 880 192096 99991 192368
rect 657 191696 99991 192096
rect 657 191416 99120 191696
rect 657 191288 99991 191416
rect 880 191008 99991 191288
rect 657 190744 99991 191008
rect 657 190464 99120 190744
rect 657 190200 99991 190464
rect 880 189920 99991 190200
rect 657 189656 99991 189920
rect 657 189376 99120 189656
rect 657 189248 99991 189376
rect 880 188968 99991 189248
rect 657 188704 99991 188968
rect 657 188424 99120 188704
rect 657 188160 99991 188424
rect 880 187880 99991 188160
rect 657 187752 99991 187880
rect 657 187472 99120 187752
rect 657 187072 99991 187472
rect 880 186800 99991 187072
rect 880 186792 99120 186800
rect 657 186520 99120 186792
rect 657 186120 99991 186520
rect 880 185840 99991 186120
rect 657 185712 99991 185840
rect 657 185432 99120 185712
rect 657 185032 99991 185432
rect 880 184760 99991 185032
rect 880 184752 99120 184760
rect 657 184480 99120 184752
rect 657 184080 99991 184480
rect 880 183808 99991 184080
rect 880 183800 99120 183808
rect 657 183528 99120 183800
rect 657 182992 99991 183528
rect 880 182720 99991 182992
rect 880 182712 99120 182720
rect 657 182440 99120 182712
rect 657 181904 99991 182440
rect 880 181768 99991 181904
rect 880 181624 99120 181768
rect 657 181488 99120 181624
rect 657 180952 99991 181488
rect 880 180816 99991 180952
rect 880 180672 99120 180816
rect 657 180536 99120 180672
rect 657 179864 99991 180536
rect 880 179584 99120 179864
rect 657 178776 99991 179584
rect 880 178496 99120 178776
rect 657 177824 99991 178496
rect 880 177544 99120 177824
rect 657 176872 99991 177544
rect 657 176736 99120 176872
rect 880 176592 99120 176736
rect 880 176456 99991 176592
rect 657 175784 99991 176456
rect 880 175504 99120 175784
rect 657 174832 99991 175504
rect 657 174696 99120 174832
rect 880 174552 99120 174696
rect 880 174416 99991 174552
rect 657 173880 99991 174416
rect 657 173608 99120 173880
rect 880 173600 99120 173608
rect 880 173328 99991 173600
rect 657 172928 99991 173328
rect 657 172656 99120 172928
rect 880 172648 99120 172656
rect 880 172376 99991 172648
rect 657 171840 99991 172376
rect 657 171568 99120 171840
rect 880 171560 99120 171568
rect 880 171288 99991 171560
rect 657 170888 99991 171288
rect 657 170608 99120 170888
rect 657 170480 99991 170608
rect 880 170200 99991 170480
rect 657 169936 99991 170200
rect 657 169656 99120 169936
rect 657 169528 99991 169656
rect 880 169248 99991 169528
rect 657 168848 99991 169248
rect 657 168568 99120 168848
rect 657 168440 99991 168568
rect 880 168160 99991 168440
rect 657 167896 99991 168160
rect 657 167616 99120 167896
rect 657 167488 99991 167616
rect 880 167208 99991 167488
rect 657 166944 99991 167208
rect 657 166664 99120 166944
rect 657 166400 99991 166664
rect 880 166120 99991 166400
rect 657 165992 99991 166120
rect 657 165712 99120 165992
rect 657 165312 99991 165712
rect 880 165032 99991 165312
rect 657 164904 99991 165032
rect 657 164624 99120 164904
rect 657 164360 99991 164624
rect 880 164080 99991 164360
rect 657 163952 99991 164080
rect 657 163672 99120 163952
rect 657 163272 99991 163672
rect 880 163000 99991 163272
rect 880 162992 99120 163000
rect 657 162720 99120 162992
rect 657 162184 99991 162720
rect 880 161912 99991 162184
rect 880 161904 99120 161912
rect 657 161632 99120 161904
rect 657 161232 99991 161632
rect 880 160960 99991 161232
rect 880 160952 99120 160960
rect 657 160680 99120 160952
rect 657 160144 99991 160680
rect 880 160008 99991 160144
rect 880 159864 99120 160008
rect 657 159728 99120 159864
rect 657 159192 99991 159728
rect 880 159056 99991 159192
rect 880 158912 99120 159056
rect 657 158776 99120 158912
rect 657 158104 99991 158776
rect 880 157968 99991 158104
rect 880 157824 99120 157968
rect 657 157688 99120 157824
rect 657 157016 99991 157688
rect 880 156736 99120 157016
rect 657 156064 99991 156736
rect 880 155784 99120 156064
rect 657 155112 99991 155784
rect 657 154976 99120 155112
rect 880 154832 99120 154976
rect 880 154696 99991 154832
rect 657 154024 99991 154696
rect 880 153744 99120 154024
rect 657 153072 99991 153744
rect 657 152936 99120 153072
rect 880 152792 99120 152936
rect 880 152656 99991 152792
rect 657 152120 99991 152656
rect 657 151848 99120 152120
rect 880 151840 99120 151848
rect 880 151568 99991 151840
rect 657 151032 99991 151568
rect 657 150896 99120 151032
rect 880 150752 99120 150896
rect 880 150616 99991 150752
rect 657 150080 99991 150616
rect 657 149808 99120 150080
rect 880 149800 99120 149808
rect 880 149528 99991 149800
rect 657 149128 99991 149528
rect 657 148848 99120 149128
rect 657 148720 99991 148848
rect 880 148440 99991 148720
rect 657 148176 99991 148440
rect 657 147896 99120 148176
rect 657 147768 99991 147896
rect 880 147488 99991 147768
rect 657 147088 99991 147488
rect 657 146808 99120 147088
rect 657 146680 99991 146808
rect 880 146400 99991 146680
rect 657 146136 99991 146400
rect 657 145856 99120 146136
rect 657 145728 99991 145856
rect 880 145448 99991 145728
rect 657 145184 99991 145448
rect 657 144904 99120 145184
rect 657 144640 99991 144904
rect 880 144360 99991 144640
rect 657 144096 99991 144360
rect 657 143816 99120 144096
rect 657 143552 99991 143816
rect 880 143272 99991 143552
rect 657 143144 99991 143272
rect 657 142864 99120 143144
rect 657 142600 99991 142864
rect 880 142320 99991 142600
rect 657 142192 99991 142320
rect 657 141912 99120 142192
rect 657 141512 99991 141912
rect 880 141240 99991 141512
rect 880 141232 99120 141240
rect 657 140960 99120 141232
rect 657 140424 99991 140960
rect 880 140152 99991 140424
rect 880 140144 99120 140152
rect 657 139872 99120 140144
rect 657 139472 99991 139872
rect 880 139200 99991 139472
rect 880 139192 99120 139200
rect 657 138920 99120 139192
rect 657 138384 99991 138920
rect 880 138248 99991 138384
rect 880 138104 99120 138248
rect 657 137968 99120 138104
rect 657 137432 99991 137968
rect 880 137160 99991 137432
rect 880 137152 99120 137160
rect 657 136880 99120 137152
rect 657 136344 99991 136880
rect 880 136208 99991 136344
rect 880 136064 99120 136208
rect 657 135928 99120 136064
rect 657 135256 99991 135928
rect 880 134976 99120 135256
rect 657 134304 99991 134976
rect 880 134024 99120 134304
rect 657 133216 99991 134024
rect 880 132936 99120 133216
rect 657 132264 99991 132936
rect 657 132128 99120 132264
rect 880 131984 99120 132128
rect 880 131848 99991 131984
rect 657 131312 99991 131848
rect 657 131176 99120 131312
rect 880 131032 99120 131176
rect 880 130896 99991 131032
rect 657 130224 99991 130896
rect 657 130088 99120 130224
rect 880 129944 99120 130088
rect 880 129808 99991 129944
rect 657 129272 99991 129808
rect 657 129136 99120 129272
rect 880 128992 99120 129136
rect 880 128856 99991 128992
rect 657 128320 99991 128856
rect 657 128048 99120 128320
rect 880 128040 99120 128048
rect 880 127768 99991 128040
rect 657 127368 99991 127768
rect 657 127088 99120 127368
rect 657 126960 99991 127088
rect 880 126680 99991 126960
rect 657 126280 99991 126680
rect 657 126008 99120 126280
rect 880 126000 99120 126008
rect 880 125728 99991 126000
rect 657 125328 99991 125728
rect 657 125048 99120 125328
rect 657 124920 99991 125048
rect 880 124640 99991 124920
rect 657 124376 99991 124640
rect 657 124096 99120 124376
rect 657 123832 99991 124096
rect 880 123552 99991 123832
rect 657 123288 99991 123552
rect 657 123008 99120 123288
rect 657 122880 99991 123008
rect 880 122600 99991 122880
rect 657 122336 99991 122600
rect 657 122056 99120 122336
rect 657 121792 99991 122056
rect 880 121512 99991 121792
rect 657 121384 99991 121512
rect 657 121104 99120 121384
rect 657 120840 99991 121104
rect 880 120560 99991 120840
rect 657 120432 99991 120560
rect 657 120152 99120 120432
rect 657 119752 99991 120152
rect 880 119472 99991 119752
rect 657 119344 99991 119472
rect 657 119064 99120 119344
rect 657 118664 99991 119064
rect 880 118392 99991 118664
rect 880 118384 99120 118392
rect 657 118112 99120 118384
rect 657 117712 99991 118112
rect 880 117440 99991 117712
rect 880 117432 99120 117440
rect 657 117160 99120 117432
rect 657 116624 99991 117160
rect 880 116488 99991 116624
rect 880 116344 99120 116488
rect 657 116208 99120 116344
rect 657 115672 99991 116208
rect 880 115400 99991 115672
rect 880 115392 99120 115400
rect 657 115120 99120 115392
rect 657 114584 99991 115120
rect 880 114448 99991 114584
rect 880 114304 99120 114448
rect 657 114168 99120 114304
rect 657 113496 99991 114168
rect 880 113216 99120 113496
rect 657 112544 99991 113216
rect 880 112408 99991 112544
rect 880 112264 99120 112408
rect 657 112128 99120 112264
rect 657 111456 99991 112128
rect 880 111176 99120 111456
rect 657 110504 99991 111176
rect 657 110368 99120 110504
rect 880 110224 99120 110368
rect 880 110088 99991 110224
rect 657 109552 99991 110088
rect 657 109416 99120 109552
rect 880 109272 99120 109416
rect 880 109136 99991 109272
rect 657 108464 99991 109136
rect 657 108328 99120 108464
rect 880 108184 99120 108328
rect 880 108048 99991 108184
rect 657 107512 99991 108048
rect 657 107376 99120 107512
rect 880 107232 99120 107376
rect 880 107096 99991 107232
rect 657 106560 99991 107096
rect 657 106288 99120 106560
rect 880 106280 99120 106288
rect 880 106008 99991 106280
rect 657 105472 99991 106008
rect 657 105200 99120 105472
rect 880 105192 99120 105200
rect 880 104920 99991 105192
rect 657 104520 99991 104920
rect 657 104248 99120 104520
rect 880 104240 99120 104248
rect 880 103968 99991 104240
rect 657 103568 99991 103968
rect 657 103288 99120 103568
rect 657 103160 99991 103288
rect 880 102880 99991 103160
rect 657 102616 99991 102880
rect 657 102336 99120 102616
rect 657 102072 99991 102336
rect 880 101792 99991 102072
rect 657 101528 99991 101792
rect 657 101248 99120 101528
rect 657 101120 99991 101248
rect 880 100840 99991 101120
rect 657 100576 99991 100840
rect 657 100296 99120 100576
rect 657 100032 99991 100296
rect 880 99752 99991 100032
rect 657 99624 99991 99752
rect 657 99344 99120 99624
rect 657 99080 99991 99344
rect 880 98800 99991 99080
rect 657 98536 99991 98800
rect 657 98256 99120 98536
rect 657 97992 99991 98256
rect 880 97712 99991 97992
rect 657 97584 99991 97712
rect 657 97304 99120 97584
rect 657 96904 99991 97304
rect 880 96632 99991 96904
rect 880 96624 99120 96632
rect 657 96352 99120 96624
rect 657 95952 99991 96352
rect 880 95680 99991 95952
rect 880 95672 99120 95680
rect 657 95400 99120 95672
rect 657 94864 99991 95400
rect 880 94592 99991 94864
rect 880 94584 99120 94592
rect 657 94312 99120 94584
rect 657 93776 99991 94312
rect 880 93640 99991 93776
rect 880 93496 99120 93640
rect 657 93360 99120 93496
rect 657 92824 99991 93360
rect 880 92688 99991 92824
rect 880 92544 99120 92688
rect 657 92408 99120 92544
rect 657 91736 99991 92408
rect 880 91600 99991 91736
rect 880 91456 99120 91600
rect 657 91320 99120 91456
rect 657 90784 99991 91320
rect 880 90648 99991 90784
rect 880 90504 99120 90648
rect 657 90368 99120 90504
rect 657 89696 99991 90368
rect 880 89416 99120 89696
rect 657 88744 99991 89416
rect 657 88608 99120 88744
rect 880 88464 99120 88608
rect 880 88328 99991 88464
rect 657 87656 99991 88328
rect 880 87376 99120 87656
rect 657 86704 99991 87376
rect 657 86568 99120 86704
rect 880 86424 99120 86568
rect 880 86288 99991 86424
rect 657 85752 99991 86288
rect 657 85480 99120 85752
rect 880 85472 99120 85480
rect 880 85200 99991 85472
rect 657 84664 99991 85200
rect 657 84528 99120 84664
rect 880 84384 99120 84528
rect 880 84248 99991 84384
rect 657 83712 99991 84248
rect 657 83440 99120 83712
rect 880 83432 99120 83440
rect 880 83160 99991 83432
rect 657 82760 99991 83160
rect 657 82488 99120 82760
rect 880 82480 99120 82488
rect 880 82208 99991 82480
rect 657 81808 99991 82208
rect 657 81528 99120 81808
rect 657 81400 99991 81528
rect 880 81120 99991 81400
rect 657 80720 99991 81120
rect 657 80440 99120 80720
rect 657 80312 99991 80440
rect 880 80032 99991 80312
rect 657 79768 99991 80032
rect 657 79488 99120 79768
rect 657 79360 99991 79488
rect 880 79080 99991 79360
rect 657 78816 99991 79080
rect 657 78536 99120 78816
rect 657 78272 99991 78536
rect 880 77992 99991 78272
rect 657 77864 99991 77992
rect 657 77584 99120 77864
rect 657 77320 99991 77584
rect 880 77040 99991 77320
rect 657 76776 99991 77040
rect 657 76496 99120 76776
rect 657 76232 99991 76496
rect 880 75952 99991 76232
rect 657 75824 99991 75952
rect 657 75544 99120 75824
rect 657 75144 99991 75544
rect 880 74872 99991 75144
rect 880 74864 99120 74872
rect 657 74592 99120 74864
rect 657 74192 99991 74592
rect 880 73912 99991 74192
rect 657 73784 99991 73912
rect 657 73504 99120 73784
rect 657 73104 99991 73504
rect 880 72832 99991 73104
rect 880 72824 99120 72832
rect 657 72552 99120 72824
rect 657 72016 99991 72552
rect 880 71880 99991 72016
rect 880 71736 99120 71880
rect 657 71600 99120 71736
rect 657 71064 99991 71600
rect 880 70928 99991 71064
rect 880 70784 99120 70928
rect 657 70648 99120 70784
rect 657 69976 99991 70648
rect 880 69840 99991 69976
rect 880 69696 99120 69840
rect 657 69560 99120 69696
rect 657 69024 99991 69560
rect 880 68888 99991 69024
rect 880 68744 99120 68888
rect 657 68608 99120 68744
rect 657 67936 99991 68608
rect 880 67656 99120 67936
rect 657 66848 99991 67656
rect 880 66568 99120 66848
rect 657 65896 99991 66568
rect 880 65616 99120 65896
rect 657 64944 99991 65616
rect 657 64808 99120 64944
rect 880 64664 99120 64808
rect 880 64528 99991 64664
rect 657 63992 99991 64528
rect 657 63720 99120 63992
rect 880 63712 99120 63720
rect 880 63440 99991 63712
rect 657 62904 99991 63440
rect 657 62768 99120 62904
rect 880 62624 99120 62768
rect 880 62488 99991 62624
rect 657 61952 99991 62488
rect 657 61680 99120 61952
rect 880 61672 99120 61680
rect 880 61400 99991 61672
rect 657 61000 99991 61400
rect 657 60728 99120 61000
rect 880 60720 99120 60728
rect 880 60448 99991 60720
rect 657 59912 99991 60448
rect 657 59640 99120 59912
rect 880 59632 99120 59640
rect 880 59360 99991 59632
rect 657 58960 99991 59360
rect 657 58680 99120 58960
rect 657 58552 99991 58680
rect 880 58272 99991 58552
rect 657 58008 99991 58272
rect 657 57728 99120 58008
rect 657 57600 99991 57728
rect 880 57320 99991 57600
rect 657 57056 99991 57320
rect 657 56776 99120 57056
rect 657 56512 99991 56776
rect 880 56232 99991 56512
rect 657 55968 99991 56232
rect 657 55688 99120 55968
rect 657 55424 99991 55688
rect 880 55144 99991 55424
rect 657 55016 99991 55144
rect 657 54736 99120 55016
rect 657 54472 99991 54736
rect 880 54192 99991 54472
rect 657 54064 99991 54192
rect 657 53784 99120 54064
rect 657 53384 99991 53784
rect 880 53104 99991 53384
rect 657 52976 99991 53104
rect 657 52696 99120 52976
rect 657 52432 99991 52696
rect 880 52152 99991 52432
rect 657 52024 99991 52152
rect 657 51744 99120 52024
rect 657 51344 99991 51744
rect 880 51072 99991 51344
rect 880 51064 99120 51072
rect 657 50792 99120 51064
rect 657 50256 99991 50792
rect 880 50120 99991 50256
rect 880 49976 99120 50120
rect 657 49840 99120 49976
rect 657 49304 99991 49840
rect 880 49032 99991 49304
rect 880 49024 99120 49032
rect 657 48752 99120 49024
rect 657 48216 99991 48752
rect 880 48080 99991 48216
rect 880 47936 99120 48080
rect 657 47800 99120 47936
rect 657 47128 99991 47800
rect 880 46848 99120 47128
rect 657 46176 99991 46848
rect 880 46040 99991 46176
rect 880 45896 99120 46040
rect 657 45760 99120 45896
rect 657 45088 99991 45760
rect 880 44808 99120 45088
rect 657 44136 99991 44808
rect 880 43856 99120 44136
rect 657 43184 99991 43856
rect 657 43048 99120 43184
rect 880 42904 99120 43048
rect 880 42768 99991 42904
rect 657 42096 99991 42768
rect 657 41960 99120 42096
rect 880 41816 99120 41960
rect 880 41680 99991 41816
rect 657 41144 99991 41680
rect 657 41008 99120 41144
rect 880 40864 99120 41008
rect 880 40728 99991 40864
rect 657 40192 99991 40728
rect 657 39920 99120 40192
rect 880 39912 99120 39920
rect 880 39640 99991 39912
rect 657 39240 99991 39640
rect 657 38968 99120 39240
rect 880 38960 99120 38968
rect 880 38688 99991 38960
rect 657 38152 99991 38688
rect 657 37880 99120 38152
rect 880 37872 99120 37880
rect 880 37600 99991 37872
rect 657 37200 99991 37600
rect 657 36920 99120 37200
rect 657 36792 99991 36920
rect 880 36512 99991 36792
rect 657 36248 99991 36512
rect 657 35968 99120 36248
rect 657 35840 99991 35968
rect 880 35560 99991 35840
rect 657 35160 99991 35560
rect 657 34880 99120 35160
rect 657 34752 99991 34880
rect 880 34472 99991 34752
rect 657 34208 99991 34472
rect 657 33928 99120 34208
rect 657 33664 99991 33928
rect 880 33384 99991 33664
rect 657 33256 99991 33384
rect 657 32976 99120 33256
rect 657 32712 99991 32976
rect 880 32432 99991 32712
rect 657 32304 99991 32432
rect 657 32024 99120 32304
rect 657 31624 99991 32024
rect 880 31344 99991 31624
rect 657 31216 99991 31344
rect 657 30936 99120 31216
rect 657 30672 99991 30936
rect 880 30392 99991 30672
rect 657 30264 99991 30392
rect 657 29984 99120 30264
rect 657 29584 99991 29984
rect 880 29312 99991 29584
rect 880 29304 99120 29312
rect 657 29032 99120 29304
rect 657 28496 99991 29032
rect 880 28224 99991 28496
rect 880 28216 99120 28224
rect 657 27944 99120 28216
rect 657 27544 99991 27944
rect 880 27272 99991 27544
rect 880 27264 99120 27272
rect 657 26992 99120 27264
rect 657 26456 99991 26992
rect 880 26320 99991 26456
rect 880 26176 99120 26320
rect 657 26040 99120 26176
rect 657 25368 99991 26040
rect 880 25088 99120 25368
rect 657 24416 99991 25088
rect 880 24280 99991 24416
rect 880 24136 99120 24280
rect 657 24000 99120 24136
rect 657 23328 99991 24000
rect 880 23048 99120 23328
rect 657 22376 99991 23048
rect 880 22096 99120 22376
rect 657 21288 99991 22096
rect 880 21008 99120 21288
rect 657 20336 99991 21008
rect 657 20200 99120 20336
rect 880 20056 99120 20200
rect 880 19920 99991 20056
rect 657 19384 99991 19920
rect 657 19248 99120 19384
rect 880 19104 99120 19248
rect 880 18968 99991 19104
rect 657 18432 99991 18968
rect 657 18160 99120 18432
rect 880 18152 99120 18160
rect 880 17880 99991 18152
rect 657 17344 99991 17880
rect 657 17072 99120 17344
rect 880 17064 99120 17072
rect 880 16792 99991 17064
rect 657 16392 99991 16792
rect 657 16120 99120 16392
rect 880 16112 99120 16120
rect 880 15840 99991 16112
rect 657 15440 99991 15840
rect 657 15160 99120 15440
rect 657 15032 99991 15160
rect 880 14752 99991 15032
rect 657 14352 99991 14752
rect 657 14080 99120 14352
rect 880 14072 99120 14080
rect 880 13800 99991 14072
rect 657 13400 99991 13800
rect 657 13120 99120 13400
rect 657 12992 99991 13120
rect 880 12712 99991 12992
rect 657 12448 99991 12712
rect 657 12168 99120 12448
rect 657 11904 99991 12168
rect 880 11624 99991 11904
rect 657 11496 99991 11624
rect 657 11216 99120 11496
rect 657 10952 99991 11216
rect 880 10672 99991 10952
rect 657 10408 99991 10672
rect 657 10128 99120 10408
rect 657 9864 99991 10128
rect 880 9584 99991 9864
rect 657 9456 99991 9584
rect 657 9176 99120 9456
rect 657 8776 99991 9176
rect 880 8504 99991 8776
rect 880 8496 99120 8504
rect 657 8224 99120 8496
rect 657 7824 99991 8224
rect 880 7544 99991 7824
rect 657 7416 99991 7544
rect 657 7136 99120 7416
rect 657 6736 99991 7136
rect 880 6464 99991 6736
rect 880 6456 99120 6464
rect 657 6184 99120 6456
rect 657 5784 99991 6184
rect 880 5512 99991 5784
rect 880 5504 99120 5512
rect 657 5232 99120 5504
rect 657 4696 99991 5232
rect 880 4560 99991 4696
rect 880 4416 99120 4560
rect 657 4280 99120 4416
rect 657 3608 99991 4280
rect 880 3472 99991 3608
rect 880 3328 99120 3472
rect 657 3192 99120 3328
rect 657 2656 99991 3192
rect 880 2520 99991 2656
rect 880 2376 99120 2520
rect 657 2240 99120 2376
rect 657 1568 99991 2240
rect 880 1288 99120 1568
rect 657 616 99991 1288
rect 880 443 99120 616
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
<< obsm4 >>
rect 1531 6835 4128 185061
rect 4608 6835 19488 185061
rect 19968 6835 34848 185061
rect 35328 6835 50208 185061
rect 50688 6835 65568 185061
rect 66048 6835 80928 185061
rect 81408 6835 96288 185061
rect 96768 6835 99853 185061
<< labels >>
rlabel metal3 s 0 12792 800 12912 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 124720 800 124840 6 addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 126760 800 126880 6 addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 130976 800 131096 6 addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 clk0
port 19 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 clk1
port 20 nsew signal output
rlabel metal2 s 1214 199200 1270 200000 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 3698 199200 3754 200000 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 6274 199200 6330 200000 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 8850 199200 8906 200000 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 11426 199200 11482 200000 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 14002 199200 14058 200000 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 16578 199200 16634 200000 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 19154 199200 19210 200000 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 99200 2320 100000 2440 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 99200 8304 100000 8424 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 99200 41896 100000 42016 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 99200 44888 100000 45008 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 99200 47880 100000 48000 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 99200 50872 100000 50992 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 99200 53864 100000 53984 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 99200 56856 100000 56976 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 99200 59712 100000 59832 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 99200 62704 100000 62824 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 99200 65696 100000 65816 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 99200 68688 100000 68808 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 99200 12248 100000 12368 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 99200 71680 100000 71800 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 99200 74672 100000 74792 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 99200 77664 100000 77784 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 99200 80520 100000 80640 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 99200 83512 100000 83632 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 99200 86504 100000 86624 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 99200 89496 100000 89616 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 99200 92488 100000 92608 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 99200 16192 100000 16312 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 99200 20136 100000 20256 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 99200 24080 100000 24200 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 99200 27072 100000 27192 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 99200 30064 100000 30184 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 99200 33056 100000 33176 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 99200 36048 100000 36168 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 99200 39040 100000 39160 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 99200 3272 100000 3392 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 99200 9256 100000 9376 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 99200 42984 100000 43104 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 99200 45840 100000 45960 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 99200 48832 100000 48952 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 99200 51824 100000 51944 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 99200 54816 100000 54936 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 99200 57808 100000 57928 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 99200 60800 100000 60920 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 99200 63792 100000 63912 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 99200 66648 100000 66768 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 99200 69640 100000 69760 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 99200 13200 100000 13320 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 99200 72632 100000 72752 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 99200 75624 100000 75744 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 99200 78616 100000 78736 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 99200 81608 100000 81728 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 99200 84464 100000 84584 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 99200 87456 100000 87576 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 99200 90448 100000 90568 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 99200 93440 100000 93560 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 99200 95480 100000 95600 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 99200 97384 100000 97504 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 99200 17144 100000 17264 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 99200 99424 100000 99544 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 99200 101328 100000 101448 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 99200 21088 100000 21208 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 99200 25168 100000 25288 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 99200 28024 100000 28144 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 99200 31016 100000 31136 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 99200 34008 100000 34128 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 99200 37000 100000 37120 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 99200 39992 100000 40112 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 99200 10208 100000 10328 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 99200 43936 100000 44056 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 99200 46928 100000 47048 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 99200 49920 100000 50040 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 99200 52776 100000 52896 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 99200 55768 100000 55888 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 99200 58760 100000 58880 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 99200 61752 100000 61872 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 99200 64744 100000 64864 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 99200 67736 100000 67856 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 99200 70728 100000 70848 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 99200 14152 100000 14272 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 99200 73584 100000 73704 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 99200 76576 100000 76696 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 99200 79568 100000 79688 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 99200 82560 100000 82680 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 99200 85552 100000 85672 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 99200 88544 100000 88664 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 99200 91400 100000 91520 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 99200 94392 100000 94512 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 99200 96432 100000 96552 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 99200 98336 100000 98456 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 99200 18232 100000 18352 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 99200 100376 100000 100496 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 99200 102416 100000 102536 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 99200 22176 100000 22296 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 99200 26120 100000 26240 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 99200 29112 100000 29232 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 99200 32104 100000 32224 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 99200 34960 100000 35080 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 99200 37952 100000 38072 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 99200 40944 100000 41064 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 99200 4360 100000 4480 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 99200 11296 100000 11416 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 99200 15240 100000 15360 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 99200 19184 100000 19304 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 99200 23128 100000 23248 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 99200 5312 100000 5432 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 99200 6264 100000 6384 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 99200 7216 100000 7336 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 csb1[1]
port 134 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 din0[0]
port 135 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 din0[10]
port 136 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 din0[11]
port 137 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 din0[12]
port 138 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 din0[13]
port 139 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 din0[14]
port 140 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 din0[15]
port 141 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 din0[16]
port 142 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 din0[17]
port 143 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 din0[18]
port 144 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 din0[19]
port 145 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 din0[1]
port 146 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 din0[20]
port 147 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 din0[21]
port 148 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 din0[22]
port 149 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 din0[23]
port 150 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 din0[24]
port 151 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 din0[25]
port 152 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 din0[26]
port 153 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 din0[27]
port 154 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 din0[28]
port 155 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 din0[29]
port 156 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 din0[2]
port 157 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 din0[30]
port 158 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 din0[31]
port 159 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 din0[3]
port 160 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 din0[4]
port 161 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 din0[5]
port 162 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 din0[6]
port 163 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 din0[7]
port 164 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 din0[8]
port 165 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 din0[9]
port 166 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 dout0[0]
port 167 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 dout0[10]
port 168 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 dout0[11]
port 169 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 dout0[12]
port 170 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 dout0[13]
port 171 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 dout0[15]
port 173 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 dout0[17]
port 175 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 dout0[18]
port 176 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 dout0[1]
port 178 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 dout0[20]
port 179 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 dout0[21]
port 180 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 dout0[22]
port 181 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 dout0[23]
port 182 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 dout0[24]
port 183 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 dout0[25]
port 184 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 dout0[26]
port 185 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 dout0[27]
port 186 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 dout0[29]
port 188 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 dout0[32]
port 192 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 dout0[33]
port 193 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 dout0[34]
port 194 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 dout0[35]
port 195 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 dout0[36]
port 196 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 dout0[37]
port 197 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 dout0[38]
port 198 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 dout0[39]
port 199 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 dout0[3]
port 200 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 dout0[40]
port 201 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 dout0[41]
port 202 nsew signal input
rlabel metal3 s 0 98880 800 99000 6 dout0[42]
port 203 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 dout0[43]
port 204 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 dout0[44]
port 205 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 dout0[45]
port 206 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 dout0[46]
port 207 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 dout0[47]
port 208 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 dout0[48]
port 209 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 dout0[49]
port 210 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 dout0[4]
port 211 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 dout0[50]
port 212 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 dout0[51]
port 213 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 dout0[52]
port 214 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 dout0[53]
port 215 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 dout0[54]
port 216 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 dout0[55]
port 217 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 dout0[56]
port 218 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 dout0[57]
port 219 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 dout0[58]
port 220 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 dout0[59]
port 221 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 dout0[5]
port 222 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 dout0[60]
port 223 nsew signal input
rlabel metal3 s 0 118464 800 118584 6 dout0[61]
port 224 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 dout0[62]
port 225 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 dout0[63]
port 226 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 dout0[6]
port 227 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 dout0[7]
port 228 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 dout0[8]
port 229 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 dout0[9]
port 230 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 dout1[0]
port 231 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 dout1[10]
port 232 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 dout1[11]
port 233 nsew signal input
rlabel metal3 s 0 146480 800 146600 6 dout1[12]
port 234 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 dout1[13]
port 235 nsew signal input
rlabel metal3 s 0 148520 800 148640 6 dout1[14]
port 236 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 dout1[15]
port 237 nsew signal input
rlabel metal3 s 0 150696 800 150816 6 dout1[16]
port 238 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 dout1[17]
port 239 nsew signal input
rlabel metal3 s 0 152736 800 152856 6 dout1[18]
port 240 nsew signal input
rlabel metal3 s 0 153824 800 153944 6 dout1[19]
port 241 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 dout1[1]
port 242 nsew signal input
rlabel metal3 s 0 154776 800 154896 6 dout1[20]
port 243 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 dout1[21]
port 244 nsew signal input
rlabel metal3 s 0 156816 800 156936 6 dout1[22]
port 245 nsew signal input
rlabel metal3 s 0 157904 800 158024 6 dout1[23]
port 246 nsew signal input
rlabel metal3 s 0 158992 800 159112 6 dout1[24]
port 247 nsew signal input
rlabel metal3 s 0 159944 800 160064 6 dout1[25]
port 248 nsew signal input
rlabel metal3 s 0 161032 800 161152 6 dout1[26]
port 249 nsew signal input
rlabel metal3 s 0 161984 800 162104 6 dout1[27]
port 250 nsew signal input
rlabel metal3 s 0 163072 800 163192 6 dout1[28]
port 251 nsew signal input
rlabel metal3 s 0 164160 800 164280 6 dout1[29]
port 252 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 dout1[2]
port 253 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 dout1[30]
port 254 nsew signal input
rlabel metal3 s 0 166200 800 166320 6 dout1[31]
port 255 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 dout1[32]
port 256 nsew signal input
rlabel metal3 s 0 168240 800 168360 6 dout1[33]
port 257 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 dout1[34]
port 258 nsew signal input
rlabel metal3 s 0 170280 800 170400 6 dout1[35]
port 259 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 dout1[36]
port 260 nsew signal input
rlabel metal3 s 0 172456 800 172576 6 dout1[37]
port 261 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 dout1[38]
port 262 nsew signal input
rlabel metal3 s 0 174496 800 174616 6 dout1[39]
port 263 nsew signal input
rlabel metal3 s 0 137232 800 137352 6 dout1[3]
port 264 nsew signal input
rlabel metal3 s 0 175584 800 175704 6 dout1[40]
port 265 nsew signal input
rlabel metal3 s 0 176536 800 176656 6 dout1[41]
port 266 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 dout1[42]
port 267 nsew signal input
rlabel metal3 s 0 178576 800 178696 6 dout1[43]
port 268 nsew signal input
rlabel metal3 s 0 179664 800 179784 6 dout1[44]
port 269 nsew signal input
rlabel metal3 s 0 180752 800 180872 6 dout1[45]
port 270 nsew signal input
rlabel metal3 s 0 181704 800 181824 6 dout1[46]
port 271 nsew signal input
rlabel metal3 s 0 182792 800 182912 6 dout1[47]
port 272 nsew signal input
rlabel metal3 s 0 183880 800 184000 6 dout1[48]
port 273 nsew signal input
rlabel metal3 s 0 184832 800 184952 6 dout1[49]
port 274 nsew signal input
rlabel metal3 s 0 138184 800 138304 6 dout1[4]
port 275 nsew signal input
rlabel metal3 s 0 185920 800 186040 6 dout1[50]
port 276 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 dout1[51]
port 277 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 dout1[52]
port 278 nsew signal input
rlabel metal3 s 0 189048 800 189168 6 dout1[53]
port 279 nsew signal input
rlabel metal3 s 0 190000 800 190120 6 dout1[54]
port 280 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 dout1[55]
port 281 nsew signal input
rlabel metal3 s 0 192176 800 192296 6 dout1[56]
port 282 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 dout1[57]
port 283 nsew signal input
rlabel metal3 s 0 194216 800 194336 6 dout1[58]
port 284 nsew signal input
rlabel metal3 s 0 195168 800 195288 6 dout1[59]
port 285 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 dout1[5]
port 286 nsew signal input
rlabel metal3 s 0 196256 800 196376 6 dout1[60]
port 287 nsew signal input
rlabel metal3 s 0 197344 800 197464 6 dout1[61]
port 288 nsew signal input
rlabel metal3 s 0 198296 800 198416 6 dout1[62]
port 289 nsew signal input
rlabel metal3 s 0 199384 800 199504 6 dout1[63]
port 290 nsew signal input
rlabel metal3 s 0 140224 800 140344 6 dout1[6]
port 291 nsew signal input
rlabel metal3 s 0 141312 800 141432 6 dout1[7]
port 292 nsew signal input
rlabel metal3 s 0 142400 800 142520 6 dout1[8]
port 293 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 dout1[9]
port 294 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 irq[0]
port 295 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 irq[10]
port 296 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 irq[11]
port 297 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 irq[12]
port 298 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 irq[13]
port 299 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 irq[14]
port 300 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 irq[15]
port 301 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 irq[1]
port 302 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 irq[2]
port 303 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 irq[3]
port 304 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 irq[4]
port 305 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 irq[5]
port 306 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 irq[6]
port 307 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 irq[7]
port 308 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 irq[8]
port 309 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 irq[9]
port 310 nsew signal input
rlabel metal3 s 0 416 800 536 6 jtag_tck
port 311 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 jtag_tdi
port 312 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 jtag_tdo
port 313 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 jtag_tms
port 314 nsew signal input
rlabel metal3 s 99200 103368 100000 103488 6 localMemory_wb_ack_o
port 315 nsew signal output
rlabel metal3 s 99200 109352 100000 109472 6 localMemory_wb_adr_i[0]
port 316 nsew signal input
rlabel metal3 s 99200 142944 100000 143064 6 localMemory_wb_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 99200 145936 100000 146056 6 localMemory_wb_adr_i[11]
port 318 nsew signal input
rlabel metal3 s 99200 148928 100000 149048 6 localMemory_wb_adr_i[12]
port 319 nsew signal input
rlabel metal3 s 99200 151920 100000 152040 6 localMemory_wb_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 99200 154912 100000 155032 6 localMemory_wb_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 99200 157768 100000 157888 6 localMemory_wb_adr_i[15]
port 322 nsew signal input
rlabel metal3 s 99200 160760 100000 160880 6 localMemory_wb_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 99200 163752 100000 163872 6 localMemory_wb_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 99200 166744 100000 166864 6 localMemory_wb_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 99200 169736 100000 169856 6 localMemory_wb_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 99200 113296 100000 113416 6 localMemory_wb_adr_i[1]
port 327 nsew signal input
rlabel metal3 s 99200 172728 100000 172848 6 localMemory_wb_adr_i[20]
port 328 nsew signal input
rlabel metal3 s 99200 175584 100000 175704 6 localMemory_wb_adr_i[21]
port 329 nsew signal input
rlabel metal3 s 99200 178576 100000 178696 6 localMemory_wb_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 99200 181568 100000 181688 6 localMemory_wb_adr_i[23]
port 331 nsew signal input
rlabel metal3 s 99200 117240 100000 117360 6 localMemory_wb_adr_i[2]
port 332 nsew signal input
rlabel metal3 s 99200 121184 100000 121304 6 localMemory_wb_adr_i[3]
port 333 nsew signal input
rlabel metal3 s 99200 125128 100000 125248 6 localMemory_wb_adr_i[4]
port 334 nsew signal input
rlabel metal3 s 99200 128120 100000 128240 6 localMemory_wb_adr_i[5]
port 335 nsew signal input
rlabel metal3 s 99200 131112 100000 131232 6 localMemory_wb_adr_i[6]
port 336 nsew signal input
rlabel metal3 s 99200 134104 100000 134224 6 localMemory_wb_adr_i[7]
port 337 nsew signal input
rlabel metal3 s 99200 136960 100000 137080 6 localMemory_wb_adr_i[8]
port 338 nsew signal input
rlabel metal3 s 99200 139952 100000 140072 6 localMemory_wb_adr_i[9]
port 339 nsew signal input
rlabel metal3 s 99200 104320 100000 104440 6 localMemory_wb_cyc_i
port 340 nsew signal input
rlabel metal3 s 99200 110304 100000 110424 6 localMemory_wb_data_i[0]
port 341 nsew signal input
rlabel metal3 s 99200 143896 100000 144016 6 localMemory_wb_data_i[10]
port 342 nsew signal input
rlabel metal3 s 99200 146888 100000 147008 6 localMemory_wb_data_i[11]
port 343 nsew signal input
rlabel metal3 s 99200 149880 100000 150000 6 localMemory_wb_data_i[12]
port 344 nsew signal input
rlabel metal3 s 99200 152872 100000 152992 6 localMemory_wb_data_i[13]
port 345 nsew signal input
rlabel metal3 s 99200 155864 100000 155984 6 localMemory_wb_data_i[14]
port 346 nsew signal input
rlabel metal3 s 99200 158856 100000 158976 6 localMemory_wb_data_i[15]
port 347 nsew signal input
rlabel metal3 s 99200 161712 100000 161832 6 localMemory_wb_data_i[16]
port 348 nsew signal input
rlabel metal3 s 99200 164704 100000 164824 6 localMemory_wb_data_i[17]
port 349 nsew signal input
rlabel metal3 s 99200 167696 100000 167816 6 localMemory_wb_data_i[18]
port 350 nsew signal input
rlabel metal3 s 99200 170688 100000 170808 6 localMemory_wb_data_i[19]
port 351 nsew signal input
rlabel metal3 s 99200 114248 100000 114368 6 localMemory_wb_data_i[1]
port 352 nsew signal input
rlabel metal3 s 99200 173680 100000 173800 6 localMemory_wb_data_i[20]
port 353 nsew signal input
rlabel metal3 s 99200 176672 100000 176792 6 localMemory_wb_data_i[21]
port 354 nsew signal input
rlabel metal3 s 99200 179664 100000 179784 6 localMemory_wb_data_i[22]
port 355 nsew signal input
rlabel metal3 s 99200 182520 100000 182640 6 localMemory_wb_data_i[23]
port 356 nsew signal input
rlabel metal3 s 99200 184560 100000 184680 6 localMemory_wb_data_i[24]
port 357 nsew signal input
rlabel metal3 s 99200 186600 100000 186720 6 localMemory_wb_data_i[25]
port 358 nsew signal input
rlabel metal3 s 99200 188504 100000 188624 6 localMemory_wb_data_i[26]
port 359 nsew signal input
rlabel metal3 s 99200 190544 100000 190664 6 localMemory_wb_data_i[27]
port 360 nsew signal input
rlabel metal3 s 99200 192448 100000 192568 6 localMemory_wb_data_i[28]
port 361 nsew signal input
rlabel metal3 s 99200 194488 100000 194608 6 localMemory_wb_data_i[29]
port 362 nsew signal input
rlabel metal3 s 99200 118192 100000 118312 6 localMemory_wb_data_i[2]
port 363 nsew signal input
rlabel metal3 s 99200 196392 100000 196512 6 localMemory_wb_data_i[30]
port 364 nsew signal input
rlabel metal3 s 99200 198432 100000 198552 6 localMemory_wb_data_i[31]
port 365 nsew signal input
rlabel metal3 s 99200 122136 100000 122256 6 localMemory_wb_data_i[3]
port 366 nsew signal input
rlabel metal3 s 99200 126080 100000 126200 6 localMemory_wb_data_i[4]
port 367 nsew signal input
rlabel metal3 s 99200 129072 100000 129192 6 localMemory_wb_data_i[5]
port 368 nsew signal input
rlabel metal3 s 99200 132064 100000 132184 6 localMemory_wb_data_i[6]
port 369 nsew signal input
rlabel metal3 s 99200 135056 100000 135176 6 localMemory_wb_data_i[7]
port 370 nsew signal input
rlabel metal3 s 99200 138048 100000 138168 6 localMemory_wb_data_i[8]
port 371 nsew signal input
rlabel metal3 s 99200 141040 100000 141160 6 localMemory_wb_data_i[9]
port 372 nsew signal input
rlabel metal3 s 99200 111256 100000 111376 6 localMemory_wb_data_o[0]
port 373 nsew signal output
rlabel metal3 s 99200 144984 100000 145104 6 localMemory_wb_data_o[10]
port 374 nsew signal output
rlabel metal3 s 99200 147976 100000 148096 6 localMemory_wb_data_o[11]
port 375 nsew signal output
rlabel metal3 s 99200 150832 100000 150952 6 localMemory_wb_data_o[12]
port 376 nsew signal output
rlabel metal3 s 99200 153824 100000 153944 6 localMemory_wb_data_o[13]
port 377 nsew signal output
rlabel metal3 s 99200 156816 100000 156936 6 localMemory_wb_data_o[14]
port 378 nsew signal output
rlabel metal3 s 99200 159808 100000 159928 6 localMemory_wb_data_o[15]
port 379 nsew signal output
rlabel metal3 s 99200 162800 100000 162920 6 localMemory_wb_data_o[16]
port 380 nsew signal output
rlabel metal3 s 99200 165792 100000 165912 6 localMemory_wb_data_o[17]
port 381 nsew signal output
rlabel metal3 s 99200 168648 100000 168768 6 localMemory_wb_data_o[18]
port 382 nsew signal output
rlabel metal3 s 99200 171640 100000 171760 6 localMemory_wb_data_o[19]
port 383 nsew signal output
rlabel metal3 s 99200 115200 100000 115320 6 localMemory_wb_data_o[1]
port 384 nsew signal output
rlabel metal3 s 99200 174632 100000 174752 6 localMemory_wb_data_o[20]
port 385 nsew signal output
rlabel metal3 s 99200 177624 100000 177744 6 localMemory_wb_data_o[21]
port 386 nsew signal output
rlabel metal3 s 99200 180616 100000 180736 6 localMemory_wb_data_o[22]
port 387 nsew signal output
rlabel metal3 s 99200 183608 100000 183728 6 localMemory_wb_data_o[23]
port 388 nsew signal output
rlabel metal3 s 99200 185512 100000 185632 6 localMemory_wb_data_o[24]
port 389 nsew signal output
rlabel metal3 s 99200 187552 100000 187672 6 localMemory_wb_data_o[25]
port 390 nsew signal output
rlabel metal3 s 99200 189456 100000 189576 6 localMemory_wb_data_o[26]
port 391 nsew signal output
rlabel metal3 s 99200 191496 100000 191616 6 localMemory_wb_data_o[27]
port 392 nsew signal output
rlabel metal3 s 99200 193536 100000 193656 6 localMemory_wb_data_o[28]
port 393 nsew signal output
rlabel metal3 s 99200 195440 100000 195560 6 localMemory_wb_data_o[29]
port 394 nsew signal output
rlabel metal3 s 99200 119144 100000 119264 6 localMemory_wb_data_o[2]
port 395 nsew signal output
rlabel metal3 s 99200 197480 100000 197600 6 localMemory_wb_data_o[30]
port 396 nsew signal output
rlabel metal3 s 99200 199384 100000 199504 6 localMemory_wb_data_o[31]
port 397 nsew signal output
rlabel metal3 s 99200 123088 100000 123208 6 localMemory_wb_data_o[3]
port 398 nsew signal output
rlabel metal3 s 99200 127168 100000 127288 6 localMemory_wb_data_o[4]
port 399 nsew signal output
rlabel metal3 s 99200 130024 100000 130144 6 localMemory_wb_data_o[5]
port 400 nsew signal output
rlabel metal3 s 99200 133016 100000 133136 6 localMemory_wb_data_o[6]
port 401 nsew signal output
rlabel metal3 s 99200 136008 100000 136128 6 localMemory_wb_data_o[7]
port 402 nsew signal output
rlabel metal3 s 99200 139000 100000 139120 6 localMemory_wb_data_o[8]
port 403 nsew signal output
rlabel metal3 s 99200 141992 100000 142112 6 localMemory_wb_data_o[9]
port 404 nsew signal output
rlabel metal3 s 99200 105272 100000 105392 6 localMemory_wb_error_o
port 405 nsew signal output
rlabel metal3 s 99200 112208 100000 112328 6 localMemory_wb_sel_i[0]
port 406 nsew signal input
rlabel metal3 s 99200 116288 100000 116408 6 localMemory_wb_sel_i[1]
port 407 nsew signal input
rlabel metal3 s 99200 120232 100000 120352 6 localMemory_wb_sel_i[2]
port 408 nsew signal input
rlabel metal3 s 99200 124176 100000 124296 6 localMemory_wb_sel_i[3]
port 409 nsew signal input
rlabel metal3 s 99200 106360 100000 106480 6 localMemory_wb_stall_o
port 410 nsew signal output
rlabel metal3 s 99200 107312 100000 107432 6 localMemory_wb_stb_i
port 411 nsew signal input
rlabel metal3 s 99200 108264 100000 108384 6 localMemory_wb_we_i
port 412 nsew signal input
rlabel metal2 s 21638 199200 21694 200000 6 manufacturerID[0]
port 413 nsew signal input
rlabel metal2 s 47306 199200 47362 200000 6 manufacturerID[10]
port 414 nsew signal input
rlabel metal2 s 24214 199200 24270 200000 6 manufacturerID[1]
port 415 nsew signal input
rlabel metal2 s 26790 199200 26846 200000 6 manufacturerID[2]
port 416 nsew signal input
rlabel metal2 s 29366 199200 29422 200000 6 manufacturerID[3]
port 417 nsew signal input
rlabel metal2 s 31942 199200 31998 200000 6 manufacturerID[4]
port 418 nsew signal input
rlabel metal2 s 34518 199200 34574 200000 6 manufacturerID[5]
port 419 nsew signal input
rlabel metal2 s 37094 199200 37150 200000 6 manufacturerID[6]
port 420 nsew signal input
rlabel metal2 s 39670 199200 39726 200000 6 manufacturerID[7]
port 421 nsew signal input
rlabel metal2 s 42154 199200 42210 200000 6 manufacturerID[8]
port 422 nsew signal input
rlabel metal2 s 44730 199200 44786 200000 6 manufacturerID[9]
port 423 nsew signal input
rlabel metal2 s 49882 199200 49938 200000 6 partID[0]
port 424 nsew signal input
rlabel metal2 s 75550 199200 75606 200000 6 partID[10]
port 425 nsew signal input
rlabel metal2 s 78126 199200 78182 200000 6 partID[11]
port 426 nsew signal input
rlabel metal2 s 80702 199200 80758 200000 6 partID[12]
port 427 nsew signal input
rlabel metal2 s 83186 199200 83242 200000 6 partID[13]
port 428 nsew signal input
rlabel metal2 s 85762 199200 85818 200000 6 partID[14]
port 429 nsew signal input
rlabel metal2 s 88338 199200 88394 200000 6 partID[15]
port 430 nsew signal input
rlabel metal2 s 52458 199200 52514 200000 6 partID[1]
port 431 nsew signal input
rlabel metal2 s 55034 199200 55090 200000 6 partID[2]
port 432 nsew signal input
rlabel metal2 s 57610 199200 57666 200000 6 partID[3]
port 433 nsew signal input
rlabel metal2 s 60186 199200 60242 200000 6 partID[4]
port 434 nsew signal input
rlabel metal2 s 62670 199200 62726 200000 6 partID[5]
port 435 nsew signal input
rlabel metal2 s 65246 199200 65302 200000 6 partID[6]
port 436 nsew signal input
rlabel metal2 s 67822 199200 67878 200000 6 partID[7]
port 437 nsew signal input
rlabel metal2 s 70398 199200 70454 200000 6 partID[8]
port 438 nsew signal input
rlabel metal2 s 72974 199200 73030 200000 6 partID[9]
port 439 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 probe_env[0]
port 440 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 probe_env[1]
port 441 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 probe_errorCode[0]
port 442 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 probe_errorCode[1]
port 443 nsew signal output
rlabel metal2 s 662 0 718 800 6 probe_isBranch
port 444 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 probe_isCompressed
port 445 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 probe_isLoad
port 446 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 probe_isStore
port 447 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 probe_jtagInstruction[0]
port 448 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 probe_jtagInstruction[1]
port 449 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 probe_jtagInstruction[2]
port 450 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 probe_jtagInstruction[3]
port 451 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 probe_jtagInstruction[4]
port 452 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 probe_opcode[0]
port 453 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 probe_opcode[1]
port 454 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 probe_opcode[2]
port 455 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 probe_opcode[3]
port 456 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 probe_opcode[4]
port 457 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 probe_opcode[5]
port 458 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 probe_opcode[6]
port 459 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 probe_programCounter[0]
port 460 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 probe_programCounter[10]
port 461 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 probe_programCounter[11]
port 462 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 probe_programCounter[12]
port 463 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 probe_programCounter[13]
port 464 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 probe_programCounter[14]
port 465 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 probe_programCounter[15]
port 466 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 probe_programCounter[16]
port 467 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 probe_programCounter[17]
port 468 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 probe_programCounter[18]
port 469 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 probe_programCounter[19]
port 470 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 probe_programCounter[1]
port 471 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 probe_programCounter[20]
port 472 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 probe_programCounter[21]
port 473 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 probe_programCounter[22]
port 474 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 probe_programCounter[23]
port 475 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 probe_programCounter[24]
port 476 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 probe_programCounter[25]
port 477 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 probe_programCounter[26]
port 478 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 probe_programCounter[27]
port 479 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 probe_programCounter[28]
port 480 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 probe_programCounter[29]
port 481 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 probe_programCounter[2]
port 482 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 probe_programCounter[30]
port 483 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 probe_programCounter[31]
port 484 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 probe_programCounter[3]
port 485 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 probe_programCounter[4]
port 486 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 probe_programCounter[5]
port 487 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 probe_programCounter[6]
port 488 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 probe_programCounter[7]
port 489 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 probe_programCounter[8]
port 490 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 probe_programCounter[9]
port 491 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 probe_state[0]
port 492 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 probe_state[1]
port 493 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 probe_takeBranch
port 494 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 495 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 495 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 495 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 495 nsew power input
rlabel metal2 s 90914 199200 90970 200000 6 versionID[0]
port 496 nsew signal input
rlabel metal2 s 93490 199200 93546 200000 6 versionID[1]
port 497 nsew signal input
rlabel metal2 s 96066 199200 96122 200000 6 versionID[2]
port 498 nsew signal input
rlabel metal2 s 98642 199200 98698 200000 6 versionID[3]
port 499 nsew signal input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 500 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 500 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 500 nsew ground input
rlabel metal3 s 99200 416 100000 536 6 wb_clk_i
port 501 nsew signal input
rlabel metal3 s 99200 1368 100000 1488 6 wb_rst_i
port 502 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 web0
port 503 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 wmask0[0]
port 504 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 wmask0[1]
port 505 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 wmask0[2]
port 506 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 wmask0[3]
port 507 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 47854972
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/finishing/ExperiarCore.magic.gds
string GDS_START 1598494
<< end >>

