magic
tech sky130A
magscale 1 2
timestamp 1683882473
<< viali >>
rect 41429 39593 41463 39627
rect 48881 39593 48915 39627
rect 1777 39457 1811 39491
rect 4261 39457 4295 39491
rect 19441 39457 19475 39491
rect 27353 39457 27387 39491
rect 56333 39457 56367 39491
rect 1593 39389 1627 39423
rect 2513 39389 2547 39423
rect 3985 39389 4019 39423
rect 27169 39389 27203 39423
rect 33885 39389 33919 39423
rect 56149 39389 56183 39423
rect 2789 39321 2823 39355
rect 33977 39253 34011 39287
rect 1593 38913 1627 38947
rect 2513 38913 2547 38947
rect 1777 38845 1811 38879
rect 2697 38845 2731 38879
rect 1593 38301 1627 38335
rect 1869 38233 1903 38267
rect 1593 37213 1627 37247
rect 1869 37145 1903 37179
rect 1593 36737 1627 36771
rect 1777 36669 1811 36703
rect 1593 35649 1627 35683
rect 1777 35581 1811 35615
rect 1593 35037 1627 35071
rect 1869 34969 1903 35003
rect 1869 34629 1903 34663
rect 1685 34561 1719 34595
rect 2421 34561 2455 34595
rect 2605 34493 2639 34527
rect 1685 33881 1719 33915
rect 1869 33881 1903 33915
rect 1593 33473 1627 33507
rect 1777 33405 1811 33439
rect 1685 32793 1719 32827
rect 1869 32793 1903 32827
rect 1593 32385 1627 32419
rect 1777 32317 1811 32351
rect 1869 31909 1903 31943
rect 1685 31773 1719 31807
rect 2421 31773 2455 31807
rect 2605 31773 2639 31807
rect 1593 31297 1627 31331
rect 1777 31229 1811 31263
rect 1685 30617 1719 30651
rect 1777 30549 1811 30583
rect 1593 30209 1627 30243
rect 2605 30209 2639 30243
rect 1777 30141 1811 30175
rect 2789 30073 2823 30107
rect 1685 29529 1719 29563
rect 2053 29529 2087 29563
rect 1593 29121 1627 29155
rect 2605 29121 2639 29155
rect 1777 29053 1811 29087
rect 2789 28985 2823 29019
rect 1685 28441 1719 28475
rect 1961 28373 1995 28407
rect 1593 28033 1627 28067
rect 2605 28033 2639 28067
rect 1777 27965 1811 27999
rect 2789 27897 2823 27931
rect 19809 27421 19843 27455
rect 19993 27421 20027 27455
rect 1685 27353 1719 27387
rect 1961 27285 1995 27319
rect 19901 27285 19935 27319
rect 19809 27081 19843 27115
rect 20637 27081 20671 27115
rect 2605 27013 2639 27047
rect 1593 26945 1627 26979
rect 14657 26945 14691 26979
rect 15393 26945 15427 26979
rect 15577 26945 15611 26979
rect 19533 26945 19567 26979
rect 20453 26945 20487 26979
rect 24317 26945 24351 26979
rect 34621 26945 34655 26979
rect 1777 26877 1811 26911
rect 14933 26877 14967 26911
rect 19625 26877 19659 26911
rect 19809 26877 19843 26911
rect 20269 26877 20303 26911
rect 24593 26877 24627 26911
rect 34897 26877 34931 26911
rect 2789 26809 2823 26843
rect 14841 26809 14875 26843
rect 14749 26741 14783 26775
rect 15393 26741 15427 26775
rect 24409 26741 24443 26775
rect 24501 26741 24535 26775
rect 34437 26741 34471 26775
rect 34805 26741 34839 26775
rect 1961 26537 1995 26571
rect 15761 26537 15795 26571
rect 15945 26537 15979 26571
rect 21373 26537 21407 26571
rect 22109 26537 22143 26571
rect 24593 26469 24627 26503
rect 33517 26469 33551 26503
rect 37749 26469 37783 26503
rect 2973 26401 3007 26435
rect 3157 26401 3191 26435
rect 6469 26401 6503 26435
rect 6561 26401 6595 26435
rect 8033 26401 8067 26435
rect 15117 26401 15151 26435
rect 20177 26401 20211 26435
rect 33609 26401 33643 26435
rect 34253 26401 34287 26435
rect 35357 26401 35391 26435
rect 35909 26401 35943 26435
rect 38485 26401 38519 26435
rect 38669 26401 38703 26435
rect 7941 26333 7975 26367
rect 13553 26333 13587 26367
rect 13737 26333 13771 26367
rect 14749 26333 14783 26367
rect 14933 26333 14967 26367
rect 20361 26333 20395 26367
rect 20453 26333 20487 26367
rect 20545 26333 20579 26367
rect 20637 26333 20671 26367
rect 22017 26333 22051 26367
rect 22293 26333 22327 26367
rect 24593 26333 24627 26367
rect 24869 26333 24903 26367
rect 31953 26333 31987 26367
rect 32321 26333 32355 26367
rect 34161 26333 34195 26367
rect 35081 26333 35115 26367
rect 35265 26333 35299 26367
rect 36277 26333 36311 26367
rect 37749 26333 37783 26367
rect 38025 26333 38059 26367
rect 38577 26333 38611 26367
rect 39037 26333 39071 26367
rect 39313 26333 39347 26367
rect 40049 26333 40083 26367
rect 40233 26333 40267 26367
rect 40325 26333 40359 26367
rect 40417 26333 40451 26367
rect 40601 26333 40635 26367
rect 1685 26265 1719 26299
rect 7849 26265 7883 26299
rect 13645 26265 13679 26299
rect 15577 26265 15611 26299
rect 15761 26265 15795 26299
rect 21189 26265 21223 26299
rect 21389 26265 21423 26299
rect 22201 26265 22235 26299
rect 24777 26265 24811 26299
rect 32689 26265 32723 26299
rect 33149 26265 33183 26299
rect 34897 26265 34931 26299
rect 36185 26265 36219 26299
rect 36394 26265 36428 26299
rect 40785 26265 40819 26299
rect 2513 26197 2547 26231
rect 2881 26197 2915 26231
rect 6009 26197 6043 26231
rect 6377 26197 6411 26231
rect 7481 26197 7515 26231
rect 21557 26197 21591 26231
rect 36553 26197 36587 26231
rect 37933 26197 37967 26231
rect 4261 25993 4295 26027
rect 8033 25993 8067 26027
rect 10701 25993 10735 26027
rect 15117 25993 15151 26027
rect 17969 25993 18003 26027
rect 35081 25993 35115 26027
rect 41429 25993 41463 26027
rect 42717 25993 42751 26027
rect 2605 25925 2639 25959
rect 17785 25925 17819 25959
rect 32689 25925 32723 25959
rect 38853 25925 38887 25959
rect 39865 25925 39899 25959
rect 1593 25857 1627 25891
rect 4169 25857 4203 25891
rect 7941 25857 7975 25891
rect 10609 25857 10643 25891
rect 14841 25857 14875 25891
rect 18061 25857 18095 25891
rect 18153 25857 18187 25891
rect 29837 25857 29871 25891
rect 29929 25857 29963 25891
rect 30113 25857 30147 25891
rect 30205 25857 30239 25891
rect 32321 25857 32355 25891
rect 32505 25857 32539 25891
rect 33609 25857 33643 25891
rect 33701 25857 33735 25891
rect 34989 25857 35023 25891
rect 35173 25857 35207 25891
rect 36001 25857 36035 25891
rect 36185 25857 36219 25891
rect 38761 25857 38795 25891
rect 38945 25857 38979 25891
rect 39221 25857 39255 25891
rect 40049 25857 40083 25891
rect 40141 25857 40175 25891
rect 41521 25857 41555 25891
rect 42625 25857 42659 25891
rect 1777 25789 1811 25823
rect 4353 25789 4387 25823
rect 10793 25789 10827 25823
rect 15117 25789 15151 25823
rect 41061 25789 41095 25823
rect 2789 25721 2823 25755
rect 33977 25721 34011 25755
rect 3801 25653 3835 25687
rect 10241 25653 10275 25687
rect 14933 25653 14967 25687
rect 18337 25653 18371 25687
rect 29653 25653 29687 25687
rect 33793 25653 33827 25687
rect 36093 25653 36127 25687
rect 40141 25653 40175 25687
rect 41245 25653 41279 25687
rect 6745 25449 6779 25483
rect 15669 25449 15703 25483
rect 22293 25449 22327 25483
rect 25973 25449 26007 25483
rect 36921 25449 36955 25483
rect 36553 25381 36587 25415
rect 10793 25313 10827 25347
rect 10885 25313 10919 25347
rect 29745 25313 29779 25347
rect 2053 25245 2087 25279
rect 2320 25245 2354 25279
rect 5365 25245 5399 25279
rect 7205 25245 7239 25279
rect 7472 25245 7506 25279
rect 14289 25245 14323 25279
rect 19441 25245 19475 25279
rect 19625 25245 19659 25279
rect 20913 25245 20947 25279
rect 21180 25245 21214 25279
rect 24593 25245 24627 25279
rect 24860 25245 24894 25279
rect 30021 25245 30055 25279
rect 37749 25245 37783 25279
rect 38025 25245 38059 25279
rect 5632 25177 5666 25211
rect 14556 25177 14590 25211
rect 36921 25177 36955 25211
rect 37565 25177 37599 25211
rect 3433 25109 3467 25143
rect 8585 25109 8619 25143
rect 10333 25109 10367 25143
rect 10701 25109 10735 25143
rect 19533 25109 19567 25143
rect 31125 25109 31159 25143
rect 37105 25109 37139 25143
rect 37933 25109 37967 25143
rect 4997 24905 5031 24939
rect 20177 24905 20211 24939
rect 29745 24905 29779 24939
rect 38485 24905 38519 24939
rect 38669 24905 38703 24939
rect 10048 24837 10082 24871
rect 32321 24837 32355 24871
rect 34621 24837 34655 24871
rect 1685 24769 1719 24803
rect 2605 24769 2639 24803
rect 3884 24769 3918 24803
rect 13369 24769 13403 24803
rect 13636 24769 13670 24803
rect 17121 24769 17155 24803
rect 19064 24769 19098 24803
rect 24225 24769 24259 24803
rect 24492 24769 24526 24803
rect 27353 24769 27387 24803
rect 29929 24769 29963 24803
rect 30205 24769 30239 24803
rect 30389 24769 30423 24803
rect 32505 24769 32539 24803
rect 32597 24769 32631 24803
rect 34253 24769 34287 24803
rect 34437 24769 34471 24803
rect 38301 24769 38335 24803
rect 38761 24769 38795 24803
rect 40868 24769 40902 24803
rect 3617 24701 3651 24735
rect 9781 24701 9815 24735
rect 16865 24701 16899 24735
rect 18797 24701 18831 24735
rect 27629 24701 27663 24735
rect 38393 24701 38427 24735
rect 40601 24701 40635 24735
rect 1961 24633 1995 24667
rect 2697 24565 2731 24599
rect 11161 24565 11195 24599
rect 14749 24565 14783 24599
rect 18245 24565 18279 24599
rect 25605 24565 25639 24599
rect 28917 24565 28951 24599
rect 32321 24565 32355 24599
rect 38117 24565 38151 24599
rect 41981 24565 42015 24599
rect 15945 24361 15979 24395
rect 16129 24361 16163 24395
rect 24777 24361 24811 24395
rect 27629 24361 27663 24395
rect 36277 24361 36311 24395
rect 38393 24361 38427 24395
rect 42349 24361 42383 24395
rect 19993 24293 20027 24327
rect 32321 24293 32355 24327
rect 21373 24225 21407 24259
rect 31953 24225 31987 24259
rect 2053 24157 2087 24191
rect 10241 24157 10275 24191
rect 10497 24157 10531 24191
rect 15577 24157 15611 24191
rect 19809 24157 19843 24191
rect 24961 24157 24995 24191
rect 25237 24157 25271 24191
rect 26249 24157 26283 24191
rect 32873 24157 32907 24191
rect 33140 24157 33174 24191
rect 34897 24157 34931 24191
rect 37013 24157 37047 24191
rect 37280 24157 37314 24191
rect 39129 24157 39163 24191
rect 39221 24157 39255 24191
rect 40969 24157 41003 24191
rect 41236 24157 41270 24191
rect 2320 24089 2354 24123
rect 15945 24089 15979 24123
rect 19441 24089 19475 24123
rect 21618 24089 21652 24123
rect 25145 24089 25179 24123
rect 26494 24089 26528 24123
rect 35142 24089 35176 24123
rect 38853 24089 38887 24123
rect 3433 24021 3467 24055
rect 11621 24021 11655 24055
rect 19625 24021 19659 24055
rect 19717 24021 19751 24055
rect 22753 24021 22787 24055
rect 32413 24021 32447 24055
rect 34253 24021 34287 24055
rect 39037 24021 39071 24055
rect 39405 24021 39439 24055
rect 1961 23817 1995 23851
rect 2513 23817 2547 23851
rect 2973 23817 3007 23851
rect 26157 23817 26191 23851
rect 31769 23817 31803 23851
rect 32505 23817 32539 23851
rect 41797 23817 41831 23851
rect 4905 23749 4939 23783
rect 16957 23749 16991 23783
rect 17157 23749 17191 23783
rect 20085 23749 20119 23783
rect 20545 23749 20579 23783
rect 28733 23749 28767 23783
rect 29377 23749 29411 23783
rect 40662 23749 40696 23783
rect 1685 23681 1719 23715
rect 2881 23681 2915 23715
rect 5181 23681 5215 23715
rect 6561 23681 6595 23715
rect 6817 23681 6851 23715
rect 20269 23681 20303 23715
rect 21005 23681 21039 23715
rect 26341 23681 26375 23715
rect 30205 23681 30239 23715
rect 31401 23681 31435 23715
rect 32321 23681 32355 23715
rect 32505 23681 32539 23715
rect 33057 23681 33091 23715
rect 3065 23613 3099 23647
rect 4997 23613 5031 23647
rect 20453 23613 20487 23647
rect 21097 23613 21131 23647
rect 26617 23613 26651 23647
rect 31493 23613 31527 23647
rect 33333 23613 33367 23647
rect 40417 23613 40451 23647
rect 17325 23545 17359 23579
rect 28365 23545 28399 23579
rect 28917 23545 28951 23579
rect 4997 23477 5031 23511
rect 5365 23477 5399 23511
rect 7941 23477 7975 23511
rect 17141 23477 17175 23511
rect 20361 23477 20395 23511
rect 26525 23477 26559 23511
rect 28733 23477 28767 23511
rect 31585 23477 31619 23511
rect 6285 23273 6319 23307
rect 7481 23273 7515 23307
rect 13553 23273 13587 23307
rect 16589 23273 16623 23307
rect 26065 23273 26099 23307
rect 26249 23273 26283 23307
rect 29745 23273 29779 23307
rect 32965 23273 32999 23307
rect 42165 23273 42199 23307
rect 17693 23205 17727 23239
rect 30113 23205 30147 23239
rect 1777 23137 1811 23171
rect 4997 23137 5031 23171
rect 6837 23137 6871 23171
rect 7665 23137 7699 23171
rect 28089 23137 28123 23171
rect 38577 23137 38611 23171
rect 1593 23069 1627 23103
rect 7481 23069 7515 23103
rect 7757 23069 7791 23103
rect 12173 23069 12207 23103
rect 16773 23069 16807 23103
rect 16865 23069 16899 23103
rect 16957 23069 16991 23103
rect 17049 23069 17083 23103
rect 17877 23069 17911 23103
rect 17969 23069 18003 23103
rect 21189 23069 21223 23103
rect 28365 23069 28399 23103
rect 28457 23069 28491 23103
rect 28549 23069 28583 23103
rect 28733 23069 28767 23103
rect 29929 23069 29963 23103
rect 30021 23069 30055 23103
rect 30205 23069 30239 23103
rect 32873 23069 32907 23103
rect 36461 23069 36495 23103
rect 36553 23069 36587 23103
rect 36645 23069 36679 23103
rect 36829 23069 36863 23103
rect 38761 23069 38795 23103
rect 40785 23069 40819 23103
rect 2605 23001 2639 23035
rect 4813 23001 4847 23035
rect 6745 23001 6779 23035
rect 12440 23001 12474 23035
rect 17693 23001 17727 23035
rect 25881 23001 25915 23035
rect 38945 23001 38979 23035
rect 41030 23001 41064 23035
rect 2697 22933 2731 22967
rect 4445 22933 4479 22967
rect 4905 22933 4939 22967
rect 6653 22933 6687 22967
rect 7941 22933 7975 22967
rect 21281 22933 21315 22967
rect 26081 22933 26115 22967
rect 36185 22933 36219 22967
rect 2421 22729 2455 22763
rect 5457 22729 5491 22763
rect 12817 22729 12851 22763
rect 13185 22729 13219 22763
rect 18797 22729 18831 22763
rect 23765 22729 23799 22763
rect 26157 22729 26191 22763
rect 29561 22729 29595 22763
rect 4344 22661 4378 22695
rect 29193 22661 29227 22695
rect 29393 22661 29427 22695
rect 31309 22661 31343 22695
rect 31493 22661 31527 22695
rect 2329 22593 2363 22627
rect 3249 22593 3283 22627
rect 4077 22593 4111 22627
rect 8033 22593 8067 22627
rect 8217 22593 8251 22627
rect 8309 22593 8343 22627
rect 9680 22593 9714 22627
rect 13001 22593 13035 22627
rect 13277 22593 13311 22627
rect 14933 22593 14967 22627
rect 15200 22593 15234 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 17325 22593 17359 22627
rect 18705 22593 18739 22627
rect 18889 22593 18923 22627
rect 22385 22593 22419 22627
rect 22652 22593 22686 22627
rect 24777 22593 24811 22627
rect 25044 22593 25078 22627
rect 2605 22525 2639 22559
rect 9413 22525 9447 22559
rect 8125 22457 8159 22491
rect 10793 22457 10827 22491
rect 16313 22457 16347 22491
rect 1961 22389 1995 22423
rect 3341 22389 3375 22423
rect 7849 22389 7883 22423
rect 17233 22389 17267 22423
rect 29377 22389 29411 22423
rect 31493 22389 31527 22423
rect 31677 22389 31711 22423
rect 3065 22185 3099 22219
rect 5181 22185 5215 22219
rect 9873 22185 9907 22219
rect 19809 22185 19843 22219
rect 23397 22185 23431 22219
rect 25145 22185 25179 22219
rect 30849 22185 30883 22219
rect 37933 22185 37967 22219
rect 19993 22117 20027 22151
rect 4997 22049 5031 22083
rect 18797 22049 18831 22083
rect 19901 22049 19935 22083
rect 35357 22049 35391 22083
rect 36553 22049 36587 22083
rect 36829 22049 36863 22083
rect 1685 21981 1719 22015
rect 1952 21981 1986 22015
rect 4261 21981 4295 22015
rect 5181 21981 5215 22015
rect 10057 21981 10091 22015
rect 10333 21981 10367 22015
rect 14473 21981 14507 22015
rect 14749 21981 14783 22015
rect 18705 21981 18739 22015
rect 19717 21981 19751 22015
rect 20177 21981 20211 22015
rect 21465 21981 21499 22015
rect 23581 21981 23615 22015
rect 23765 21981 23799 22015
rect 23857 21981 23891 22015
rect 25329 21981 25363 22015
rect 25605 21981 25639 22015
rect 29929 21981 29963 22015
rect 30205 21981 30239 22015
rect 32965 21981 32999 22015
rect 40233 21981 40267 22015
rect 4077 21913 4111 21947
rect 4905 21913 4939 21947
rect 21732 21913 21766 21947
rect 25513 21913 25547 21947
rect 30665 21913 30699 21947
rect 33232 21913 33266 21947
rect 34989 21913 35023 21947
rect 35173 21913 35207 21947
rect 40500 21913 40534 21947
rect 5365 21845 5399 21879
rect 10241 21845 10275 21879
rect 14289 21845 14323 21879
rect 14657 21845 14691 21879
rect 19441 21845 19475 21879
rect 22845 21845 22879 21879
rect 29745 21845 29779 21879
rect 30113 21845 30147 21879
rect 30865 21845 30899 21879
rect 31033 21845 31067 21879
rect 34345 21845 34379 21879
rect 41613 21845 41647 21879
rect 9505 21641 9539 21675
rect 33333 21641 33367 21675
rect 33701 21641 33735 21675
rect 37841 21641 37875 21675
rect 40601 21641 40635 21675
rect 40969 21641 41003 21675
rect 11897 21573 11931 21607
rect 13176 21573 13210 21607
rect 17417 21573 17451 21607
rect 17633 21573 17667 21607
rect 19441 21573 19475 21607
rect 22109 21573 22143 21607
rect 22477 21573 22511 21607
rect 28908 21573 28942 21607
rect 37473 21573 37507 21607
rect 37673 21573 37707 21607
rect 41705 21573 41739 21607
rect 1593 21505 1627 21539
rect 2513 21505 2547 21539
rect 5089 21505 5123 21539
rect 6561 21505 6595 21539
rect 7021 21505 7055 21539
rect 9321 21505 9355 21539
rect 9597 21505 9631 21539
rect 11989 21505 12023 21539
rect 12909 21505 12943 21539
rect 19349 21505 19383 21539
rect 21097 21505 21131 21539
rect 25973 21505 26007 21539
rect 30665 21505 30699 21539
rect 33517 21505 33551 21539
rect 33793 21505 33827 21539
rect 34253 21505 34287 21539
rect 34437 21505 34471 21539
rect 40785 21505 40819 21539
rect 41061 21505 41095 21539
rect 41521 21505 41555 21539
rect 1777 21437 1811 21471
rect 2697 21437 2731 21471
rect 5181 21437 5215 21471
rect 6929 21437 6963 21471
rect 26065 21437 26099 21471
rect 26157 21437 26191 21471
rect 26249 21437 26283 21471
rect 27353 21437 27387 21471
rect 27445 21437 27479 21471
rect 27537 21437 27571 21471
rect 27629 21437 27663 21471
rect 28641 21437 28675 21471
rect 30849 21437 30883 21471
rect 34345 21437 34379 21471
rect 14289 21369 14323 21403
rect 5181 21301 5215 21335
rect 5457 21301 5491 21335
rect 6653 21301 6687 21335
rect 7205 21301 7239 21335
rect 9137 21301 9171 21335
rect 11713 21301 11747 21335
rect 12173 21301 12207 21335
rect 17601 21301 17635 21335
rect 17785 21301 17819 21335
rect 21189 21301 21223 21335
rect 25789 21301 25823 21335
rect 27169 21301 27203 21335
rect 30021 21301 30055 21335
rect 37657 21301 37691 21335
rect 38117 21301 38151 21335
rect 41889 21301 41923 21335
rect 7757 21097 7791 21131
rect 11989 21097 12023 21131
rect 17969 21097 18003 21131
rect 18521 21097 18555 21131
rect 22201 21097 22235 21131
rect 23489 21097 23523 21131
rect 34345 21097 34379 21131
rect 44557 21097 44591 21131
rect 45201 21097 45235 21131
rect 30205 21029 30239 21063
rect 30573 21029 30607 21063
rect 31217 21029 31251 21063
rect 42349 21029 42383 21063
rect 2605 20961 2639 20995
rect 21741 20961 21775 20995
rect 23857 20961 23891 20995
rect 25973 20961 26007 20995
rect 27169 20961 27203 20995
rect 32965 20961 32999 20995
rect 40969 20961 41003 20995
rect 6377 20893 6411 20927
rect 9873 20893 9907 20927
rect 10609 20893 10643 20927
rect 17601 20893 17635 20927
rect 18429 20893 18463 20927
rect 18613 20893 18647 20927
rect 21005 20893 21039 20927
rect 21189 20893 21223 20927
rect 21281 20893 21315 20927
rect 22385 20893 22419 20927
rect 22569 20893 22603 20927
rect 22661 20893 22695 20927
rect 23673 20893 23707 20927
rect 23765 20893 23799 20927
rect 23949 20893 23983 20927
rect 26065 20893 26099 20927
rect 26157 20893 26191 20927
rect 26249 20893 26283 20927
rect 26985 20893 27019 20927
rect 27077 20893 27111 20927
rect 27261 20893 27295 20927
rect 30389 20893 30423 20927
rect 30665 20893 30699 20927
rect 31217 20893 31251 20927
rect 31401 20893 31435 20927
rect 33232 20893 33266 20927
rect 34897 20893 34931 20927
rect 36645 20893 36679 20927
rect 36912 20893 36946 20927
rect 38945 20893 38979 20927
rect 41236 20893 41270 20927
rect 44465 20893 44499 20927
rect 44649 20893 44683 20927
rect 45477 20893 45511 20927
rect 45569 20893 45603 20927
rect 45661 20893 45695 20927
rect 45845 20893 45879 20927
rect 2421 20825 2455 20859
rect 6644 20825 6678 20859
rect 9137 20825 9171 20859
rect 10876 20825 10910 20859
rect 15209 20825 15243 20859
rect 15945 20825 15979 20859
rect 17785 20825 17819 20859
rect 38577 20825 38611 20859
rect 38761 20825 38795 20859
rect 1961 20757 1995 20791
rect 2329 20757 2363 20791
rect 25789 20757 25823 20791
rect 26801 20757 26835 20791
rect 34989 20757 35023 20791
rect 38025 20757 38059 20791
rect 3341 20553 3375 20587
rect 6653 20553 6687 20587
rect 7021 20553 7055 20587
rect 9689 20553 9723 20587
rect 12357 20553 12391 20587
rect 14381 20553 14415 20587
rect 27169 20553 27203 20587
rect 30113 20553 30147 20587
rect 33701 20553 33735 20587
rect 2228 20485 2262 20519
rect 8576 20485 8610 20519
rect 12081 20485 12115 20519
rect 15200 20485 15234 20519
rect 34161 20485 34195 20519
rect 1961 20417 1995 20451
rect 3893 20417 3927 20451
rect 11713 20417 11747 20451
rect 11806 20417 11840 20451
rect 11989 20417 12023 20451
rect 12219 20417 12253 20451
rect 13001 20417 13035 20451
rect 13268 20417 13302 20451
rect 18245 20417 18279 20451
rect 19073 20417 19107 20451
rect 19340 20417 19374 20451
rect 25973 20417 26007 20451
rect 28989 20417 29023 20451
rect 30573 20417 30607 20451
rect 34069 20417 34103 20451
rect 34897 20417 34931 20451
rect 35081 20417 35115 20451
rect 37473 20417 37507 20451
rect 37740 20417 37774 20451
rect 40693 20417 40727 20451
rect 40960 20417 40994 20451
rect 7113 20349 7147 20383
rect 7297 20349 7331 20383
rect 8309 20349 8343 20383
rect 14933 20349 14967 20383
rect 18337 20349 18371 20383
rect 25789 20349 25823 20383
rect 26065 20349 26099 20383
rect 26157 20349 26191 20383
rect 26249 20349 26283 20383
rect 27353 20349 27387 20383
rect 27445 20349 27479 20383
rect 27537 20349 27571 20383
rect 27629 20349 27663 20383
rect 28733 20349 28767 20383
rect 30849 20349 30883 20383
rect 34253 20349 34287 20383
rect 16313 20281 16347 20315
rect 20453 20281 20487 20315
rect 3985 20213 4019 20247
rect 18613 20213 18647 20247
rect 34989 20213 35023 20247
rect 38853 20213 38887 20247
rect 42073 20213 42107 20247
rect 10517 20009 10551 20043
rect 13737 20009 13771 20043
rect 16865 20009 16899 20043
rect 19441 20009 19475 20043
rect 24593 20009 24627 20043
rect 25973 20009 26007 20043
rect 28733 20009 28767 20043
rect 37749 20009 37783 20043
rect 41429 20009 41463 20043
rect 5457 19941 5491 19975
rect 2789 19873 2823 19907
rect 5328 19873 5362 19907
rect 5549 19873 5583 19907
rect 6469 19873 6503 19907
rect 11253 19873 11287 19907
rect 16957 19873 16991 19907
rect 26433 19873 26467 19907
rect 30941 19873 30975 19907
rect 37105 19873 37139 19907
rect 38301 19873 38335 19907
rect 45201 19873 45235 19907
rect 1685 19805 1719 19839
rect 2513 19805 2547 19839
rect 5181 19805 5215 19839
rect 6377 19805 6411 19839
rect 6653 19805 6687 19839
rect 9873 19805 9907 19839
rect 10701 19805 10735 19839
rect 10793 19805 10827 19839
rect 13093 19805 13127 19839
rect 13186 19805 13220 19839
rect 13461 19805 13495 19839
rect 13558 19805 13592 19839
rect 15853 19805 15887 19839
rect 16681 19805 16715 19839
rect 19441 19805 19475 19839
rect 19625 19805 19659 19839
rect 20821 19805 20855 19839
rect 21373 19805 21407 19839
rect 23673 19805 23707 19839
rect 23949 19805 23983 19839
rect 24777 19805 24811 19839
rect 24869 19805 24903 19839
rect 24961 19805 24995 19839
rect 25053 19805 25087 19839
rect 26157 19805 26191 19839
rect 26249 19805 26283 19839
rect 26341 19805 26375 19839
rect 28917 19805 28951 19839
rect 29193 19805 29227 19839
rect 34161 19805 34195 19839
rect 37933 19805 37967 19839
rect 38025 19805 38059 19839
rect 38393 19805 38427 19839
rect 41429 19805 41463 19839
rect 41613 19805 41647 19839
rect 45477 19805 45511 19839
rect 45569 19805 45603 19839
rect 45661 19805 45695 19839
rect 45845 19805 45879 19839
rect 4077 19737 4111 19771
rect 4445 19737 4479 19771
rect 7113 19737 7147 19771
rect 9137 19737 9171 19771
rect 13369 19737 13403 19771
rect 15117 19737 15151 19771
rect 23857 19737 23891 19771
rect 30205 19737 30239 19771
rect 33977 19737 34011 19771
rect 36369 19737 36403 19771
rect 1961 19669 1995 19703
rect 5825 19669 5859 19703
rect 16497 19669 16531 19703
rect 20913 19669 20947 19703
rect 23489 19669 23523 19703
rect 29101 19669 29135 19703
rect 34345 19669 34379 19703
rect 2697 19465 2731 19499
rect 6009 19465 6043 19499
rect 7205 19465 7239 19499
rect 9873 19465 9907 19499
rect 16221 19465 16255 19499
rect 24409 19465 24443 19499
rect 26065 19465 26099 19499
rect 29377 19465 29411 19499
rect 32597 19465 32631 19499
rect 44925 19465 44959 19499
rect 2605 19397 2639 19431
rect 6929 19397 6963 19431
rect 15108 19397 15142 19431
rect 23296 19397 23330 19431
rect 37749 19397 37783 19431
rect 37841 19397 37875 19431
rect 3525 19329 3559 19363
rect 5641 19329 5675 19363
rect 6561 19329 6595 19363
rect 6654 19329 6688 19363
rect 6837 19329 6871 19363
rect 7067 19329 7101 19363
rect 8493 19329 8527 19363
rect 8760 19329 8794 19363
rect 14841 19329 14875 19363
rect 23029 19329 23063 19363
rect 29193 19329 29227 19363
rect 29377 19329 29411 19363
rect 29844 19329 29878 19363
rect 30104 19329 30138 19363
rect 32413 19329 32447 19363
rect 32597 19329 32631 19363
rect 33977 19329 34011 19363
rect 34161 19329 34195 19363
rect 34989 19329 35023 19363
rect 35265 19329 35299 19363
rect 36277 19329 36311 19363
rect 36645 19329 36679 19363
rect 37473 19329 37507 19363
rect 37621 19329 37655 19363
rect 37979 19329 38013 19363
rect 40969 19329 41003 19363
rect 41153 19329 41187 19363
rect 43085 19329 43119 19363
rect 43361 19329 43395 19363
rect 43913 19329 43947 19363
rect 44097 19329 44131 19363
rect 44741 19329 44775 19363
rect 44925 19329 44959 19363
rect 2789 19261 2823 19295
rect 3709 19261 3743 19295
rect 5733 19261 5767 19295
rect 26249 19261 26283 19295
rect 26341 19261 26375 19295
rect 26433 19261 26467 19295
rect 26525 19261 26559 19295
rect 27353 19261 27387 19295
rect 27445 19261 27479 19295
rect 27537 19261 27571 19295
rect 27629 19261 27663 19295
rect 34253 19261 34287 19295
rect 35173 19261 35207 19295
rect 35817 19261 35851 19295
rect 42901 19261 42935 19295
rect 43177 19261 43211 19295
rect 44005 19261 44039 19295
rect 27169 19193 27203 19227
rect 36553 19193 36587 19227
rect 38117 19193 38151 19227
rect 43269 19193 43303 19227
rect 2237 19125 2271 19159
rect 5641 19125 5675 19159
rect 31217 19125 31251 19159
rect 34805 19125 34839 19159
rect 40969 19125 41003 19159
rect 3249 18921 3283 18955
rect 6561 18921 6595 18955
rect 10149 18921 10183 18955
rect 11529 18921 11563 18955
rect 13369 18921 13403 18955
rect 22569 18921 22603 18955
rect 31401 18921 31435 18955
rect 44465 18921 44499 18955
rect 20637 18853 20671 18887
rect 26433 18853 26467 18887
rect 42441 18853 42475 18887
rect 42717 18853 42751 18887
rect 44649 18853 44683 18887
rect 12909 18785 12943 18819
rect 21189 18785 21223 18819
rect 22753 18785 22787 18819
rect 22937 18785 22971 18819
rect 26617 18785 26651 18819
rect 45201 18785 45235 18819
rect 45937 18785 45971 18819
rect 1869 18717 1903 18751
rect 2136 18717 2170 18751
rect 5181 18717 5215 18751
rect 5448 18717 5482 18751
rect 9505 18717 9539 18751
rect 9653 18717 9687 18751
rect 9970 18717 10004 18751
rect 11805 18717 11839 18751
rect 13185 18717 13219 18751
rect 19533 18717 19567 18751
rect 19809 18717 19843 18751
rect 20453 18717 20487 18751
rect 21373 18717 21407 18751
rect 21465 18717 21499 18751
rect 21557 18717 21591 18751
rect 21649 18717 21683 18751
rect 22845 18717 22879 18751
rect 23029 18717 23063 18751
rect 26709 18717 26743 18751
rect 26801 18717 26835 18751
rect 26893 18717 26927 18751
rect 31585 18717 31619 18751
rect 31677 18717 31711 18751
rect 36369 18717 36403 18751
rect 40233 18717 40267 18751
rect 40500 18717 40534 18751
rect 42625 18717 42659 18751
rect 42809 18717 42843 18751
rect 42901 18717 42935 18751
rect 45385 18717 45419 18751
rect 45477 18717 45511 18751
rect 9781 18649 9815 18683
rect 9873 18649 9907 18683
rect 11713 18649 11747 18683
rect 12265 18649 12299 18683
rect 13093 18649 13127 18683
rect 30021 18649 30055 18683
rect 30757 18649 30791 18683
rect 31953 18649 31987 18683
rect 32045 18649 32079 18683
rect 37105 18649 37139 18683
rect 44281 18649 44315 18683
rect 44497 18649 44531 18683
rect 45569 18649 45603 18683
rect 41613 18581 41647 18615
rect 19717 18377 19751 18411
rect 24409 18377 24443 18411
rect 40601 18377 40635 18411
rect 43913 18377 43947 18411
rect 44649 18377 44683 18411
rect 1869 18309 1903 18343
rect 2605 18309 2639 18343
rect 40325 18309 40359 18343
rect 43637 18309 43671 18343
rect 1593 18241 1627 18275
rect 17049 18241 17083 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 18604 18241 18638 18275
rect 22017 18241 22051 18275
rect 22273 18241 22307 18275
rect 24685 18241 24719 18275
rect 24869 18241 24903 18275
rect 25697 18241 25731 18275
rect 25789 18241 25823 18275
rect 30656 18241 30690 18275
rect 32413 18241 32447 18275
rect 32597 18241 32631 18275
rect 37473 18241 37507 18275
rect 37657 18241 37691 18275
rect 39957 18241 39991 18275
rect 40105 18241 40139 18275
rect 40233 18241 40267 18275
rect 40463 18241 40497 18275
rect 43269 18241 43303 18275
rect 43417 18241 43451 18275
rect 43545 18241 43579 18275
rect 43734 18241 43768 18275
rect 44465 18241 44499 18275
rect 44741 18241 44775 18275
rect 18337 18173 18371 18207
rect 24593 18173 24627 18207
rect 24777 18173 24811 18207
rect 25605 18173 25639 18207
rect 25881 18173 25915 18207
rect 30389 18173 30423 18207
rect 2789 18105 2823 18139
rect 25421 18105 25455 18139
rect 32413 18105 32447 18139
rect 44465 18105 44499 18139
rect 16865 18037 16899 18071
rect 23397 18037 23431 18071
rect 31769 18037 31803 18071
rect 37473 18037 37507 18071
rect 5365 17833 5399 17867
rect 17785 17833 17819 17867
rect 19441 17833 19475 17867
rect 21649 17833 21683 17867
rect 30665 17833 30699 17867
rect 35725 17833 35759 17867
rect 40693 17833 40727 17867
rect 8585 17765 8619 17799
rect 3985 17697 4019 17731
rect 16405 17697 16439 17731
rect 31217 17697 31251 17731
rect 36553 17697 36587 17731
rect 2513 17629 2547 17663
rect 7205 17629 7239 17663
rect 10793 17629 10827 17663
rect 14473 17629 14507 17663
rect 14657 17629 14691 17663
rect 14749 17629 14783 17663
rect 18245 17629 18279 17663
rect 19625 17629 19659 17663
rect 19901 17629 19935 17663
rect 21833 17629 21867 17663
rect 22017 17629 22051 17663
rect 22109 17629 22143 17663
rect 30849 17629 30883 17663
rect 30941 17629 30975 17663
rect 32873 17629 32907 17663
rect 34897 17629 34931 17663
rect 35633 17629 35667 17663
rect 35817 17629 35851 17663
rect 36820 17629 36854 17663
rect 40049 17629 40083 17663
rect 40197 17629 40231 17663
rect 40555 17629 40589 17663
rect 1685 17561 1719 17595
rect 2789 17561 2823 17595
rect 4252 17561 4286 17595
rect 7472 17561 7506 17595
rect 11060 17561 11094 17595
rect 16672 17561 16706 17595
rect 19809 17561 19843 17595
rect 31309 17561 31343 17595
rect 33140 17561 33174 17595
rect 40325 17561 40359 17595
rect 40417 17561 40451 17595
rect 1961 17493 1995 17527
rect 12173 17493 12207 17527
rect 14289 17493 14323 17527
rect 18429 17493 18463 17527
rect 34253 17493 34287 17527
rect 35081 17493 35115 17527
rect 37933 17493 37967 17527
rect 2329 17289 2363 17323
rect 4997 17289 5031 17323
rect 8953 17289 8987 17323
rect 11713 17289 11747 17323
rect 16957 17289 16991 17323
rect 19349 17289 19383 17323
rect 23581 17289 23615 17323
rect 33885 17289 33919 17323
rect 36737 17289 36771 17323
rect 37473 17289 37507 17323
rect 45753 17289 45787 17323
rect 45845 17289 45879 17323
rect 3249 17221 3283 17255
rect 8217 17221 8251 17255
rect 9321 17221 9355 17255
rect 12081 17221 12115 17255
rect 13268 17221 13302 17255
rect 34437 17221 34471 17255
rect 34529 17221 34563 17255
rect 44005 17221 44039 17255
rect 44097 17221 44131 17255
rect 4353 17153 4387 17187
rect 4501 17153 4535 17187
rect 4629 17153 4663 17187
rect 4721 17153 4755 17187
rect 4859 17153 4893 17187
rect 7849 17153 7883 17187
rect 9137 17153 9171 17187
rect 9413 17153 9447 17187
rect 11897 17153 11931 17187
rect 12173 17153 12207 17187
rect 15945 17153 15979 17187
rect 17325 17153 17359 17187
rect 17417 17153 17451 17187
rect 17969 17153 18003 17187
rect 18236 17153 18270 17187
rect 23765 17153 23799 17187
rect 23857 17153 23891 17187
rect 25053 17153 25087 17187
rect 27169 17153 27203 17187
rect 27436 17153 27470 17187
rect 29285 17153 29319 17187
rect 29469 17153 29503 17187
rect 32321 17153 32355 17187
rect 32873 17153 32907 17187
rect 34069 17153 34103 17187
rect 34161 17153 34195 17187
rect 34989 17153 35023 17187
rect 36093 17153 36127 17187
rect 36241 17153 36275 17187
rect 36369 17153 36403 17187
rect 36461 17153 36495 17187
rect 36599 17153 36633 17187
rect 37657 17153 37691 17187
rect 37933 17153 37967 17187
rect 43729 17153 43763 17187
rect 43822 17153 43856 17187
rect 44194 17153 44228 17187
rect 45661 17153 45695 17187
rect 46673 17153 46707 17187
rect 46857 17153 46891 17187
rect 46949 17153 46983 17187
rect 2421 17085 2455 17119
rect 2605 17085 2639 17119
rect 13001 17085 13035 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 23949 17085 23983 17119
rect 24041 17085 24075 17119
rect 24777 17085 24811 17119
rect 24869 17085 24903 17119
rect 24961 17085 24995 17119
rect 33333 17085 33367 17119
rect 35265 17085 35299 17119
rect 37749 17085 37783 17119
rect 14381 17017 14415 17051
rect 32597 17017 32631 17051
rect 37841 17017 37875 17051
rect 45477 17017 45511 17051
rect 46489 17017 46523 17051
rect 1961 16949 1995 16983
rect 3341 16949 3375 16983
rect 16221 16949 16255 16983
rect 24593 16949 24627 16983
rect 28549 16949 28583 16983
rect 29377 16949 29411 16983
rect 44373 16949 44407 16983
rect 46029 16949 46063 16983
rect 6285 16745 6319 16779
rect 9413 16745 9447 16779
rect 23305 16745 23339 16779
rect 27353 16745 27387 16779
rect 28917 16745 28951 16779
rect 36645 16745 36679 16779
rect 43545 16745 43579 16779
rect 4261 16677 4295 16711
rect 47961 16677 47995 16711
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 6745 16609 6779 16643
rect 10149 16609 10183 16643
rect 14841 16609 14875 16643
rect 16681 16609 16715 16643
rect 16865 16609 16899 16643
rect 18429 16609 18463 16643
rect 23489 16609 23523 16643
rect 23581 16609 23615 16643
rect 25329 16609 25363 16643
rect 27537 16609 27571 16643
rect 29101 16609 29135 16643
rect 29745 16609 29779 16643
rect 37289 16609 37323 16643
rect 38025 16609 38059 16643
rect 40325 16609 40359 16643
rect 42165 16609 42199 16643
rect 46305 16609 46339 16643
rect 47501 16609 47535 16643
rect 3433 16541 3467 16575
rect 5641 16541 5675 16575
rect 5789 16541 5823 16575
rect 5917 16541 5951 16575
rect 6009 16541 6043 16575
rect 6147 16541 6181 16575
rect 7012 16541 7046 16575
rect 9689 16541 9723 16575
rect 15025 16541 15059 16575
rect 15301 16541 15335 16575
rect 16590 16541 16624 16575
rect 16773 16541 16807 16575
rect 18061 16541 18095 16575
rect 23673 16541 23707 16575
rect 23765 16541 23799 16575
rect 25053 16541 25087 16575
rect 25145 16541 25179 16575
rect 25237 16541 25271 16575
rect 27629 16541 27663 16575
rect 27905 16541 27939 16575
rect 28825 16541 28859 16575
rect 34897 16541 34931 16575
rect 35081 16541 35115 16575
rect 36645 16541 36679 16575
rect 36829 16541 36863 16575
rect 45937 16541 45971 16575
rect 46121 16541 46155 16575
rect 46397 16541 46431 16575
rect 47593 16541 47627 16575
rect 4077 16473 4111 16507
rect 9597 16473 9631 16507
rect 17877 16473 17911 16507
rect 27997 16473 28031 16507
rect 29101 16473 29135 16507
rect 29990 16473 30024 16507
rect 37565 16473 37599 16507
rect 37657 16473 37691 16507
rect 40570 16473 40604 16507
rect 42432 16473 42466 16507
rect 8125 16405 8159 16439
rect 15209 16405 15243 16439
rect 16405 16405 16439 16439
rect 24869 16405 24903 16439
rect 31125 16405 31159 16439
rect 34989 16405 35023 16439
rect 37473 16405 37507 16439
rect 41705 16405 41739 16439
rect 3433 16201 3467 16235
rect 14381 16201 14415 16235
rect 16313 16201 16347 16235
rect 18153 16201 18187 16235
rect 18521 16201 18555 16235
rect 34529 16201 34563 16235
rect 37841 16201 37875 16235
rect 40049 16201 40083 16235
rect 40417 16201 40451 16235
rect 45569 16201 45603 16235
rect 1869 16133 1903 16167
rect 15200 16133 15234 16167
rect 17049 16133 17083 16167
rect 26065 16133 26099 16167
rect 29837 16133 29871 16167
rect 36645 16133 36679 16167
rect 37473 16133 37507 16167
rect 37673 16133 37707 16167
rect 1593 16065 1627 16099
rect 3341 16065 3375 16099
rect 6561 16065 6595 16099
rect 7665 16065 7699 16099
rect 7921 16065 7955 16099
rect 13268 16065 13302 16099
rect 14933 16065 14967 16099
rect 16957 16065 16991 16099
rect 18337 16065 18371 16099
rect 18613 16065 18647 16099
rect 19625 16065 19659 16099
rect 20637 16065 20671 16099
rect 20729 16065 20763 16099
rect 20913 16065 20947 16099
rect 22273 16065 22307 16099
rect 24501 16065 24535 16099
rect 24685 16065 24719 16099
rect 25881 16065 25915 16099
rect 26157 16065 26191 16099
rect 29469 16065 29503 16099
rect 30573 16065 30607 16099
rect 30757 16065 30791 16099
rect 33885 16065 33919 16099
rect 33978 16065 34012 16099
rect 34161 16065 34195 16099
rect 34253 16065 34287 16099
rect 34391 16065 34425 16099
rect 36829 16065 36863 16099
rect 36921 16065 36955 16099
rect 40233 16065 40267 16099
rect 40509 16065 40543 16099
rect 43545 16065 43579 16099
rect 43638 16065 43672 16099
rect 43821 16065 43855 16099
rect 43913 16065 43947 16099
rect 44010 16065 44044 16099
rect 46029 16065 46063 16099
rect 3617 15997 3651 16031
rect 6745 15997 6779 16031
rect 13001 15997 13035 16031
rect 19441 15997 19475 16031
rect 19717 15997 19751 16031
rect 19809 15997 19843 16031
rect 19901 15997 19935 16031
rect 20453 15997 20487 16031
rect 20821 15997 20855 16031
rect 22017 15997 22051 16031
rect 26617 15997 26651 16031
rect 45753 15997 45787 16031
rect 45845 15997 45879 16031
rect 45937 15997 45971 16031
rect 44189 15929 44223 15963
rect 2973 15861 3007 15895
rect 9045 15861 9079 15895
rect 23397 15861 23431 15895
rect 24593 15861 24627 15895
rect 30573 15861 30607 15895
rect 36645 15861 36679 15895
rect 37657 15861 37691 15895
rect 7389 15657 7423 15691
rect 14933 15657 14967 15691
rect 22109 15657 22143 15691
rect 29745 15657 29779 15691
rect 33885 15657 33919 15691
rect 27445 15589 27479 15623
rect 36829 15589 36863 15623
rect 36921 15589 36955 15623
rect 7849 15521 7883 15555
rect 8033 15521 8067 15555
rect 17509 15521 17543 15555
rect 20177 15521 20211 15555
rect 21281 15521 21315 15555
rect 22661 15521 22695 15555
rect 41153 15521 41187 15555
rect 1593 15453 1627 15487
rect 14289 15453 14323 15487
rect 14437 15453 14471 15487
rect 14657 15453 14691 15487
rect 14754 15453 14788 15487
rect 19993 15453 20027 15487
rect 21005 15453 21039 15487
rect 22293 15453 22327 15487
rect 22385 15453 22419 15487
rect 24593 15453 24627 15487
rect 27721 15453 27755 15487
rect 29929 15453 29963 15487
rect 30021 15453 30055 15487
rect 30205 15453 30239 15487
rect 30297 15453 30331 15487
rect 33241 15453 33275 15487
rect 33334 15453 33368 15487
rect 33706 15453 33740 15487
rect 36737 15453 36771 15487
rect 37013 15453 37047 15487
rect 1869 15385 1903 15419
rect 2605 15385 2639 15419
rect 2789 15385 2823 15419
rect 14565 15385 14599 15419
rect 17776 15385 17810 15419
rect 22753 15385 22787 15419
rect 24869 15385 24903 15419
rect 27445 15385 27479 15419
rect 33517 15385 33551 15419
rect 33609 15385 33643 15419
rect 41420 15385 41454 15419
rect 7757 15317 7791 15351
rect 18889 15317 18923 15351
rect 27629 15317 27663 15351
rect 36553 15317 36587 15351
rect 42533 15317 42567 15351
rect 11069 15113 11103 15147
rect 19533 15113 19567 15147
rect 26617 15113 26651 15147
rect 27813 15113 27847 15147
rect 38853 15113 38887 15147
rect 42625 15113 42659 15147
rect 42993 15113 43027 15147
rect 1685 15045 1719 15079
rect 2964 15045 2998 15079
rect 19901 15045 19935 15079
rect 28089 15045 28123 15079
rect 31033 15045 31067 15079
rect 31401 15045 31435 15079
rect 32566 15045 32600 15079
rect 36535 15045 36569 15079
rect 44005 15045 44039 15079
rect 1869 14977 1903 15011
rect 7104 14977 7138 15011
rect 9689 14977 9723 15011
rect 9956 14977 9990 15011
rect 19717 14977 19751 15011
rect 19993 14977 20027 15011
rect 23213 14977 23247 15011
rect 23949 14977 23983 15011
rect 24216 14977 24250 15011
rect 25973 14977 26007 15011
rect 26121 14977 26155 15011
rect 26249 14977 26283 15011
rect 26341 14977 26375 15011
rect 26438 14977 26472 15011
rect 27813 14977 27847 15011
rect 27905 14977 27939 15011
rect 31217 14977 31251 15011
rect 32321 14977 32355 15011
rect 35817 14977 35851 15011
rect 36001 14977 36035 15011
rect 37473 14977 37507 15011
rect 37729 14977 37763 15011
rect 42809 14977 42843 15011
rect 43085 14977 43119 15011
rect 43729 14977 43763 15011
rect 43822 14977 43856 15011
rect 44097 14977 44131 15011
rect 44194 14977 44228 15011
rect 45109 14977 45143 15011
rect 2697 14909 2731 14943
rect 6837 14909 6871 14943
rect 22845 14909 22879 14943
rect 23029 14909 23063 14943
rect 23121 14909 23155 14943
rect 23305 14909 23339 14943
rect 36829 14909 36863 14943
rect 45201 14909 45235 14943
rect 25329 14841 25363 14875
rect 35817 14841 35851 14875
rect 44373 14841 44407 14875
rect 45477 14841 45511 14875
rect 4077 14773 4111 14807
rect 8217 14773 8251 14807
rect 33701 14773 33735 14807
rect 7021 14569 7055 14603
rect 11805 14569 11839 14603
rect 36645 14569 36679 14603
rect 12725 14501 12759 14535
rect 17601 14501 17635 14535
rect 18245 14501 18279 14535
rect 24685 14501 24719 14535
rect 24777 14501 24811 14535
rect 26709 14501 26743 14535
rect 26801 14501 26835 14535
rect 40141 14501 40175 14535
rect 3985 14433 4019 14467
rect 7665 14433 7699 14467
rect 13461 14433 13495 14467
rect 24869 14433 24903 14467
rect 25697 14433 25731 14467
rect 26893 14433 26927 14467
rect 28273 14433 28307 14467
rect 31217 14433 31251 14467
rect 1593 14365 1627 14399
rect 2605 14365 2639 14399
rect 4261 14365 4295 14399
rect 7481 14365 7515 14399
rect 11161 14365 11195 14399
rect 11309 14365 11343 14399
rect 11529 14365 11563 14399
rect 11667 14365 11701 14399
rect 13001 14365 13035 14399
rect 16221 14365 16255 14399
rect 18061 14365 18095 14399
rect 24593 14365 24627 14399
rect 25881 14365 25915 14399
rect 26157 14365 26191 14399
rect 26617 14365 26651 14399
rect 30941 14365 30975 14399
rect 36553 14365 36587 14399
rect 36737 14365 36771 14399
rect 40417 14365 40451 14399
rect 41153 14365 41187 14399
rect 41337 14365 41371 14399
rect 1869 14297 1903 14331
rect 2789 14297 2823 14331
rect 5641 14297 5675 14331
rect 11437 14297 11471 14331
rect 12909 14297 12943 14331
rect 16488 14297 16522 14331
rect 22017 14297 22051 14331
rect 27537 14297 27571 14331
rect 27813 14297 27847 14331
rect 27905 14297 27939 14331
rect 31033 14297 31067 14331
rect 40141 14297 40175 14331
rect 7389 14229 7423 14263
rect 23305 14229 23339 14263
rect 26065 14229 26099 14263
rect 27721 14229 27755 14263
rect 30573 14229 30607 14263
rect 40325 14229 40359 14263
rect 41245 14229 41279 14263
rect 4077 14025 4111 14059
rect 4445 14025 4479 14059
rect 15117 14025 15151 14059
rect 17049 14025 17083 14059
rect 17417 14025 17451 14059
rect 20913 14025 20947 14059
rect 23673 14025 23707 14059
rect 30757 14025 30791 14059
rect 33793 14025 33827 14059
rect 38025 14025 38059 14059
rect 41061 14025 41095 14059
rect 33425 13957 33459 13991
rect 37749 13957 37783 13991
rect 1685 13889 1719 13923
rect 1952 13889 1986 13923
rect 4537 13889 4571 13923
rect 8300 13889 8334 13923
rect 11989 13889 12023 13923
rect 12173 13889 12207 13923
rect 12725 13889 12759 13923
rect 13737 13889 13771 13923
rect 14004 13889 14038 13923
rect 17233 13889 17267 13923
rect 17509 13889 17543 13923
rect 21189 13889 21223 13923
rect 21281 13889 21315 13923
rect 22017 13889 22051 13923
rect 23857 13889 23891 13923
rect 23949 13889 23983 13923
rect 24041 13889 24075 13923
rect 29377 13889 29411 13923
rect 29644 13889 29678 13923
rect 33149 13889 33183 13923
rect 33297 13889 33331 13923
rect 33517 13889 33551 13923
rect 33614 13889 33648 13923
rect 37473 13889 37507 13923
rect 37657 13889 37691 13923
rect 37841 13889 37875 13923
rect 38853 13889 38887 13923
rect 39681 13889 39715 13923
rect 39937 13889 39971 13923
rect 4721 13821 4755 13855
rect 8033 13821 8067 13855
rect 11713 13821 11747 13855
rect 11897 13821 11931 13855
rect 12081 13821 12115 13855
rect 12909 13821 12943 13855
rect 21097 13821 21131 13855
rect 21373 13821 21407 13855
rect 22201 13821 22235 13855
rect 24133 13821 24167 13855
rect 38669 13821 38703 13855
rect 39037 13821 39071 13855
rect 3065 13685 3099 13719
rect 9413 13685 9447 13719
rect 1961 13481 1995 13515
rect 9137 13481 9171 13515
rect 11989 13481 12023 13515
rect 14473 13481 14507 13515
rect 16773 13481 16807 13515
rect 21649 13481 21683 13515
rect 27537 13481 27571 13515
rect 29929 13481 29963 13515
rect 30297 13481 30331 13515
rect 2605 13345 2639 13379
rect 9689 13345 9723 13379
rect 12265 13345 12299 13379
rect 12449 13345 12483 13379
rect 16405 13345 16439 13379
rect 21833 13345 21867 13379
rect 22017 13345 22051 13379
rect 30389 13345 30423 13379
rect 30941 13345 30975 13379
rect 37381 13345 37415 13379
rect 2421 13277 2455 13311
rect 4261 13277 4295 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 6009 13277 6043 13311
rect 12173 13277 12207 13311
rect 12357 13277 12391 13311
rect 14657 13277 14691 13311
rect 14841 13277 14875 13311
rect 14933 13277 14967 13311
rect 16589 13277 16623 13311
rect 17509 13277 17543 13311
rect 21925 13277 21959 13311
rect 22109 13277 22143 13311
rect 22661 13277 22695 13311
rect 22937 13277 22971 13311
rect 27261 13277 27295 13311
rect 27353 13277 27387 13311
rect 30113 13277 30147 13311
rect 30849 13277 30883 13311
rect 31677 13277 31711 13311
rect 32045 13277 32079 13311
rect 35725 13277 35759 13311
rect 36001 13277 36035 13311
rect 36093 13277 36127 13311
rect 37105 13277 37139 13311
rect 41521 13277 41555 13311
rect 41777 13277 41811 13311
rect 3249 13209 3283 13243
rect 4077 13209 4111 13243
rect 5457 13209 5491 13243
rect 6254 13209 6288 13243
rect 17776 13209 17810 13243
rect 31861 13209 31895 13243
rect 31953 13209 31987 13243
rect 35909 13209 35943 13243
rect 2329 13141 2363 13175
rect 3341 13141 3375 13175
rect 7389 13141 7423 13175
rect 9505 13141 9539 13175
rect 9597 13141 9631 13175
rect 18889 13141 18923 13175
rect 32229 13141 32263 13175
rect 36277 13141 36311 13175
rect 42901 13141 42935 13175
rect 13093 12937 13127 12971
rect 18521 12937 18555 12971
rect 24869 12937 24903 12971
rect 27629 12937 27663 12971
rect 32781 12937 32815 12971
rect 37473 12937 37507 12971
rect 37841 12937 37875 12971
rect 2605 12869 2639 12903
rect 2789 12869 2823 12903
rect 18889 12869 18923 12903
rect 26341 12869 26375 12903
rect 1593 12801 1627 12835
rect 9045 12801 9079 12835
rect 9505 12801 9539 12835
rect 11713 12801 11747 12835
rect 11980 12801 12014 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 18705 12801 18739 12835
rect 18981 12801 19015 12835
rect 22201 12801 22235 12835
rect 22293 12801 22327 12835
rect 23756 12801 23790 12835
rect 25973 12801 26007 12835
rect 27169 12801 27203 12835
rect 27997 12801 28031 12835
rect 28273 12801 28307 12835
rect 28917 12801 28951 12835
rect 31585 12801 31619 12835
rect 33149 12801 33183 12835
rect 33241 12801 33275 12835
rect 35624 12801 35658 12835
rect 37933 12801 37967 12835
rect 40693 12801 40727 12835
rect 40877 12801 40911 12835
rect 1777 12733 1811 12767
rect 9137 12733 9171 12767
rect 22569 12733 22603 12767
rect 22661 12733 22695 12767
rect 23489 12733 23523 12767
rect 29193 12733 29227 12767
rect 31401 12733 31435 12767
rect 33425 12733 33459 12767
rect 35357 12733 35391 12767
rect 38025 12733 38059 12767
rect 8769 12597 8803 12631
rect 9229 12597 9263 12631
rect 9321 12597 9355 12631
rect 16865 12597 16899 12631
rect 22017 12597 22051 12631
rect 27261 12597 27295 12631
rect 31769 12597 31803 12631
rect 36737 12597 36771 12631
rect 40693 12597 40727 12631
rect 11897 12393 11931 12427
rect 17417 12393 17451 12427
rect 22477 12393 22511 12427
rect 24593 12393 24627 12427
rect 27905 12393 27939 12427
rect 29009 12393 29043 12427
rect 35817 12393 35851 12427
rect 36553 12393 36587 12427
rect 10609 12325 10643 12359
rect 25789 12325 25823 12359
rect 39221 12325 39255 12359
rect 16313 12257 16347 12291
rect 21097 12257 21131 12291
rect 27537 12257 27571 12291
rect 37013 12257 37047 12291
rect 37197 12257 37231 12291
rect 1685 12189 1719 12223
rect 3985 12189 4019 12223
rect 7205 12189 7239 12223
rect 7573 12189 7607 12223
rect 7849 12189 7883 12223
rect 8493 12189 8527 12223
rect 12081 12189 12115 12223
rect 12357 12189 12391 12223
rect 14381 12189 14415 12223
rect 16681 12189 16715 12223
rect 17417 12189 17451 12223
rect 17601 12189 17635 12223
rect 20085 12189 20119 12223
rect 21364 12189 21398 12223
rect 24777 12189 24811 12223
rect 24961 12189 24995 12223
rect 25053 12189 25087 12223
rect 26065 12189 26099 12223
rect 26525 12189 26559 12223
rect 26709 12189 26743 12223
rect 26801 12189 26835 12223
rect 26985 12189 27019 12223
rect 27077 12189 27111 12223
rect 27721 12189 27755 12223
rect 28365 12189 28399 12223
rect 28458 12189 28492 12223
rect 28830 12189 28864 12223
rect 31769 12189 31803 12223
rect 32025 12189 32059 12223
rect 35449 12189 35483 12223
rect 35633 12189 35667 12223
rect 36921 12189 36955 12223
rect 38669 12189 38703 12223
rect 39037 12189 39071 12223
rect 40049 12189 40083 12223
rect 40233 12189 40267 12223
rect 41337 12189 41371 12223
rect 41593 12189 41627 12223
rect 2605 12121 2639 12155
rect 2789 12121 2823 12155
rect 4230 12121 4264 12155
rect 10333 12121 10367 12155
rect 14648 12121 14682 12155
rect 20361 12121 20395 12155
rect 25789 12121 25823 12155
rect 28641 12121 28675 12155
rect 28733 12121 28767 12155
rect 38853 12121 38887 12155
rect 38945 12121 38979 12155
rect 1961 12053 1995 12087
rect 5365 12053 5399 12087
rect 8309 12053 8343 12087
rect 10793 12053 10827 12087
rect 12265 12053 12299 12087
rect 15761 12053 15795 12087
rect 16497 12053 16531 12087
rect 16589 12053 16623 12087
rect 16865 12053 16899 12087
rect 25973 12053 26007 12087
rect 33149 12053 33183 12087
rect 40417 12053 40451 12087
rect 42717 12053 42751 12087
rect 3433 11849 3467 11883
rect 3893 11849 3927 11883
rect 7297 11849 7331 11883
rect 10241 11849 10275 11883
rect 15577 11849 15611 11883
rect 17065 11849 17099 11883
rect 17233 11849 17267 11883
rect 22201 11849 22235 11883
rect 28549 11849 28583 11883
rect 29929 11849 29963 11883
rect 40141 11849 40175 11883
rect 2605 11781 2639 11815
rect 2789 11781 2823 11815
rect 15945 11781 15979 11815
rect 16865 11781 16899 11815
rect 20177 11781 20211 11815
rect 39773 11781 39807 11815
rect 39865 11781 39899 11815
rect 1593 11713 1627 11747
rect 3801 11713 3835 11747
rect 4905 11713 4939 11747
rect 5089 11713 5123 11747
rect 7205 11713 7239 11747
rect 8125 11713 8159 11747
rect 8309 11713 8343 11747
rect 9873 11713 9907 11747
rect 15761 11713 15795 11747
rect 16037 11713 16071 11747
rect 17693 11713 17727 11747
rect 17877 11713 17911 11747
rect 20085 11713 20119 11747
rect 20269 11713 20303 11747
rect 22017 11713 22051 11747
rect 22201 11713 22235 11747
rect 25881 11713 25915 11747
rect 27425 11713 27459 11747
rect 29745 11713 29779 11747
rect 30021 11713 30055 11747
rect 37841 11713 37875 11747
rect 38577 11713 38611 11747
rect 38761 11713 38795 11747
rect 38853 11713 38887 11747
rect 39589 11713 39623 11747
rect 39957 11713 39991 11747
rect 1777 11645 1811 11679
rect 3985 11645 4019 11679
rect 9965 11645 9999 11679
rect 20729 11645 20763 11679
rect 25513 11645 25547 11679
rect 25697 11645 25731 11679
rect 25789 11645 25823 11679
rect 25973 11645 26007 11679
rect 27169 11645 27203 11679
rect 5273 11577 5307 11611
rect 38577 11577 38611 11611
rect 8125 11509 8159 11543
rect 9873 11509 9907 11543
rect 17049 11509 17083 11543
rect 17693 11509 17727 11543
rect 29745 11509 29779 11543
rect 38025 11509 38059 11543
rect 4997 11305 5031 11339
rect 5273 11305 5307 11339
rect 13001 11305 13035 11339
rect 30389 11305 30423 11339
rect 39405 11305 39439 11339
rect 3065 11237 3099 11271
rect 10333 11237 10367 11271
rect 32597 11237 32631 11271
rect 42717 11237 42751 11271
rect 4997 11169 5031 11203
rect 7849 11169 7883 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 15853 11169 15887 11203
rect 16037 11169 16071 11203
rect 22385 11169 22419 11203
rect 38117 11169 38151 11203
rect 44281 11169 44315 11203
rect 1685 11101 1719 11135
rect 4905 11101 4939 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 8401 11101 8435 11135
rect 9689 11101 9723 11135
rect 10057 11101 10091 11135
rect 10425 11101 10459 11135
rect 11621 11101 11655 11135
rect 14473 11101 14507 11135
rect 16129 11101 16163 11135
rect 16221 11101 16255 11135
rect 16313 11101 16347 11135
rect 18429 11101 18463 11135
rect 18613 11101 18647 11135
rect 21373 11101 21407 11135
rect 21649 11101 21683 11135
rect 22109 11101 22143 11135
rect 24961 11101 24995 11135
rect 25237 11101 25271 11135
rect 29837 11101 29871 11135
rect 30205 11101 30239 11135
rect 32781 11101 32815 11135
rect 32873 11101 32907 11135
rect 37657 11101 37691 11135
rect 37841 11101 37875 11135
rect 38853 11101 38887 11135
rect 39129 11101 39163 11135
rect 39221 11101 39255 11135
rect 41337 11101 41371 11135
rect 44097 11101 44131 11135
rect 1952 11033 1986 11067
rect 11888 11033 11922 11067
rect 15209 11033 15243 11067
rect 21557 11033 21591 11067
rect 30021 11033 30055 11067
rect 30113 11033 30147 11067
rect 32597 11033 32631 11067
rect 37749 11033 37783 11067
rect 37959 11033 37993 11067
rect 39037 11033 39071 11067
rect 41604 11033 41638 11067
rect 44189 11033 44223 11067
rect 7021 10965 7055 10999
rect 18521 10965 18555 10999
rect 21189 10965 21223 10999
rect 24777 10965 24811 10999
rect 25145 10965 25179 10999
rect 37473 10965 37507 10999
rect 43729 10965 43763 10999
rect 1961 10761 1995 10795
rect 2329 10761 2363 10795
rect 12265 10761 12299 10795
rect 12633 10761 12667 10795
rect 19533 10761 19567 10795
rect 25237 10761 25271 10795
rect 25697 10761 25731 10795
rect 30481 10761 30515 10795
rect 37749 10761 37783 10795
rect 42993 10761 43027 10795
rect 44281 10761 44315 10795
rect 2421 10693 2455 10727
rect 5825 10693 5859 10727
rect 8033 10693 8067 10727
rect 9413 10693 9447 10727
rect 15209 10693 15243 10727
rect 17141 10693 17175 10727
rect 24124 10693 24158 10727
rect 30113 10693 30147 10727
rect 30205 10693 30239 10727
rect 31217 10693 31251 10727
rect 40938 10693 40972 10727
rect 43361 10693 43395 10727
rect 3249 10625 3283 10659
rect 5549 10625 5583 10659
rect 5733 10625 5767 10659
rect 10149 10625 10183 10659
rect 12449 10625 12483 10659
rect 12725 10625 12759 10659
rect 14473 10625 14507 10659
rect 16865 10625 16899 10659
rect 18420 10625 18454 10659
rect 23857 10625 23891 10659
rect 26065 10625 26099 10659
rect 26157 10625 26191 10659
rect 29929 10625 29963 10659
rect 30297 10625 30331 10659
rect 31125 10625 31159 10659
rect 31309 10625 31343 10659
rect 31447 10625 31481 10659
rect 32321 10625 32355 10659
rect 33977 10625 34011 10659
rect 34161 10625 34195 10659
rect 38117 10625 38151 10659
rect 43177 10625 43211 10659
rect 43269 10625 43303 10659
rect 43479 10625 43513 10659
rect 44189 10625 44223 10659
rect 2513 10557 2547 10591
rect 7297 10557 7331 10591
rect 7389 10557 7423 10591
rect 7481 10557 7515 10591
rect 8769 10557 8803 10591
rect 18153 10557 18187 10591
rect 25881 10557 25915 10591
rect 25973 10557 26007 10591
rect 31585 10557 31619 10591
rect 32505 10557 32539 10591
rect 38209 10557 38243 10591
rect 38393 10557 38427 10591
rect 40693 10557 40727 10591
rect 43637 10557 43671 10591
rect 3341 10421 3375 10455
rect 7113 10421 7147 10455
rect 30941 10421 30975 10455
rect 33977 10421 34011 10455
rect 42073 10421 42107 10455
rect 22385 10217 22419 10251
rect 24593 10217 24627 10251
rect 27261 10217 27295 10251
rect 28457 10217 28491 10251
rect 36737 10217 36771 10251
rect 43177 10217 43211 10251
rect 16589 10149 16623 10183
rect 18429 10149 18463 10183
rect 27905 10149 27939 10183
rect 28641 10149 28675 10183
rect 39037 10149 39071 10183
rect 2973 10081 3007 10115
rect 3065 10081 3099 10115
rect 7481 10081 7515 10115
rect 12357 10081 12391 10115
rect 16773 10081 16807 10115
rect 16957 10081 16991 10115
rect 21005 10081 21039 10115
rect 30849 10081 30883 10115
rect 32045 10081 32079 10115
rect 35357 10081 35391 10115
rect 43729 10081 43763 10115
rect 1593 10013 1627 10047
rect 6009 10013 6043 10047
rect 7113 10013 7147 10047
rect 7849 10013 7883 10047
rect 9505 10013 9539 10047
rect 10517 10013 10551 10047
rect 10977 10013 11011 10047
rect 14473 10013 14507 10047
rect 14749 10013 14783 10047
rect 16865 10013 16899 10047
rect 17049 10013 17083 10047
rect 18613 10013 18647 10047
rect 18889 10013 18923 10047
rect 19441 10013 19475 10047
rect 21272 10013 21306 10047
rect 24777 10013 24811 10047
rect 24869 10013 24903 10047
rect 27169 10013 27203 10047
rect 27353 10013 27387 10047
rect 30113 10013 30147 10047
rect 32301 10013 32335 10047
rect 37197 10013 37231 10047
rect 37464 10013 37498 10047
rect 39313 10013 39347 10047
rect 1869 9945 1903 9979
rect 6561 9945 6595 9979
rect 9781 9945 9815 9979
rect 12624 9945 12658 9979
rect 14289 9945 14323 9979
rect 19717 9945 19751 9979
rect 25329 9945 25363 9979
rect 28273 9945 28307 9979
rect 28489 9945 28523 9979
rect 35602 9945 35636 9979
rect 39037 9945 39071 9979
rect 39221 9945 39255 9979
rect 2513 9877 2547 9911
rect 2881 9877 2915 9911
rect 13737 9877 13771 9911
rect 14657 9877 14691 9911
rect 18797 9877 18831 9911
rect 33425 9877 33459 9911
rect 38577 9877 38611 9911
rect 43545 9877 43579 9911
rect 43637 9877 43671 9911
rect 8217 9673 8251 9707
rect 39405 9673 39439 9707
rect 7021 9605 7055 9639
rect 9413 9605 9447 9639
rect 9618 9605 9652 9639
rect 10701 9605 10735 9639
rect 17110 9605 17144 9639
rect 20913 9605 20947 9639
rect 25145 9605 25179 9639
rect 25973 9605 26007 9639
rect 29009 9605 29043 9639
rect 30113 9605 30147 9639
rect 36001 9605 36035 9639
rect 39957 9605 39991 9639
rect 40938 9605 40972 9639
rect 2145 9537 2179 9571
rect 2412 9537 2446 9571
rect 4629 9537 4663 9571
rect 4896 9537 4930 9571
rect 6653 9537 6687 9571
rect 8125 9537 8159 9571
rect 8493 9537 8527 9571
rect 10333 9537 10367 9571
rect 12173 9537 12207 9571
rect 12265 9537 12299 9571
rect 15301 9537 15335 9571
rect 15485 9537 15519 9571
rect 21005 9537 21039 9571
rect 22385 9537 22419 9571
rect 22477 9537 22511 9571
rect 25329 9537 25363 9571
rect 26249 9537 26283 9571
rect 26341 9537 26375 9571
rect 26433 9537 26467 9571
rect 26617 9537 26651 9571
rect 27445 9537 27479 9571
rect 27538 9537 27572 9571
rect 27721 9537 27755 9571
rect 27813 9537 27847 9571
rect 27951 9537 27985 9571
rect 28641 9537 28675 9571
rect 31493 9537 31527 9571
rect 31677 9537 31711 9571
rect 32321 9537 32355 9571
rect 32505 9537 32539 9571
rect 33793 9537 33827 9571
rect 38853 9537 38887 9571
rect 39037 9537 39071 9571
rect 39129 9537 39163 9571
rect 39221 9537 39255 9571
rect 39865 9537 39899 9571
rect 40049 9537 40083 9571
rect 8309 9469 8343 9503
rect 16865 9469 16899 9503
rect 22201 9469 22235 9503
rect 22293 9469 22327 9503
rect 30941 9469 30975 9503
rect 33885 9469 33919 9503
rect 34069 9469 34103 9503
rect 36737 9469 36771 9503
rect 40693 9469 40727 9503
rect 6009 9401 6043 9435
rect 28089 9401 28123 9435
rect 42073 9401 42107 9435
rect 3525 9333 3559 9367
rect 8401 9333 8435 9367
rect 9597 9333 9631 9367
rect 9781 9333 9815 9367
rect 11989 9333 12023 9367
rect 12449 9333 12483 9367
rect 15393 9333 15427 9367
rect 18245 9333 18279 9367
rect 20729 9333 20763 9367
rect 21189 9333 21223 9367
rect 22017 9333 22051 9367
rect 25513 9333 25547 9367
rect 31493 9333 31527 9367
rect 32321 9333 32355 9367
rect 33425 9333 33459 9367
rect 2513 9129 2547 9163
rect 3249 9129 3283 9163
rect 5457 9129 5491 9163
rect 7481 9129 7515 9163
rect 8125 9129 8159 9163
rect 1869 9061 1903 9095
rect 12817 9061 12851 9095
rect 16405 9061 16439 9095
rect 17785 9061 17819 9095
rect 21281 9061 21315 9095
rect 21465 8993 21499 9027
rect 21649 8993 21683 9027
rect 37197 8993 37231 9027
rect 40233 8993 40267 9027
rect 2421 8925 2455 8959
rect 3157 8925 3191 8959
rect 5641 8925 5675 8959
rect 5917 8925 5951 8959
rect 8125 8925 8159 8959
rect 9873 8925 9907 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 11437 8925 11471 8959
rect 16589 8925 16623 8959
rect 16681 8925 16715 8959
rect 16957 8925 16991 8959
rect 19441 8925 19475 8959
rect 21557 8925 21591 8959
rect 21741 8925 21775 8959
rect 26249 8925 26283 8959
rect 26525 8925 26559 8959
rect 28365 8925 28399 8959
rect 29745 8925 29779 8959
rect 31953 8925 31987 8959
rect 36461 8925 36495 8959
rect 40049 8925 40083 8959
rect 1685 8857 1719 8891
rect 7297 8857 7331 8891
rect 7497 8857 7531 8891
rect 10609 8857 10643 8891
rect 11704 8857 11738 8891
rect 17049 8857 17083 8891
rect 17601 8857 17635 8891
rect 19717 8857 19751 8891
rect 28641 8857 28675 8891
rect 30012 8857 30046 8891
rect 31585 8857 31619 8891
rect 31769 8857 31803 8891
rect 35633 8857 35667 8891
rect 5825 8789 5859 8823
rect 7665 8789 7699 8823
rect 26065 8789 26099 8823
rect 26433 8789 26467 8823
rect 31125 8789 31159 8823
rect 35909 8789 35943 8823
rect 8769 8585 8803 8619
rect 10609 8585 10643 8619
rect 12081 8585 12115 8619
rect 13829 8585 13863 8619
rect 17049 8585 17083 8619
rect 19901 8585 19935 8619
rect 24041 8585 24075 8619
rect 39497 8585 39531 8619
rect 2605 8517 2639 8551
rect 2789 8517 2823 8551
rect 12633 8517 12667 8551
rect 32873 8517 32907 8551
rect 33609 8517 33643 8551
rect 36461 8517 36495 8551
rect 39313 8517 39347 8551
rect 1593 8449 1627 8483
rect 5273 8449 5307 8483
rect 7297 8449 7331 8483
rect 7757 8449 7791 8483
rect 8978 8449 9012 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 12725 8449 12759 8483
rect 14105 8449 14139 8483
rect 14197 8449 14231 8483
rect 14841 8449 14875 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 18153 8449 18187 8483
rect 18245 8449 18279 8483
rect 18337 8449 18371 8483
rect 20361 8449 20395 8483
rect 21097 8449 21131 8483
rect 21281 8449 21315 8483
rect 22661 8449 22695 8483
rect 22917 8449 22951 8483
rect 25145 8449 25179 8483
rect 25412 8449 25446 8483
rect 32413 8449 32447 8483
rect 33333 8449 33367 8483
rect 35449 8449 35483 8483
rect 35541 8449 35575 8483
rect 35633 8449 35667 8483
rect 35817 8449 35851 8483
rect 36277 8449 36311 8483
rect 36553 8449 36587 8483
rect 36645 8449 36679 8483
rect 37657 8449 37691 8483
rect 39589 8449 39623 8483
rect 40233 8449 40267 8483
rect 40877 8449 40911 8483
rect 41061 8449 41095 8483
rect 1777 8381 1811 8415
rect 5089 8381 5123 8415
rect 7941 8381 7975 8415
rect 8493 8381 8527 8415
rect 8861 8381 8895 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 11713 8381 11747 8415
rect 14013 8381 14047 8415
rect 14289 8381 14323 8415
rect 15117 8381 15151 8415
rect 18797 8381 18831 8415
rect 20085 8381 20119 8415
rect 20177 8381 20211 8415
rect 20269 8381 20303 8415
rect 21189 8381 21223 8415
rect 21373 8381 21407 8415
rect 32321 8381 32355 8415
rect 37473 8381 37507 8415
rect 40049 8381 40083 8415
rect 40417 8381 40451 8415
rect 40969 8381 41003 8415
rect 5457 8313 5491 8347
rect 9137 8313 9171 8347
rect 20913 8313 20947 8347
rect 26525 8313 26559 8347
rect 36829 8313 36863 8347
rect 39313 8313 39347 8347
rect 10241 8245 10275 8279
rect 35173 8245 35207 8279
rect 37841 8245 37875 8279
rect 3065 8041 3099 8075
rect 5365 8041 5399 8075
rect 11069 8041 11103 8075
rect 18337 8041 18371 8075
rect 21649 8041 21683 8075
rect 22385 8041 22419 8075
rect 27261 8041 27295 8075
rect 10241 7973 10275 8007
rect 23305 7973 23339 8007
rect 31769 7973 31803 8007
rect 13645 7905 13679 7939
rect 19441 7905 19475 7939
rect 23581 7905 23615 7939
rect 23673 7905 23707 7939
rect 25881 7905 25915 7939
rect 35173 7905 35207 7939
rect 35357 7905 35391 7939
rect 1685 7837 1719 7871
rect 3985 7837 4019 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 10057 7837 10091 7871
rect 10977 7837 11011 7871
rect 13369 7837 13403 7871
rect 13461 7837 13495 7871
rect 13553 7837 13587 7871
rect 14381 7837 14415 7871
rect 14565 7837 14599 7871
rect 18521 7837 18555 7871
rect 18613 7837 18647 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 23489 7837 23523 7871
rect 23765 7837 23799 7871
rect 26148 7837 26182 7871
rect 31585 7837 31619 7871
rect 31677 7837 31711 7871
rect 32321 7837 32355 7871
rect 32597 7837 32631 7871
rect 32689 7837 32723 7871
rect 33333 7837 33367 7871
rect 35081 7837 35115 7871
rect 35265 7837 35299 7871
rect 36001 7837 36035 7871
rect 36268 7837 36302 7871
rect 40049 7837 40083 7871
rect 40417 7837 40451 7871
rect 41245 7837 41279 7871
rect 41512 7837 41546 7871
rect 1952 7769 1986 7803
rect 4252 7769 4286 7803
rect 7849 7769 7883 7803
rect 14473 7769 14507 7803
rect 15025 7769 15059 7803
rect 19686 7769 19720 7803
rect 21373 7769 21407 7803
rect 22753 7769 22787 7803
rect 32505 7769 32539 7803
rect 33609 7769 33643 7803
rect 40233 7769 40267 7803
rect 40325 7769 40359 7803
rect 13185 7701 13219 7735
rect 20821 7701 20855 7735
rect 32873 7701 32907 7735
rect 34897 7701 34931 7735
rect 37381 7701 37415 7735
rect 40601 7701 40635 7735
rect 42625 7701 42659 7735
rect 1961 7497 1995 7531
rect 2329 7497 2363 7531
rect 2421 7497 2455 7531
rect 3341 7497 3375 7531
rect 4537 7497 4571 7531
rect 4905 7497 4939 7531
rect 9413 7497 9447 7531
rect 14841 7497 14875 7531
rect 19165 7497 19199 7531
rect 19533 7497 19567 7531
rect 32413 7497 32447 7531
rect 33517 7497 33551 7531
rect 37749 7497 37783 7531
rect 3249 7429 3283 7463
rect 11713 7429 11747 7463
rect 11929 7429 11963 7463
rect 4721 7361 4755 7395
rect 4997 7361 5031 7395
rect 7021 7361 7055 7395
rect 9321 7361 9355 7395
rect 10701 7361 10735 7395
rect 15025 7361 15059 7395
rect 15209 7361 15243 7395
rect 19349 7361 19383 7395
rect 19625 7361 19659 7395
rect 22937 7361 22971 7395
rect 32597 7361 32631 7395
rect 32689 7361 32723 7395
rect 32965 7361 32999 7395
rect 33425 7361 33459 7395
rect 33609 7361 33643 7395
rect 38117 7361 38151 7395
rect 42809 7361 42843 7395
rect 2513 7293 2547 7327
rect 7113 7293 7147 7327
rect 9597 7293 9631 7327
rect 10885 7293 10919 7327
rect 15117 7293 15151 7327
rect 15301 7293 15335 7327
rect 23029 7293 23063 7327
rect 23121 7293 23155 7327
rect 23213 7293 23247 7327
rect 38209 7293 38243 7327
rect 38393 7293 38427 7327
rect 42625 7293 42659 7327
rect 7297 7157 7331 7191
rect 8953 7157 8987 7191
rect 11897 7157 11931 7191
rect 12081 7157 12115 7191
rect 22753 7157 22787 7191
rect 32873 7157 32907 7191
rect 42993 7157 43027 7191
rect 16681 6953 16715 6987
rect 2697 6817 2731 6851
rect 4261 6817 4295 6851
rect 22017 6817 22051 6851
rect 24685 6817 24719 6851
rect 30021 6817 30055 6851
rect 30941 6817 30975 6851
rect 31309 6817 31343 6851
rect 36645 6817 36679 6851
rect 4077 6749 4111 6783
rect 8125 6749 8159 6783
rect 10149 6749 10183 6783
rect 11529 6749 11563 6783
rect 15301 6749 15335 6783
rect 17325 6749 17359 6783
rect 17601 6749 17635 6783
rect 22284 6749 22318 6783
rect 24593 6749 24627 6783
rect 29745 6749 29779 6783
rect 29929 6749 29963 6783
rect 30113 6749 30147 6783
rect 30297 6749 30331 6783
rect 31125 6749 31159 6783
rect 31217 6749 31251 6783
rect 31401 6749 31435 6783
rect 32045 6749 32079 6783
rect 32229 6749 32263 6783
rect 32873 6749 32907 6783
rect 33140 6749 33174 6783
rect 35541 6749 35575 6783
rect 35633 6749 35667 6783
rect 41337 6749 41371 6783
rect 41604 6749 41638 6783
rect 44005 6749 44039 6783
rect 44097 6749 44131 6783
rect 44189 6749 44223 6783
rect 44373 6749 44407 6783
rect 8401 6681 8435 6715
rect 10885 6681 10919 6715
rect 11796 6681 11830 6715
rect 15568 6681 15602 6715
rect 17141 6681 17175 6715
rect 32321 6681 32355 6715
rect 36277 6681 36311 6715
rect 36461 6681 36495 6715
rect 2145 6613 2179 6647
rect 2513 6613 2547 6647
rect 2605 6613 2639 6647
rect 12909 6613 12943 6647
rect 17509 6613 17543 6647
rect 23397 6613 23431 6647
rect 30481 6613 30515 6647
rect 34253 6613 34287 6647
rect 35817 6613 35851 6647
rect 42717 6613 42751 6647
rect 43729 6613 43763 6647
rect 8493 6409 8527 6443
rect 10333 6409 10367 6443
rect 11805 6409 11839 6443
rect 38209 6409 38243 6443
rect 42625 6409 42659 6443
rect 44281 6409 44315 6443
rect 2136 6341 2170 6375
rect 4077 6341 4111 6375
rect 7297 6341 7331 6375
rect 13921 6341 13955 6375
rect 14121 6341 14155 6375
rect 22385 6341 22419 6375
rect 37933 6341 37967 6375
rect 43913 6341 43947 6375
rect 3801 6273 3835 6307
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 9413 6273 9447 6307
rect 9781 6273 9815 6307
rect 10517 6273 10551 6307
rect 10609 6273 10643 6307
rect 10701 6273 10735 6307
rect 10839 6273 10873 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 12265 6273 12299 6307
rect 19349 6273 19383 6307
rect 22017 6273 22051 6307
rect 22110 6273 22144 6307
rect 22293 6273 22327 6307
rect 22523 6273 22557 6307
rect 25329 6273 25363 6307
rect 25513 6273 25547 6307
rect 25605 6273 25639 6307
rect 28273 6273 28307 6307
rect 28540 6273 28574 6307
rect 33977 6273 34011 6307
rect 34069 6273 34103 6307
rect 37657 6273 37691 6307
rect 37841 6273 37875 6307
rect 38025 6273 38059 6307
rect 38925 6273 38959 6307
rect 42901 6273 42935 6307
rect 42993 6273 43027 6307
rect 43085 6273 43119 6307
rect 44097 6273 44131 6307
rect 1869 6205 1903 6239
rect 8585 6205 8619 6239
rect 8677 6205 8711 6239
rect 10977 6205 11011 6239
rect 19073 6205 19107 6239
rect 19165 6205 19199 6239
rect 19257 6205 19291 6239
rect 38669 6205 38703 6239
rect 42809 6205 42843 6239
rect 3249 6137 3283 6171
rect 22661 6137 22695 6171
rect 34253 6137 34287 6171
rect 5181 6069 5215 6103
rect 8125 6069 8159 6103
rect 14105 6069 14139 6103
rect 14289 6069 14323 6103
rect 18889 6069 18923 6103
rect 25145 6069 25179 6103
rect 29653 6069 29687 6103
rect 40049 6069 40083 6103
rect 4169 5865 4203 5899
rect 7021 5865 7055 5899
rect 7941 5865 7975 5899
rect 12357 5865 12391 5899
rect 18797 5865 18831 5899
rect 23029 5865 23063 5899
rect 40601 5865 40635 5899
rect 1777 5729 1811 5763
rect 5457 5729 5491 5763
rect 10425 5729 10459 5763
rect 19441 5729 19475 5763
rect 25973 5729 26007 5763
rect 33885 5729 33919 5763
rect 41153 5729 41187 5763
rect 43637 5729 43671 5763
rect 1593 5661 1627 5695
rect 2697 5661 2731 5695
rect 5733 5661 5767 5695
rect 8217 5661 8251 5695
rect 10149 5661 10183 5695
rect 11069 5661 11103 5695
rect 11162 5661 11196 5695
rect 11437 5661 11471 5695
rect 11534 5661 11568 5695
rect 14473 5661 14507 5695
rect 14749 5661 14783 5695
rect 18429 5661 18463 5695
rect 19697 5661 19731 5695
rect 22845 5661 22879 5695
rect 26229 5661 26263 5695
rect 30297 5661 30331 5695
rect 33425 5661 33459 5695
rect 33609 5661 33643 5695
rect 33747 5661 33781 5695
rect 36369 5661 36403 5695
rect 36625 5661 36659 5695
rect 40049 5661 40083 5695
rect 40233 5661 40267 5695
rect 40417 5661 40451 5695
rect 43177 5661 43211 5695
rect 43479 5661 43513 5695
rect 3065 5593 3099 5627
rect 4077 5593 4111 5627
rect 4813 5593 4847 5627
rect 7573 5593 7607 5627
rect 11345 5593 11379 5627
rect 12173 5593 12207 5627
rect 12373 5593 12407 5627
rect 14657 5593 14691 5627
rect 18613 5593 18647 5627
rect 22661 5593 22695 5627
rect 30542 5593 30576 5627
rect 33517 5593 33551 5627
rect 40325 5593 40359 5627
rect 41420 5593 41454 5627
rect 42993 5593 43027 5627
rect 43269 5593 43303 5627
rect 43361 5593 43395 5627
rect 4905 5525 4939 5559
rect 7950 5525 7984 5559
rect 11713 5525 11747 5559
rect 12541 5525 12575 5559
rect 14289 5525 14323 5559
rect 20821 5525 20855 5559
rect 27353 5525 27387 5559
rect 31677 5525 31711 5559
rect 33241 5525 33275 5559
rect 37749 5525 37783 5559
rect 42533 5525 42567 5559
rect 14657 5321 14691 5355
rect 18797 5321 18831 5355
rect 23949 5321 23983 5355
rect 27813 5321 27847 5355
rect 30481 5321 30515 5355
rect 35357 5321 35391 5355
rect 36277 5321 36311 5355
rect 44097 5321 44131 5355
rect 45201 5321 45235 5355
rect 5917 5253 5951 5287
rect 8033 5253 8067 5287
rect 8217 5253 8251 5287
rect 16865 5253 16899 5287
rect 17081 5253 17115 5287
rect 23765 5253 23799 5287
rect 24133 5253 24167 5287
rect 27445 5253 27479 5287
rect 34222 5253 34256 5287
rect 41521 5253 41555 5287
rect 1593 5185 1627 5219
rect 2513 5185 2547 5219
rect 3893 5185 3927 5219
rect 4169 5185 4203 5219
rect 4353 5185 4387 5219
rect 5365 5185 5399 5219
rect 6745 5185 6779 5219
rect 10701 5185 10735 5219
rect 10885 5185 10919 5219
rect 10977 5185 11011 5219
rect 13277 5185 13311 5219
rect 13544 5185 13578 5219
rect 15761 5185 15795 5219
rect 16037 5185 16071 5219
rect 18613 5185 18647 5219
rect 18797 5185 18831 5219
rect 22661 5185 22695 5219
rect 22845 5185 22879 5219
rect 24041 5185 24075 5219
rect 24501 5185 24535 5219
rect 27169 5185 27203 5219
rect 27317 5185 27351 5219
rect 27537 5185 27571 5219
rect 27634 5185 27668 5219
rect 29745 5185 29779 5219
rect 29929 5185 29963 5219
rect 30113 5185 30147 5219
rect 30297 5185 30331 5219
rect 41337 5185 41371 5219
rect 41429 5185 41463 5219
rect 41639 5185 41673 5219
rect 41797 5185 41831 5219
rect 44005 5185 44039 5219
rect 1777 5117 1811 5151
rect 6561 5117 6595 5151
rect 6929 5117 6963 5151
rect 7021 5117 7055 5151
rect 15853 5117 15887 5151
rect 30021 5117 30055 5151
rect 33977 5117 34011 5151
rect 36369 5117 36403 5151
rect 36553 5117 36587 5151
rect 44189 5117 44223 5151
rect 45293 5117 45327 5151
rect 45385 5117 45419 5151
rect 2697 5049 2731 5083
rect 15945 5049 15979 5083
rect 17233 5049 17267 5083
rect 22661 5049 22695 5083
rect 35909 5049 35943 5083
rect 43637 5049 43671 5083
rect 3709 4981 3743 5015
rect 8401 4981 8435 5015
rect 10517 4981 10551 5015
rect 15577 4981 15611 5015
rect 17049 4981 17083 5015
rect 41153 4981 41187 5015
rect 44833 4981 44867 5015
rect 3065 4777 3099 4811
rect 5089 4777 5123 4811
rect 8585 4777 8619 4811
rect 11621 4777 11655 4811
rect 16037 4777 16071 4811
rect 22109 4777 22143 4811
rect 22753 4777 22787 4811
rect 27537 4777 27571 4811
rect 30297 4777 30331 4811
rect 22293 4709 22327 4743
rect 38761 4709 38795 4743
rect 19717 4641 19751 4675
rect 20545 4641 20579 4675
rect 26157 4641 26191 4675
rect 29929 4641 29963 4675
rect 39313 4641 39347 4675
rect 1685 4573 1719 4607
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 7205 4573 7239 4607
rect 10241 4573 10275 4607
rect 10508 4573 10542 4607
rect 16221 4573 16255 4607
rect 16313 4573 16347 4607
rect 19625 4573 19659 4607
rect 19809 4573 19843 4607
rect 19901 4573 19935 4607
rect 20453 4573 20487 4607
rect 23029 4573 23063 4607
rect 30113 4573 30147 4607
rect 37841 4573 37875 4607
rect 38025 4573 38059 4607
rect 38143 4573 38177 4607
rect 38301 4573 38335 4607
rect 41613 4573 41647 4607
rect 41705 4573 41739 4607
rect 41797 4573 41831 4607
rect 42073 4573 42107 4607
rect 1952 4505 1986 4539
rect 4077 4505 4111 4539
rect 6285 4505 6319 4539
rect 7472 4505 7506 4539
rect 16037 4505 16071 4539
rect 17969 4505 18003 4539
rect 18245 4505 18279 4539
rect 18337 4505 18371 4539
rect 18705 4505 18739 4539
rect 21925 4505 21959 4539
rect 22125 4505 22159 4539
rect 22753 4505 22787 4539
rect 26424 4505 26458 4539
rect 37933 4505 37967 4539
rect 41915 4505 41949 4539
rect 4169 4437 4203 4471
rect 6377 4437 6411 4471
rect 18153 4437 18187 4471
rect 19441 4437 19475 4471
rect 22937 4437 22971 4471
rect 37657 4437 37691 4471
rect 39129 4437 39163 4471
rect 39221 4437 39255 4471
rect 41429 4437 41463 4471
rect 3433 4233 3467 4267
rect 44005 4233 44039 4267
rect 4261 4165 4295 4199
rect 17233 4165 17267 4199
rect 17877 4165 17911 4199
rect 34713 4165 34747 4199
rect 38853 4165 38887 4199
rect 42993 4165 43027 4199
rect 43111 4165 43145 4199
rect 44373 4165 44407 4199
rect 45569 4165 45603 4199
rect 1593 4097 1627 4131
rect 2513 4097 2547 4131
rect 3249 4097 3283 4131
rect 4077 4097 4111 4131
rect 4721 4097 4755 4131
rect 4905 4097 4939 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 6929 4097 6963 4131
rect 11897 4097 11931 4131
rect 11990 4097 12024 4131
rect 12173 4097 12207 4131
rect 12265 4097 12299 4131
rect 12403 4097 12437 4131
rect 14657 4097 14691 4131
rect 14841 4097 14875 4131
rect 18061 4097 18095 4131
rect 18245 4097 18279 4131
rect 20361 4097 20395 4131
rect 23765 4097 23799 4131
rect 29285 4097 29319 4131
rect 29469 4097 29503 4131
rect 29837 4097 29871 4131
rect 30021 4097 30055 4131
rect 30941 4097 30975 4131
rect 31034 4097 31068 4131
rect 31217 4097 31251 4131
rect 31309 4097 31343 4131
rect 31447 4097 31481 4131
rect 33057 4097 33091 4131
rect 39037 4097 39071 4131
rect 42809 4097 42843 4131
rect 42901 4097 42935 4131
rect 44465 4097 44499 4131
rect 45661 4097 45695 4131
rect 1777 4029 1811 4063
rect 5365 4029 5399 4063
rect 5549 4029 5583 4063
rect 7205 4029 7239 4063
rect 8309 4029 8343 4063
rect 20545 4029 20579 4063
rect 23857 4029 23891 4063
rect 29561 4029 29595 4063
rect 29653 4029 29687 4063
rect 32873 4029 32907 4063
rect 34897 4029 34931 4063
rect 43269 4029 43303 4063
rect 44649 4029 44683 4063
rect 45753 4029 45787 4063
rect 2697 3961 2731 3995
rect 4813 3961 4847 3995
rect 31585 3961 31619 3995
rect 45201 3961 45235 3995
rect 12541 3893 12575 3927
rect 14657 3893 14691 3927
rect 17325 3893 17359 3927
rect 24133 3893 24167 3927
rect 33241 3893 33275 3927
rect 42625 3893 42659 3927
rect 1961 3689 1995 3723
rect 2697 3689 2731 3723
rect 7205 3689 7239 3723
rect 11713 3689 11747 3723
rect 16865 3689 16899 3723
rect 17969 3689 18003 3723
rect 21097 3689 21131 3723
rect 30205 3689 30239 3723
rect 39497 3689 39531 3723
rect 42441 3689 42475 3723
rect 4813 3621 4847 3655
rect 6561 3621 6595 3655
rect 27169 3621 27203 3655
rect 29193 3621 29227 3655
rect 40417 3621 40451 3655
rect 7757 3553 7791 3587
rect 10241 3553 10275 3587
rect 19717 3553 19751 3587
rect 27629 3553 27663 3587
rect 31953 3553 31987 3587
rect 35909 3553 35943 3587
rect 2513 3485 2547 3519
rect 3433 3485 3467 3519
rect 4629 3485 4663 3519
rect 4905 3485 4939 3519
rect 5457 3485 5491 3519
rect 5641 3485 5675 3519
rect 7113 3485 7147 3519
rect 8585 3485 8619 3519
rect 10425 3485 10459 3519
rect 12265 3485 12299 3519
rect 12449 3485 12483 3519
rect 12633 3485 12667 3519
rect 13093 3485 13127 3519
rect 13186 3485 13220 3519
rect 13369 3485 13403 3519
rect 13599 3485 13633 3519
rect 16221 3485 16255 3519
rect 16314 3485 16348 3519
rect 16597 3485 16631 3519
rect 16727 3485 16761 3519
rect 17325 3485 17359 3519
rect 17418 3485 17452 3519
rect 17831 3485 17865 3519
rect 20453 3485 20487 3519
rect 20546 3485 20580 3519
rect 20918 3485 20952 3519
rect 22661 3485 22695 3519
rect 23765 3485 23799 3519
rect 24041 3485 24075 3519
rect 25789 3485 25823 3519
rect 27813 3485 27847 3519
rect 28549 3485 28583 3519
rect 28642 3485 28676 3519
rect 28917 3485 28951 3519
rect 29055 3485 29089 3519
rect 30757 3485 30791 3519
rect 30941 3485 30975 3519
rect 31033 3485 31067 3519
rect 31125 3485 31159 3519
rect 31309 3485 31343 3519
rect 35173 3485 35207 3519
rect 35265 3485 35299 3519
rect 38117 3485 38151 3519
rect 38384 3485 38418 3519
rect 41061 3485 41095 3519
rect 41328 3485 41362 3519
rect 57161 3485 57195 3519
rect 1685 3417 1719 3451
rect 6377 3417 6411 3451
rect 10609 3417 10643 3451
rect 11621 3417 11655 3451
rect 13461 3417 13495 3451
rect 14473 3417 14507 3451
rect 16497 3417 16531 3451
rect 17601 3417 17635 3451
rect 17693 3417 17727 3451
rect 19533 3417 19567 3451
rect 20729 3417 20763 3451
rect 20821 3417 20855 3451
rect 21833 3417 21867 3451
rect 22937 3417 22971 3451
rect 26056 3417 26090 3451
rect 27997 3417 28031 3451
rect 28825 3417 28859 3451
rect 30113 3417 30147 3451
rect 31493 3417 31527 3451
rect 32198 3417 32232 3451
rect 35449 3417 35483 3451
rect 36154 3417 36188 3451
rect 40233 3417 40267 3451
rect 57437 3417 57471 3451
rect 4445 3349 4479 3383
rect 5825 3349 5859 3383
rect 13737 3349 13771 3383
rect 14565 3349 14599 3383
rect 21925 3349 21959 3383
rect 23581 3349 23615 3383
rect 23949 3349 23983 3383
rect 33333 3349 33367 3383
rect 37289 3349 37323 3383
rect 4997 3145 5031 3179
rect 21465 3145 21499 3179
rect 23949 3145 23983 3179
rect 27445 3145 27479 3179
rect 28181 3145 28215 3179
rect 30113 3145 30147 3179
rect 35265 3145 35299 3179
rect 37657 3145 37691 3179
rect 39589 3145 39623 3179
rect 42809 3145 42843 3179
rect 43545 3145 43579 3179
rect 44465 3145 44499 3179
rect 45845 3145 45879 3179
rect 47961 3145 47995 3179
rect 54125 3145 54159 3179
rect 55965 3145 55999 3179
rect 8493 3077 8527 3111
rect 10057 3077 10091 3111
rect 14188 3077 14222 3111
rect 19248 3077 19282 3111
rect 28089 3077 28123 3111
rect 31309 3077 31343 3111
rect 32597 3077 32631 3111
rect 33425 3077 33459 3111
rect 37565 3077 37599 3111
rect 42717 3077 42751 3111
rect 56977 3077 57011 3111
rect 1593 3009 1627 3043
rect 2697 3009 2731 3043
rect 3617 3009 3651 3043
rect 3884 3009 3918 3043
rect 5457 3009 5491 3043
rect 5641 3009 5675 3043
rect 7021 3009 7055 3043
rect 8309 3009 8343 3043
rect 9137 3009 9171 3043
rect 9781 3009 9815 3043
rect 10977 3009 11011 3043
rect 12357 3009 12391 3043
rect 13001 3009 13035 3043
rect 13921 3009 13955 3043
rect 15853 3009 15887 3043
rect 17141 3009 17175 3043
rect 18061 3009 18095 3043
rect 18981 3009 19015 3043
rect 20821 3009 20855 3043
rect 20914 3009 20948 3043
rect 21097 3009 21131 3043
rect 21189 3009 21223 3043
rect 21327 3009 21361 3043
rect 22569 3009 22603 3043
rect 22836 3009 22870 3043
rect 24961 3009 24995 3043
rect 27353 3009 27387 3043
rect 29000 3009 29034 3043
rect 30573 3009 30607 3043
rect 30757 3007 30791 3041
rect 30941 3009 30975 3043
rect 31125 3009 31159 3043
rect 32413 3009 32447 3043
rect 33241 3009 33275 3043
rect 33885 3009 33919 3043
rect 34141 3009 34175 3043
rect 36461 3009 36495 3043
rect 38209 3009 38243 3043
rect 38465 3009 38499 3043
rect 40601 3009 40635 3043
rect 40868 3009 40902 3043
rect 43453 3009 43487 3043
rect 44373 3009 44407 3043
rect 45753 3009 45787 3043
rect 47869 3009 47903 3043
rect 48881 3009 48915 3043
rect 50261 3009 50295 3043
rect 51641 3009 51675 3043
rect 54033 3009 54067 3043
rect 54861 3009 54895 3043
rect 55873 3009 55907 3043
rect 56701 3009 56735 3043
rect 1777 2941 1811 2975
rect 2973 2941 3007 2975
rect 7205 2941 7239 2975
rect 8953 2941 8987 2975
rect 10793 2941 10827 2975
rect 12173 2941 12207 2975
rect 13185 2941 13219 2975
rect 16037 2941 16071 2975
rect 17417 2941 17451 2975
rect 18337 2941 18371 2975
rect 25145 2941 25179 2975
rect 28733 2941 28767 2975
rect 30843 2941 30877 2975
rect 36645 2941 36679 2975
rect 49065 2941 49099 2975
rect 50445 2941 50479 2975
rect 51825 2941 51859 2975
rect 55045 2941 55079 2975
rect 5825 2873 5859 2907
rect 11161 2873 11195 2907
rect 41981 2873 42015 2907
rect 9321 2805 9355 2839
rect 12541 2805 12575 2839
rect 15301 2805 15335 2839
rect 20361 2805 20395 2839
rect 35541 2601 35575 2635
rect 38945 2601 38979 2635
rect 53113 2601 53147 2635
rect 24869 2533 24903 2567
rect 26617 2533 26651 2567
rect 50721 2465 50755 2499
rect 2053 2397 2087 2431
rect 2973 2397 3007 2431
rect 4261 2397 4295 2431
rect 5181 2397 5215 2431
rect 7021 2397 7055 2431
rect 7941 2397 7975 2431
rect 9781 2397 9815 2431
rect 10701 2397 10735 2431
rect 12357 2397 12391 2431
rect 13277 2397 13311 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 24685 2397 24719 2431
rect 25421 2397 25455 2431
rect 27169 2397 27203 2431
rect 28181 2397 28215 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 32321 2397 32355 2431
rect 33701 2397 33735 2431
rect 34897 2397 34931 2431
rect 34990 2397 35024 2431
rect 35265 2397 35299 2431
rect 35362 2397 35396 2431
rect 36001 2397 36035 2431
rect 37841 2397 37875 2431
rect 40049 2397 40083 2431
rect 40969 2397 41003 2431
rect 42625 2397 42659 2431
rect 43545 2397 43579 2431
rect 45201 2397 45235 2431
rect 46121 2397 46155 2431
rect 47777 2397 47811 2431
rect 53849 2397 53883 2431
rect 55505 2397 55539 2431
rect 56425 2397 56459 2431
rect 2329 2329 2363 2363
rect 3249 2329 3283 2363
rect 4537 2329 4571 2363
rect 5457 2329 5491 2363
rect 7297 2329 7331 2363
rect 8217 2329 8251 2363
rect 10057 2329 10091 2363
rect 10977 2329 11011 2363
rect 12633 2329 12667 2363
rect 13553 2329 13587 2363
rect 15209 2329 15243 2363
rect 16129 2329 16163 2363
rect 17785 2329 17819 2363
rect 18705 2329 18739 2363
rect 20361 2329 20395 2363
rect 21281 2329 21315 2363
rect 22937 2329 22971 2363
rect 23857 2329 23891 2363
rect 25697 2329 25731 2363
rect 26433 2329 26467 2363
rect 27445 2329 27479 2363
rect 28457 2329 28491 2363
rect 30021 2329 30055 2363
rect 31217 2329 31251 2363
rect 32597 2329 32631 2363
rect 33977 2329 34011 2363
rect 35173 2329 35207 2363
rect 36277 2329 36311 2363
rect 38117 2329 38151 2363
rect 38853 2329 38887 2363
rect 40325 2329 40359 2363
rect 41245 2329 41279 2363
rect 42901 2329 42935 2363
rect 43821 2329 43855 2363
rect 45477 2329 45511 2363
rect 46397 2329 46431 2363
rect 48053 2329 48087 2363
rect 48789 2329 48823 2363
rect 50445 2329 50479 2363
rect 51365 2329 51399 2363
rect 53021 2329 53055 2363
rect 54125 2329 54159 2363
rect 55781 2329 55815 2363
rect 56701 2329 56735 2363
rect 9137 2261 9171 2295
rect 11713 2261 11747 2295
rect 14289 2261 14323 2295
rect 48881 2261 48915 2295
rect 51457 2261 51491 2295
<< metal1 >>
rect 3878 41080 3884 41132
rect 3936 41120 3942 41132
rect 4614 41120 4620 41132
rect 3936 41092 4620 41120
rect 3936 41080 3942 41092
rect 4614 41080 4620 41092
rect 4672 41080 4678 41132
rect 18782 41080 18788 41132
rect 18840 41120 18846 41132
rect 19426 41120 19432 41132
rect 18840 41092 19432 41120
rect 18840 41080 18846 41092
rect 19426 41080 19432 41092
rect 19484 41080 19490 41132
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 41414 39584 41420 39636
rect 41472 39584 41478 39636
rect 48590 39584 48596 39636
rect 48648 39624 48654 39636
rect 48869 39627 48927 39633
rect 48869 39624 48881 39627
rect 48648 39596 48881 39624
rect 48648 39584 48654 39596
rect 48869 39593 48881 39596
rect 48915 39593 48927 39627
rect 48869 39587 48927 39593
rect 934 39448 940 39500
rect 992 39488 998 39500
rect 1765 39491 1823 39497
rect 1765 39488 1777 39491
rect 992 39460 1777 39488
rect 992 39448 998 39460
rect 1765 39457 1777 39460
rect 1811 39457 1823 39491
rect 3418 39488 3424 39500
rect 1765 39451 1823 39457
rect 2424 39460 3424 39488
rect 1581 39423 1639 39429
rect 1581 39389 1593 39423
rect 1627 39420 1639 39423
rect 2424 39420 2452 39460
rect 3418 39448 3424 39460
rect 3476 39448 3482 39500
rect 4249 39491 4307 39497
rect 4249 39457 4261 39491
rect 4295 39488 4307 39491
rect 4614 39488 4620 39500
rect 4295 39460 4620 39488
rect 4295 39457 4307 39460
rect 4249 39451 4307 39457
rect 4614 39448 4620 39460
rect 4672 39448 4678 39500
rect 19426 39448 19432 39500
rect 19484 39448 19490 39500
rect 26234 39448 26240 39500
rect 26292 39488 26298 39500
rect 27341 39491 27399 39497
rect 27341 39488 27353 39491
rect 26292 39460 27353 39488
rect 26292 39448 26298 39460
rect 27341 39457 27353 39460
rect 27387 39457 27399 39491
rect 27341 39451 27399 39457
rect 56042 39448 56048 39500
rect 56100 39488 56106 39500
rect 56321 39491 56379 39497
rect 56321 39488 56333 39491
rect 56100 39460 56333 39488
rect 56100 39448 56106 39460
rect 56321 39457 56333 39460
rect 56367 39457 56379 39491
rect 56321 39451 56379 39457
rect 1627 39392 2452 39420
rect 1627 39389 1639 39392
rect 1581 39383 1639 39389
rect 2498 39380 2504 39432
rect 2556 39380 2562 39432
rect 3973 39423 4031 39429
rect 3973 39389 3985 39423
rect 4019 39420 4031 39423
rect 4019 39392 6914 39420
rect 4019 39389 4031 39392
rect 3973 39383 4031 39389
rect 1026 39312 1032 39364
rect 1084 39352 1090 39364
rect 2777 39355 2835 39361
rect 2777 39352 2789 39355
rect 1084 39324 2789 39352
rect 1084 39312 1090 39324
rect 2777 39321 2789 39324
rect 2823 39321 2835 39355
rect 6886 39352 6914 39392
rect 27154 39380 27160 39432
rect 27212 39380 27218 39432
rect 33686 39380 33692 39432
rect 33744 39420 33750 39432
rect 33873 39423 33931 39429
rect 33873 39420 33885 39423
rect 33744 39392 33885 39420
rect 33744 39380 33750 39392
rect 33873 39389 33885 39392
rect 33919 39389 33931 39423
rect 33873 39383 33931 39389
rect 42150 39380 42156 39432
rect 42208 39420 42214 39432
rect 56137 39423 56195 39429
rect 56137 39420 56149 39423
rect 42208 39392 56149 39420
rect 42208 39380 42214 39392
rect 56137 39389 56149 39392
rect 56183 39389 56195 39423
rect 56137 39383 56195 39389
rect 28258 39352 28264 39364
rect 6886 39324 28264 39352
rect 2777 39315 2835 39321
rect 28258 39312 28264 39324
rect 28316 39312 28322 39364
rect 33318 39244 33324 39296
rect 33376 39284 33382 39296
rect 33965 39287 34023 39293
rect 33965 39284 33977 39287
rect 33376 39256 33977 39284
rect 33376 39244 33382 39256
rect 33965 39253 33977 39256
rect 34011 39253 34023 39287
rect 33965 39247 34023 39253
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 7650 39012 7656 39024
rect 1596 38984 7656 39012
rect 1596 38953 1624 38984
rect 7650 38972 7656 38984
rect 7708 38972 7714 39024
rect 1581 38947 1639 38953
rect 1581 38913 1593 38947
rect 1627 38913 1639 38947
rect 1581 38907 1639 38913
rect 2501 38947 2559 38953
rect 2501 38913 2513 38947
rect 2547 38944 2559 38947
rect 6178 38944 6184 38956
rect 2547 38916 6184 38944
rect 2547 38913 2559 38916
rect 2501 38907 2559 38913
rect 6178 38904 6184 38916
rect 6236 38904 6242 38956
rect 934 38836 940 38888
rect 992 38876 998 38888
rect 1765 38879 1823 38885
rect 1765 38876 1777 38879
rect 992 38848 1777 38876
rect 992 38836 998 38848
rect 1765 38845 1777 38848
rect 1811 38845 1823 38879
rect 1765 38839 1823 38845
rect 2685 38879 2743 38885
rect 2685 38845 2697 38879
rect 2731 38845 2743 38879
rect 2685 38839 2743 38845
rect 1118 38768 1124 38820
rect 1176 38808 1182 38820
rect 2700 38808 2728 38839
rect 1176 38780 2728 38808
rect 1176 38768 1182 38780
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1581 38335 1639 38341
rect 1581 38301 1593 38335
rect 1627 38332 1639 38335
rect 10318 38332 10324 38344
rect 1627 38304 10324 38332
rect 1627 38301 1639 38304
rect 1581 38295 1639 38301
rect 10318 38292 10324 38304
rect 10376 38292 10382 38344
rect 934 38224 940 38276
rect 992 38264 998 38276
rect 1857 38267 1915 38273
rect 1857 38264 1869 38267
rect 992 38236 1869 38264
rect 992 38224 998 38236
rect 1857 38233 1869 38236
rect 1903 38233 1915 38267
rect 1857 38227 1915 38233
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 6178 37884 6184 37936
rect 6236 37924 6242 37936
rect 14274 37924 14280 37936
rect 6236 37896 14280 37924
rect 6236 37884 6242 37896
rect 14274 37884 14280 37896
rect 14332 37884 14338 37936
rect 2498 37612 2504 37664
rect 2556 37652 2562 37664
rect 5994 37652 6000 37664
rect 2556 37624 6000 37652
rect 2556 37612 2562 37624
rect 5994 37612 6000 37624
rect 6052 37612 6058 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 3418 37408 3424 37460
rect 3476 37448 3482 37460
rect 5350 37448 5356 37460
rect 3476 37420 5356 37448
rect 3476 37408 3482 37420
rect 5350 37408 5356 37420
rect 5408 37408 5414 37460
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 4062 37244 4068 37256
rect 1627 37216 4068 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 4062 37204 4068 37216
rect 4120 37204 4126 37256
rect 934 37136 940 37188
rect 992 37176 998 37188
rect 1857 37179 1915 37185
rect 1857 37176 1869 37179
rect 992 37148 1869 37176
rect 992 37136 998 37148
rect 1857 37145 1869 37148
rect 1903 37145 1915 37179
rect 1857 37139 1915 37145
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 11974 36768 11980 36780
rect 1627 36740 11980 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 11974 36728 11980 36740
rect 12032 36728 12038 36780
rect 934 36660 940 36712
rect 992 36700 998 36712
rect 1765 36703 1823 36709
rect 1765 36700 1777 36703
rect 992 36672 1777 36700
rect 992 36660 998 36672
rect 1765 36669 1777 36672
rect 1811 36669 1823 36703
rect 1765 36663 1823 36669
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1581 35683 1639 35689
rect 1581 35649 1593 35683
rect 1627 35680 1639 35683
rect 11698 35680 11704 35692
rect 1627 35652 11704 35680
rect 1627 35649 1639 35652
rect 1581 35643 1639 35649
rect 11698 35640 11704 35652
rect 11756 35640 11762 35692
rect 934 35572 940 35624
rect 992 35612 998 35624
rect 1765 35615 1823 35621
rect 1765 35612 1777 35615
rect 992 35584 1777 35612
rect 992 35572 998 35584
rect 1765 35581 1777 35584
rect 1811 35581 1823 35615
rect 1765 35575 1823 35581
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1581 35071 1639 35077
rect 1581 35037 1593 35071
rect 1627 35068 1639 35071
rect 5534 35068 5540 35080
rect 1627 35040 5540 35068
rect 1627 35037 1639 35040
rect 1581 35031 1639 35037
rect 5534 35028 5540 35040
rect 5592 35028 5598 35080
rect 934 34960 940 35012
rect 992 35000 998 35012
rect 1857 35003 1915 35009
rect 1857 35000 1869 35003
rect 992 34972 1869 35000
rect 992 34960 998 34972
rect 1857 34969 1869 34972
rect 1903 34969 1915 35003
rect 1857 34963 1915 34969
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1857 34663 1915 34669
rect 1857 34629 1869 34663
rect 1903 34660 1915 34663
rect 4614 34660 4620 34672
rect 1903 34632 4620 34660
rect 1903 34629 1915 34632
rect 1857 34623 1915 34629
rect 4614 34620 4620 34632
rect 4672 34620 4678 34672
rect 1026 34552 1032 34604
rect 1084 34592 1090 34604
rect 1673 34595 1731 34601
rect 1673 34592 1685 34595
rect 1084 34564 1685 34592
rect 1084 34552 1090 34564
rect 1673 34561 1685 34564
rect 1719 34561 1731 34595
rect 1673 34555 1731 34561
rect 2409 34595 2467 34601
rect 2409 34561 2421 34595
rect 2455 34561 2467 34595
rect 2409 34555 2467 34561
rect 934 34484 940 34536
rect 992 34524 998 34536
rect 2424 34524 2452 34555
rect 992 34496 2452 34524
rect 2593 34527 2651 34533
rect 992 34484 998 34496
rect 2593 34493 2605 34527
rect 2639 34524 2651 34527
rect 2682 34524 2688 34536
rect 2639 34496 2688 34524
rect 2639 34493 2651 34496
rect 2593 34487 2651 34493
rect 2682 34484 2688 34496
rect 2740 34484 2746 34536
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1118 33872 1124 33924
rect 1176 33912 1182 33924
rect 1673 33915 1731 33921
rect 1673 33912 1685 33915
rect 1176 33884 1685 33912
rect 1176 33872 1182 33884
rect 1673 33881 1685 33884
rect 1719 33881 1731 33915
rect 1673 33875 1731 33881
rect 1857 33915 1915 33921
rect 1857 33881 1869 33915
rect 1903 33912 1915 33915
rect 2130 33912 2136 33924
rect 1903 33884 2136 33912
rect 1903 33881 1915 33884
rect 1857 33875 1915 33881
rect 2130 33872 2136 33884
rect 2188 33872 2194 33924
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1581 33507 1639 33513
rect 1581 33473 1593 33507
rect 1627 33504 1639 33507
rect 23750 33504 23756 33516
rect 1627 33476 23756 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 23750 33464 23756 33476
rect 23808 33464 23814 33516
rect 934 33396 940 33448
rect 992 33436 998 33448
rect 1765 33439 1823 33445
rect 1765 33436 1777 33439
rect 992 33408 1777 33436
rect 992 33396 998 33408
rect 1765 33405 1777 33408
rect 1811 33405 1823 33439
rect 1765 33399 1823 33405
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 934 32784 940 32836
rect 992 32824 998 32836
rect 1673 32827 1731 32833
rect 1673 32824 1685 32827
rect 992 32796 1685 32824
rect 992 32784 998 32796
rect 1673 32793 1685 32796
rect 1719 32793 1731 32827
rect 1673 32787 1731 32793
rect 1857 32827 1915 32833
rect 1857 32793 1869 32827
rect 1903 32824 1915 32827
rect 2498 32824 2504 32836
rect 1903 32796 2504 32824
rect 1903 32793 1915 32796
rect 1857 32787 1915 32793
rect 2498 32784 2504 32796
rect 2556 32784 2562 32836
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 5534 32444 5540 32496
rect 5592 32484 5598 32496
rect 22830 32484 22836 32496
rect 5592 32456 22836 32484
rect 5592 32444 5598 32456
rect 22830 32444 22836 32456
rect 22888 32444 22894 32496
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 12434 32416 12440 32428
rect 1627 32388 12440 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 12434 32376 12440 32388
rect 12492 32376 12498 32428
rect 934 32308 940 32360
rect 992 32348 998 32360
rect 1765 32351 1823 32357
rect 1765 32348 1777 32351
rect 992 32320 1777 32348
rect 992 32308 998 32320
rect 1765 32317 1777 32320
rect 1811 32317 1823 32351
rect 1765 32311 1823 32317
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1857 31943 1915 31949
rect 1857 31909 1869 31943
rect 1903 31940 1915 31943
rect 1903 31912 4016 31940
rect 1903 31909 1915 31912
rect 1857 31903 1915 31909
rect 1026 31832 1032 31884
rect 1084 31872 1090 31884
rect 3988 31872 4016 31912
rect 4062 31900 4068 31952
rect 4120 31940 4126 31952
rect 6178 31940 6184 31952
rect 4120 31912 6184 31940
rect 4120 31900 4126 31912
rect 6178 31900 6184 31912
rect 6236 31900 6242 31952
rect 6638 31872 6644 31884
rect 1084 31844 2452 31872
rect 3988 31844 6644 31872
rect 1084 31832 1090 31844
rect 934 31764 940 31816
rect 992 31804 998 31816
rect 2424 31813 2452 31844
rect 6638 31832 6644 31844
rect 6696 31832 6702 31884
rect 1673 31807 1731 31813
rect 1673 31804 1685 31807
rect 992 31776 1685 31804
rect 992 31764 998 31776
rect 1673 31773 1685 31776
rect 1719 31773 1731 31807
rect 1673 31767 1731 31773
rect 2409 31807 2467 31813
rect 2409 31773 2421 31807
rect 2455 31773 2467 31807
rect 2409 31767 2467 31773
rect 2590 31764 2596 31816
rect 2648 31764 2654 31816
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1581 31331 1639 31337
rect 1581 31297 1593 31331
rect 1627 31328 1639 31331
rect 26050 31328 26056 31340
rect 1627 31300 26056 31328
rect 1627 31297 1639 31300
rect 1581 31291 1639 31297
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 934 31220 940 31272
rect 992 31260 998 31272
rect 1765 31263 1823 31269
rect 1765 31260 1777 31263
rect 992 31232 1777 31260
rect 992 31220 998 31232
rect 1765 31229 1777 31232
rect 1811 31229 1823 31263
rect 1765 31223 1823 31229
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 934 30608 940 30660
rect 992 30648 998 30660
rect 1673 30651 1731 30657
rect 1673 30648 1685 30651
rect 992 30620 1685 30648
rect 992 30608 998 30620
rect 1673 30617 1685 30620
rect 1719 30617 1731 30651
rect 1673 30611 1731 30617
rect 1765 30583 1823 30589
rect 1765 30549 1777 30583
rect 1811 30580 1823 30583
rect 1854 30580 1860 30592
rect 1811 30552 1860 30580
rect 1811 30549 1823 30552
rect 1765 30543 1823 30549
rect 1854 30540 1860 30552
rect 1912 30540 1918 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 10410 30308 10416 30320
rect 1596 30280 10416 30308
rect 1596 30249 1624 30280
rect 10410 30268 10416 30280
rect 10468 30268 10474 30320
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30209 1639 30243
rect 1581 30203 1639 30209
rect 2593 30243 2651 30249
rect 2593 30209 2605 30243
rect 2639 30209 2651 30243
rect 2593 30203 2651 30209
rect 934 30132 940 30184
rect 992 30172 998 30184
rect 1765 30175 1823 30181
rect 1765 30172 1777 30175
rect 992 30144 1777 30172
rect 992 30132 998 30144
rect 1765 30141 1777 30144
rect 1811 30141 1823 30175
rect 1765 30135 1823 30141
rect 1026 30064 1032 30116
rect 1084 30104 1090 30116
rect 2608 30104 2636 30203
rect 1084 30076 2636 30104
rect 2777 30107 2835 30113
rect 1084 30064 1090 30076
rect 2777 30073 2789 30107
rect 2823 30104 2835 30107
rect 10778 30104 10784 30116
rect 2823 30076 10784 30104
rect 2823 30073 2835 30076
rect 2777 30067 2835 30073
rect 10778 30064 10784 30076
rect 10836 30064 10842 30116
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 12434 29588 12440 29640
rect 12492 29628 12498 29640
rect 25590 29628 25596 29640
rect 12492 29600 25596 29628
rect 12492 29588 12498 29600
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 934 29520 940 29572
rect 992 29560 998 29572
rect 1673 29563 1731 29569
rect 1673 29560 1685 29563
rect 992 29532 1685 29560
rect 992 29520 998 29532
rect 1673 29529 1685 29532
rect 1719 29529 1731 29563
rect 1673 29523 1731 29529
rect 2041 29563 2099 29569
rect 2041 29529 2053 29563
rect 2087 29560 2099 29563
rect 2406 29560 2412 29572
rect 2087 29532 2412 29560
rect 2087 29529 2099 29532
rect 2041 29523 2099 29529
rect 2406 29520 2412 29532
rect 2464 29520 2470 29572
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 13538 29220 13544 29232
rect 1596 29192 13544 29220
rect 1596 29161 1624 29192
rect 13538 29180 13544 29192
rect 13596 29180 13602 29232
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29121 1639 29155
rect 1581 29115 1639 29121
rect 2593 29155 2651 29161
rect 2593 29121 2605 29155
rect 2639 29121 2651 29155
rect 2593 29115 2651 29121
rect 1026 29044 1032 29096
rect 1084 29084 1090 29096
rect 1765 29087 1823 29093
rect 1765 29084 1777 29087
rect 1084 29056 1777 29084
rect 1084 29044 1090 29056
rect 1765 29053 1777 29056
rect 1811 29053 1823 29087
rect 1765 29047 1823 29053
rect 934 28976 940 29028
rect 992 29016 998 29028
rect 2608 29016 2636 29115
rect 992 28988 2636 29016
rect 2777 29019 2835 29025
rect 992 28976 998 28988
rect 2777 28985 2789 29019
rect 2823 29016 2835 29019
rect 6454 29016 6460 29028
rect 2823 28988 6460 29016
rect 2823 28985 2835 28988
rect 2777 28979 2835 28985
rect 6454 28976 6460 28988
rect 6512 28976 6518 29028
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 934 28432 940 28484
rect 992 28472 998 28484
rect 1673 28475 1731 28481
rect 1673 28472 1685 28475
rect 992 28444 1685 28472
rect 992 28432 998 28444
rect 1673 28441 1685 28444
rect 1719 28441 1731 28475
rect 1673 28435 1731 28441
rect 4614 28432 4620 28484
rect 4672 28472 4678 28484
rect 10686 28472 10692 28484
rect 4672 28444 10692 28472
rect 4672 28432 4678 28444
rect 10686 28432 10692 28444
rect 10744 28432 10750 28484
rect 1949 28407 2007 28413
rect 1949 28373 1961 28407
rect 1995 28404 2007 28407
rect 31938 28404 31944 28416
rect 1995 28376 31944 28404
rect 1995 28373 2007 28376
rect 1949 28367 2007 28373
rect 31938 28364 31944 28376
rect 31996 28364 32002 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 4062 28132 4068 28144
rect 1596 28104 4068 28132
rect 1596 28073 1624 28104
rect 4062 28092 4068 28104
rect 4120 28092 4126 28144
rect 1581 28067 1639 28073
rect 1581 28033 1593 28067
rect 1627 28033 1639 28067
rect 2593 28067 2651 28073
rect 2593 28064 2605 28067
rect 1581 28027 1639 28033
rect 1688 28036 2605 28064
rect 934 27956 940 28008
rect 992 27996 998 28008
rect 1688 27996 1716 28036
rect 2593 28033 2605 28036
rect 2639 28033 2651 28067
rect 2593 28027 2651 28033
rect 992 27968 1716 27996
rect 1765 27999 1823 28005
rect 992 27956 998 27968
rect 1765 27965 1777 27999
rect 1811 27965 1823 27999
rect 1765 27959 1823 27965
rect 1026 27888 1032 27940
rect 1084 27928 1090 27940
rect 1780 27928 1808 27959
rect 1084 27900 1808 27928
rect 2777 27931 2835 27937
rect 1084 27888 1090 27900
rect 2777 27897 2789 27931
rect 2823 27928 2835 27931
rect 4614 27928 4620 27940
rect 2823 27900 4620 27928
rect 2823 27897 2835 27900
rect 2777 27891 2835 27897
rect 4614 27888 4620 27900
rect 4672 27888 4678 27940
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 10318 27548 10324 27600
rect 10376 27588 10382 27600
rect 11238 27588 11244 27600
rect 10376 27560 11244 27588
rect 10376 27548 10382 27560
rect 11238 27548 11244 27560
rect 11296 27548 11302 27600
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19981 27455 20039 27461
rect 19981 27421 19993 27455
rect 20027 27452 20039 27455
rect 20622 27452 20628 27464
rect 20027 27424 20628 27452
rect 20027 27421 20039 27424
rect 19981 27415 20039 27421
rect 934 27344 940 27396
rect 992 27384 998 27396
rect 1673 27387 1731 27393
rect 1673 27384 1685 27387
rect 992 27356 1685 27384
rect 992 27344 998 27356
rect 1673 27353 1685 27356
rect 1719 27353 1731 27387
rect 19812 27384 19840 27415
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 19812 27356 20024 27384
rect 1673 27347 1731 27353
rect 19996 27328 20024 27356
rect 1946 27276 1952 27328
rect 2004 27276 2010 27328
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19889 27319 19947 27325
rect 19889 27316 19901 27319
rect 19116 27288 19901 27316
rect 19116 27276 19122 27288
rect 19889 27285 19901 27288
rect 19935 27285 19947 27319
rect 19889 27279 19947 27285
rect 19978 27276 19984 27328
rect 20036 27276 20042 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1946 27072 1952 27124
rect 2004 27112 2010 27124
rect 19334 27112 19340 27124
rect 2004 27084 19340 27112
rect 2004 27072 2010 27084
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 19797 27115 19855 27121
rect 19797 27081 19809 27115
rect 19843 27112 19855 27115
rect 19978 27112 19984 27124
rect 19843 27084 19984 27112
rect 19843 27081 19855 27084
rect 19797 27075 19855 27081
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 20622 27072 20628 27124
rect 20680 27072 20686 27124
rect 1026 27004 1032 27056
rect 1084 27044 1090 27056
rect 2593 27047 2651 27053
rect 2593 27044 2605 27047
rect 1084 27016 2605 27044
rect 1084 27004 1090 27016
rect 2593 27013 2605 27016
rect 2639 27013 2651 27047
rect 2593 27007 2651 27013
rect 5258 27004 5264 27056
rect 5316 27044 5322 27056
rect 33778 27044 33784 27056
rect 5316 27016 33784 27044
rect 5316 27004 5322 27016
rect 33778 27004 33784 27016
rect 33836 27004 33842 27056
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26976 1639 26979
rect 3970 26976 3976 26988
rect 1627 26948 3976 26976
rect 1627 26945 1639 26948
rect 1581 26939 1639 26945
rect 3970 26936 3976 26948
rect 4028 26936 4034 26988
rect 14642 26936 14648 26988
rect 14700 26936 14706 26988
rect 15381 26979 15439 26985
rect 15381 26976 15393 26979
rect 14844 26948 15393 26976
rect 1118 26868 1124 26920
rect 1176 26908 1182 26920
rect 1765 26911 1823 26917
rect 1765 26908 1777 26911
rect 1176 26880 1777 26908
rect 1176 26868 1182 26880
rect 1765 26877 1777 26880
rect 1811 26877 1823 26911
rect 1765 26871 1823 26877
rect 4062 26868 4068 26920
rect 4120 26908 4126 26920
rect 14090 26908 14096 26920
rect 4120 26880 14096 26908
rect 4120 26868 4126 26880
rect 14090 26868 14096 26880
rect 14148 26868 14154 26920
rect 2774 26800 2780 26852
rect 2832 26800 2838 26852
rect 14844 26849 14872 26948
rect 15381 26945 15393 26948
rect 15427 26945 15439 26979
rect 15381 26939 15439 26945
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 15930 26976 15936 26988
rect 15611 26948 15936 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 20346 26976 20352 26988
rect 19628 26948 20352 26976
rect 14918 26868 14924 26920
rect 14976 26868 14982 26920
rect 15948 26908 15976 26936
rect 19628 26917 19656 26948
rect 20346 26936 20352 26948
rect 20404 26976 20410 26988
rect 20441 26979 20499 26985
rect 20441 26976 20453 26979
rect 20404 26948 20453 26976
rect 20404 26936 20410 26948
rect 20441 26945 20453 26948
rect 20487 26945 20499 26979
rect 20441 26939 20499 26945
rect 24305 26979 24363 26985
rect 24305 26945 24317 26979
rect 24351 26976 24363 26979
rect 24946 26976 24952 26988
rect 24351 26948 24952 26976
rect 24351 26945 24363 26948
rect 24305 26939 24363 26945
rect 24946 26936 24952 26948
rect 25004 26936 25010 26988
rect 34606 26936 34612 26988
rect 34664 26936 34670 26988
rect 19613 26911 19671 26917
rect 19613 26908 19625 26911
rect 15948 26880 19625 26908
rect 19613 26877 19625 26880
rect 19659 26877 19671 26911
rect 19613 26871 19671 26877
rect 19794 26868 19800 26920
rect 19852 26868 19858 26920
rect 20257 26911 20315 26917
rect 20257 26877 20269 26911
rect 20303 26908 20315 26911
rect 24581 26911 24639 26917
rect 24581 26908 24593 26911
rect 20303 26880 20484 26908
rect 20303 26877 20315 26880
rect 20257 26871 20315 26877
rect 20456 26852 20484 26880
rect 20548 26880 24593 26908
rect 14829 26843 14887 26849
rect 14829 26809 14841 26843
rect 14875 26809 14887 26843
rect 14829 26803 14887 26809
rect 19518 26800 19524 26852
rect 19576 26840 19582 26852
rect 20438 26840 20444 26852
rect 19576 26812 20444 26840
rect 19576 26800 19582 26812
rect 20438 26800 20444 26812
rect 20496 26800 20502 26852
rect 20548 26784 20576 26880
rect 24581 26877 24593 26880
rect 24627 26877 24639 26911
rect 24581 26871 24639 26877
rect 34146 26868 34152 26920
rect 34204 26908 34210 26920
rect 34885 26911 34943 26917
rect 34885 26908 34897 26911
rect 34204 26880 34897 26908
rect 34204 26868 34210 26880
rect 34885 26877 34897 26880
rect 34931 26908 34943 26911
rect 36354 26908 36360 26920
rect 34931 26880 36360 26908
rect 34931 26877 34943 26880
rect 34885 26871 34943 26877
rect 36354 26868 36360 26880
rect 36412 26868 36418 26920
rect 14734 26732 14740 26784
rect 14792 26732 14798 26784
rect 15378 26732 15384 26784
rect 15436 26732 15442 26784
rect 19794 26732 19800 26784
rect 19852 26772 19858 26784
rect 20530 26772 20536 26784
rect 19852 26744 20536 26772
rect 19852 26732 19858 26744
rect 20530 26732 20536 26744
rect 20588 26732 20594 26784
rect 20622 26732 20628 26784
rect 20680 26772 20686 26784
rect 22002 26772 22008 26784
rect 20680 26744 22008 26772
rect 20680 26732 20686 26744
rect 22002 26732 22008 26744
rect 22060 26772 22066 26784
rect 24394 26772 24400 26784
rect 22060 26744 24400 26772
rect 22060 26732 22066 26744
rect 24394 26732 24400 26744
rect 24452 26732 24458 26784
rect 24489 26775 24547 26781
rect 24489 26741 24501 26775
rect 24535 26772 24547 26775
rect 24578 26772 24584 26784
rect 24535 26744 24584 26772
rect 24535 26741 24547 26744
rect 24489 26735 24547 26741
rect 24578 26732 24584 26744
rect 24636 26732 24642 26784
rect 34422 26732 34428 26784
rect 34480 26732 34486 26784
rect 34790 26732 34796 26784
rect 34848 26732 34854 26784
rect 35802 26732 35808 26784
rect 35860 26772 35866 26784
rect 38010 26772 38016 26784
rect 35860 26744 38016 26772
rect 35860 26732 35866 26744
rect 38010 26732 38016 26744
rect 38068 26732 38074 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1949 26571 2007 26577
rect 1949 26537 1961 26571
rect 1995 26568 2007 26571
rect 5258 26568 5264 26580
rect 1995 26540 5264 26568
rect 1995 26537 2007 26540
rect 1949 26531 2007 26537
rect 5258 26528 5264 26540
rect 5316 26528 5322 26580
rect 14826 26528 14832 26580
rect 14884 26568 14890 26580
rect 15749 26571 15807 26577
rect 15749 26568 15761 26571
rect 14884 26540 15761 26568
rect 14884 26528 14890 26540
rect 15749 26537 15761 26540
rect 15795 26537 15807 26571
rect 15749 26531 15807 26537
rect 15930 26528 15936 26580
rect 15988 26528 15994 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 21361 26571 21419 26577
rect 21361 26568 21373 26571
rect 20128 26540 21373 26568
rect 20128 26528 20134 26540
rect 21361 26537 21373 26540
rect 21407 26568 21419 26571
rect 22097 26571 22155 26577
rect 22097 26568 22109 26571
rect 21407 26540 22109 26568
rect 21407 26537 21419 26540
rect 21361 26531 21419 26537
rect 22097 26537 22109 26540
rect 22143 26537 22155 26571
rect 22097 26531 22155 26537
rect 37826 26528 37832 26580
rect 37884 26568 37890 26580
rect 37884 26540 39344 26568
rect 37884 26528 37890 26540
rect 14734 26460 14740 26512
rect 14792 26460 14798 26512
rect 20622 26460 20628 26512
rect 20680 26500 20686 26512
rect 24581 26503 24639 26509
rect 20680 26472 22324 26500
rect 20680 26460 20686 26472
rect 2498 26392 2504 26444
rect 2556 26432 2562 26444
rect 2961 26435 3019 26441
rect 2961 26432 2973 26435
rect 2556 26404 2973 26432
rect 2556 26392 2562 26404
rect 2961 26401 2973 26404
rect 3007 26401 3019 26435
rect 2961 26395 3019 26401
rect 3145 26435 3203 26441
rect 3145 26401 3157 26435
rect 3191 26432 3203 26435
rect 4338 26432 4344 26444
rect 3191 26404 4344 26432
rect 3191 26401 3203 26404
rect 3145 26395 3203 26401
rect 4338 26392 4344 26404
rect 4396 26392 4402 26444
rect 6454 26392 6460 26444
rect 6512 26392 6518 26444
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26432 6607 26435
rect 8018 26432 8024 26444
rect 6595 26404 8024 26432
rect 6595 26401 6607 26404
rect 6549 26395 6607 26401
rect 4356 26364 4384 26392
rect 6564 26364 6592 26395
rect 8018 26392 8024 26404
rect 8076 26392 8082 26444
rect 14752 26432 14780 26460
rect 15105 26435 15163 26441
rect 15105 26432 15117 26435
rect 13740 26404 15117 26432
rect 4356 26336 6592 26364
rect 6638 26324 6644 26376
rect 6696 26364 6702 26376
rect 13740 26373 13768 26404
rect 15105 26401 15117 26404
rect 15151 26401 15163 26435
rect 15105 26395 15163 26401
rect 20165 26435 20223 26441
rect 20165 26401 20177 26435
rect 20211 26432 20223 26435
rect 20211 26404 21312 26432
rect 20211 26401 20223 26404
rect 20165 26395 20223 26401
rect 7929 26367 7987 26373
rect 7929 26364 7941 26367
rect 6696 26336 7941 26364
rect 6696 26324 6702 26336
rect 7929 26333 7941 26336
rect 7975 26333 7987 26367
rect 7929 26327 7987 26333
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13725 26367 13783 26373
rect 13725 26333 13737 26367
rect 13771 26333 13783 26367
rect 13725 26327 13783 26333
rect 934 26256 940 26308
rect 992 26296 998 26308
rect 1673 26299 1731 26305
rect 1673 26296 1685 26299
rect 992 26268 1685 26296
rect 992 26256 998 26268
rect 1673 26265 1685 26268
rect 1719 26265 1731 26299
rect 1673 26259 1731 26265
rect 7650 26256 7656 26308
rect 7708 26296 7714 26308
rect 7837 26299 7895 26305
rect 7837 26296 7849 26299
rect 7708 26268 7849 26296
rect 7708 26256 7714 26268
rect 7837 26265 7849 26268
rect 7883 26265 7895 26299
rect 7837 26259 7895 26265
rect 2314 26188 2320 26240
rect 2372 26228 2378 26240
rect 2501 26231 2559 26237
rect 2501 26228 2513 26231
rect 2372 26200 2513 26228
rect 2372 26188 2378 26200
rect 2501 26197 2513 26200
rect 2547 26197 2559 26231
rect 2501 26191 2559 26197
rect 2869 26231 2927 26237
rect 2869 26197 2881 26231
rect 2915 26228 2927 26231
rect 3418 26228 3424 26240
rect 2915 26200 3424 26228
rect 2915 26197 2927 26200
rect 2869 26191 2927 26197
rect 3418 26188 3424 26200
rect 3476 26188 3482 26240
rect 5994 26188 6000 26240
rect 6052 26188 6058 26240
rect 6362 26188 6368 26240
rect 6420 26188 6426 26240
rect 7466 26188 7472 26240
rect 7524 26188 7530 26240
rect 13556 26228 13584 26327
rect 14734 26324 14740 26376
rect 14792 26324 14798 26376
rect 14921 26367 14979 26373
rect 14921 26333 14933 26367
rect 14967 26364 14979 26367
rect 15010 26364 15016 26376
rect 14967 26336 15016 26364
rect 14967 26333 14979 26336
rect 14921 26327 14979 26333
rect 15010 26324 15016 26336
rect 15068 26364 15074 26376
rect 15068 26336 15700 26364
rect 15068 26324 15074 26336
rect 15672 26308 15700 26336
rect 20346 26324 20352 26376
rect 20404 26324 20410 26376
rect 20438 26324 20444 26376
rect 20496 26324 20502 26376
rect 20533 26367 20591 26373
rect 20533 26333 20545 26367
rect 20579 26333 20591 26367
rect 20533 26327 20591 26333
rect 13630 26256 13636 26308
rect 13688 26256 13694 26308
rect 14642 26256 14648 26308
rect 14700 26296 14706 26308
rect 15565 26299 15623 26305
rect 15565 26296 15577 26299
rect 14700 26268 15577 26296
rect 14700 26256 14706 26268
rect 15565 26265 15577 26268
rect 15611 26265 15623 26299
rect 15565 26259 15623 26265
rect 15102 26228 15108 26240
rect 13556 26200 15108 26228
rect 15102 26188 15108 26200
rect 15160 26188 15166 26240
rect 15580 26228 15608 26259
rect 15654 26256 15660 26308
rect 15712 26296 15718 26308
rect 15749 26299 15807 26305
rect 15749 26296 15761 26299
rect 15712 26268 15761 26296
rect 15712 26256 15718 26268
rect 15749 26265 15761 26268
rect 15795 26265 15807 26299
rect 15749 26259 15807 26265
rect 19242 26256 19248 26308
rect 19300 26296 19306 26308
rect 20548 26296 20576 26327
rect 20622 26324 20628 26376
rect 20680 26324 20686 26376
rect 20714 26324 20720 26376
rect 20772 26364 20778 26376
rect 20772 26336 21220 26364
rect 20772 26324 20778 26336
rect 21192 26305 21220 26336
rect 21177 26299 21235 26305
rect 19300 26268 21128 26296
rect 19300 26256 19306 26268
rect 15838 26228 15844 26240
rect 15580 26200 15844 26228
rect 15838 26188 15844 26200
rect 15896 26188 15902 26240
rect 21100 26228 21128 26268
rect 21177 26265 21189 26299
rect 21223 26265 21235 26299
rect 21284 26296 21312 26404
rect 22296 26376 22324 26472
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 24854 26500 24860 26512
rect 24627 26472 24860 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 24854 26460 24860 26472
rect 24912 26460 24918 26512
rect 33502 26460 33508 26512
rect 33560 26500 33566 26512
rect 37737 26503 37795 26509
rect 33560 26472 35940 26500
rect 33560 26460 33566 26472
rect 24394 26392 24400 26444
rect 24452 26432 24458 26444
rect 24452 26404 24900 26432
rect 24452 26392 24458 26404
rect 22002 26324 22008 26376
rect 22060 26324 22066 26376
rect 22278 26324 22284 26376
rect 22336 26324 22342 26376
rect 24578 26324 24584 26376
rect 24636 26324 24642 26376
rect 24872 26373 24900 26404
rect 28258 26392 28264 26444
rect 28316 26432 28322 26444
rect 28718 26432 28724 26444
rect 28316 26404 28724 26432
rect 28316 26392 28322 26404
rect 28718 26392 28724 26404
rect 28776 26432 28782 26444
rect 28776 26404 32260 26432
rect 28776 26392 28782 26404
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26333 24915 26367
rect 24857 26327 24915 26333
rect 31941 26367 31999 26373
rect 31941 26333 31953 26367
rect 31987 26364 31999 26367
rect 32122 26364 32128 26376
rect 31987 26336 32128 26364
rect 31987 26333 31999 26336
rect 31941 26327 31999 26333
rect 32122 26324 32128 26336
rect 32180 26324 32186 26376
rect 21377 26299 21435 26305
rect 21377 26296 21389 26299
rect 21284 26268 21389 26296
rect 21177 26259 21235 26265
rect 21377 26265 21389 26268
rect 21423 26265 21435 26299
rect 22189 26299 22247 26305
rect 22189 26296 22201 26299
rect 21377 26259 21435 26265
rect 21468 26268 21956 26296
rect 21468 26228 21496 26268
rect 21100 26200 21496 26228
rect 21542 26188 21548 26240
rect 21600 26188 21606 26240
rect 21928 26228 21956 26268
rect 22066 26268 22201 26296
rect 22066 26228 22094 26268
rect 22189 26265 22201 26268
rect 22235 26296 22247 26299
rect 24765 26299 24823 26305
rect 24765 26296 24777 26299
rect 22235 26268 24777 26296
rect 22235 26265 22247 26268
rect 22189 26259 22247 26265
rect 24765 26265 24777 26268
rect 24811 26296 24823 26299
rect 24946 26296 24952 26308
rect 24811 26268 24952 26296
rect 24811 26265 24823 26268
rect 24765 26259 24823 26265
rect 24946 26256 24952 26268
rect 25004 26296 25010 26308
rect 25958 26296 25964 26308
rect 25004 26268 25964 26296
rect 25004 26256 25010 26268
rect 25958 26256 25964 26268
rect 26016 26256 26022 26308
rect 32232 26296 32260 26404
rect 32490 26392 32496 26444
rect 32548 26432 32554 26444
rect 35912 26441 35940 26472
rect 37737 26469 37749 26503
rect 37783 26500 37795 26503
rect 39316 26500 39344 26540
rect 40310 26500 40316 26512
rect 37783 26472 38516 26500
rect 37783 26469 37795 26472
rect 37737 26463 37795 26469
rect 38488 26441 38516 26472
rect 39316 26472 40316 26500
rect 33597 26435 33655 26441
rect 33597 26432 33609 26435
rect 32548 26404 33609 26432
rect 32548 26392 32554 26404
rect 33597 26401 33609 26404
rect 33643 26401 33655 26435
rect 33597 26395 33655 26401
rect 34241 26435 34299 26441
rect 34241 26401 34253 26435
rect 34287 26432 34299 26435
rect 35345 26435 35403 26441
rect 35345 26432 35357 26435
rect 34287 26404 35357 26432
rect 34287 26401 34299 26404
rect 34241 26395 34299 26401
rect 35345 26401 35357 26404
rect 35391 26401 35403 26435
rect 35345 26395 35403 26401
rect 35897 26435 35955 26441
rect 35897 26401 35909 26435
rect 35943 26432 35955 26435
rect 38473 26435 38531 26441
rect 35943 26404 38148 26432
rect 35943 26401 35955 26404
rect 35897 26395 35955 26401
rect 32306 26324 32312 26376
rect 32364 26324 32370 26376
rect 34146 26324 34152 26376
rect 34204 26324 34210 26376
rect 34422 26324 34428 26376
rect 34480 26364 34486 26376
rect 35069 26367 35127 26373
rect 35069 26364 35081 26367
rect 34480 26336 35081 26364
rect 34480 26324 34486 26336
rect 35069 26333 35081 26336
rect 35115 26333 35127 26367
rect 35069 26327 35127 26333
rect 35250 26324 35256 26376
rect 35308 26324 35314 26376
rect 36265 26367 36323 26373
rect 36265 26333 36277 26367
rect 36311 26364 36323 26367
rect 37642 26364 37648 26376
rect 36311 26336 37648 26364
rect 36311 26333 36323 26336
rect 36265 26327 36323 26333
rect 37642 26324 37648 26336
rect 37700 26324 37706 26376
rect 37737 26367 37795 26373
rect 37737 26333 37749 26367
rect 37783 26364 37795 26367
rect 37826 26364 37832 26376
rect 37783 26336 37832 26364
rect 37783 26333 37795 26336
rect 37737 26327 37795 26333
rect 37826 26324 37832 26336
rect 37884 26324 37890 26376
rect 38010 26324 38016 26376
rect 38068 26324 38074 26376
rect 38120 26364 38148 26404
rect 38473 26401 38485 26435
rect 38519 26401 38531 26435
rect 38473 26395 38531 26401
rect 38657 26435 38715 26441
rect 38657 26401 38669 26435
rect 38703 26432 38715 26435
rect 38838 26432 38844 26444
rect 38703 26404 38844 26432
rect 38703 26401 38715 26404
rect 38657 26395 38715 26401
rect 38838 26392 38844 26404
rect 38896 26432 38902 26444
rect 39206 26432 39212 26444
rect 38896 26404 39212 26432
rect 38896 26392 38902 26404
rect 39206 26392 39212 26404
rect 39264 26392 39270 26444
rect 39316 26373 39344 26472
rect 40310 26460 40316 26472
rect 40368 26460 40374 26512
rect 39390 26392 39396 26444
rect 39448 26432 39454 26444
rect 39448 26404 40632 26432
rect 39448 26392 39454 26404
rect 38565 26367 38623 26373
rect 38565 26364 38577 26367
rect 38120 26336 38577 26364
rect 38565 26333 38577 26336
rect 38611 26333 38623 26367
rect 38565 26327 38623 26333
rect 39025 26367 39083 26373
rect 39025 26333 39037 26367
rect 39071 26333 39083 26367
rect 39025 26327 39083 26333
rect 39301 26367 39359 26373
rect 39301 26333 39313 26367
rect 39347 26333 39359 26367
rect 39301 26327 39359 26333
rect 32674 26296 32680 26308
rect 32232 26268 32680 26296
rect 32674 26256 32680 26268
rect 32732 26256 32738 26308
rect 33137 26299 33195 26305
rect 33137 26265 33149 26299
rect 33183 26296 33195 26299
rect 33686 26296 33692 26308
rect 33183 26268 33692 26296
rect 33183 26265 33195 26268
rect 33137 26259 33195 26265
rect 33686 26256 33692 26268
rect 33744 26256 33750 26308
rect 34790 26256 34796 26308
rect 34848 26296 34854 26308
rect 34885 26299 34943 26305
rect 34885 26296 34897 26299
rect 34848 26268 34897 26296
rect 34848 26256 34854 26268
rect 34885 26265 34897 26268
rect 34931 26265 34943 26299
rect 34885 26259 34943 26265
rect 34974 26256 34980 26308
rect 35032 26296 35038 26308
rect 36173 26299 36231 26305
rect 36173 26296 36185 26299
rect 35032 26268 36185 26296
rect 35032 26256 35038 26268
rect 36173 26265 36185 26268
rect 36219 26265 36231 26299
rect 36173 26259 36231 26265
rect 36354 26256 36360 26308
rect 36412 26305 36418 26308
rect 36412 26299 36440 26305
rect 36428 26265 36440 26299
rect 39040 26296 39068 26327
rect 40034 26324 40040 26376
rect 40092 26324 40098 26376
rect 40218 26324 40224 26376
rect 40276 26324 40282 26376
rect 40313 26367 40371 26373
rect 40313 26333 40325 26367
rect 40359 26333 40371 26367
rect 40313 26327 40371 26333
rect 40126 26296 40132 26308
rect 36412 26259 36440 26265
rect 38028 26268 40132 26296
rect 36412 26256 36418 26259
rect 21928 26200 22094 26228
rect 36538 26188 36544 26240
rect 36596 26188 36602 26240
rect 37921 26231 37979 26237
rect 37921 26197 37933 26231
rect 37967 26228 37979 26231
rect 38028 26228 38056 26268
rect 40126 26256 40132 26268
rect 40184 26256 40190 26308
rect 37967 26200 38056 26228
rect 37967 26197 37979 26200
rect 37921 26191 37979 26197
rect 38746 26188 38752 26240
rect 38804 26228 38810 26240
rect 40034 26228 40040 26240
rect 38804 26200 40040 26228
rect 38804 26188 38810 26200
rect 40034 26188 40040 26200
rect 40092 26228 40098 26240
rect 40328 26228 40356 26327
rect 40402 26324 40408 26376
rect 40460 26324 40466 26376
rect 40604 26373 40632 26404
rect 40589 26367 40647 26373
rect 40589 26333 40601 26367
rect 40635 26333 40647 26367
rect 40589 26327 40647 26333
rect 40773 26299 40831 26305
rect 40773 26265 40785 26299
rect 40819 26296 40831 26299
rect 40862 26296 40868 26308
rect 40819 26268 40868 26296
rect 40819 26265 40831 26268
rect 40773 26259 40831 26265
rect 40862 26256 40868 26268
rect 40920 26256 40926 26308
rect 40092 26200 40356 26228
rect 40092 26188 40098 26200
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 4249 26027 4307 26033
rect 4249 25993 4261 26027
rect 4295 26024 4307 26027
rect 4614 26024 4620 26036
rect 4295 25996 4620 26024
rect 4295 25993 4307 25996
rect 4249 25987 4307 25993
rect 4614 25984 4620 25996
rect 4672 25984 4678 26036
rect 8018 25984 8024 26036
rect 8076 25984 8082 26036
rect 10686 25984 10692 26036
rect 10744 25984 10750 26036
rect 15102 25984 15108 26036
rect 15160 25984 15166 26036
rect 17957 26027 18015 26033
rect 17957 25993 17969 26027
rect 18003 26024 18015 26027
rect 20438 26024 20444 26036
rect 18003 25996 20444 26024
rect 18003 25993 18015 25996
rect 17957 25987 18015 25993
rect 20438 25984 20444 25996
rect 20496 25984 20502 26036
rect 34882 25984 34888 26036
rect 34940 26024 34946 26036
rect 35069 26027 35127 26033
rect 35069 26024 35081 26027
rect 34940 25996 35081 26024
rect 34940 25984 34946 25996
rect 35069 25993 35081 25996
rect 35115 25993 35127 26027
rect 35069 25987 35127 25993
rect 36538 25984 36544 26036
rect 36596 26024 36602 26036
rect 36596 25996 39896 26024
rect 36596 25984 36602 25996
rect 1118 25916 1124 25968
rect 1176 25956 1182 25968
rect 2593 25959 2651 25965
rect 2593 25956 2605 25959
rect 1176 25928 2605 25956
rect 1176 25916 1182 25928
rect 2593 25925 2605 25928
rect 2639 25925 2651 25959
rect 2593 25919 2651 25925
rect 17773 25959 17831 25965
rect 17773 25925 17785 25959
rect 17819 25956 17831 25959
rect 19242 25956 19248 25968
rect 17819 25928 19248 25956
rect 17819 25925 17831 25928
rect 17773 25919 17831 25925
rect 19242 25916 19248 25928
rect 19300 25916 19306 25968
rect 30282 25956 30288 25968
rect 29840 25928 30288 25956
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 4157 25891 4215 25897
rect 1627 25860 4108 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 1026 25780 1032 25832
rect 1084 25820 1090 25832
rect 1765 25823 1823 25829
rect 1765 25820 1777 25823
rect 1084 25792 1777 25820
rect 1084 25780 1090 25792
rect 1765 25789 1777 25792
rect 1811 25789 1823 25823
rect 1765 25783 1823 25789
rect 2777 25755 2835 25761
rect 2777 25721 2789 25755
rect 2823 25752 2835 25755
rect 4080 25752 4108 25860
rect 4157 25857 4169 25891
rect 4203 25888 4215 25891
rect 4982 25888 4988 25900
rect 4203 25860 4988 25888
rect 4203 25857 4215 25860
rect 4157 25851 4215 25857
rect 4982 25848 4988 25860
rect 5040 25848 5046 25900
rect 7374 25848 7380 25900
rect 7432 25888 7438 25900
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 7432 25860 7941 25888
rect 7432 25848 7438 25860
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25888 10655 25891
rect 10686 25888 10692 25900
rect 10643 25860 10692 25888
rect 10643 25857 10655 25860
rect 10597 25851 10655 25857
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 14734 25848 14740 25900
rect 14792 25888 14798 25900
rect 14829 25891 14887 25897
rect 14829 25888 14841 25891
rect 14792 25860 14841 25888
rect 14792 25848 14798 25860
rect 14829 25857 14841 25860
rect 14875 25857 14887 25891
rect 14829 25851 14887 25857
rect 15838 25848 15844 25900
rect 15896 25888 15902 25900
rect 29840 25897 29868 25928
rect 30282 25916 30288 25928
rect 30340 25956 30346 25968
rect 32677 25959 32735 25965
rect 32677 25956 32689 25959
rect 30340 25928 32689 25956
rect 30340 25916 30346 25928
rect 32677 25925 32689 25928
rect 32723 25925 32735 25959
rect 37366 25956 37372 25968
rect 32677 25919 32735 25925
rect 33704 25928 37372 25956
rect 33704 25900 33732 25928
rect 18049 25891 18107 25897
rect 18049 25888 18061 25891
rect 15896 25860 18061 25888
rect 15896 25848 15902 25860
rect 18049 25857 18061 25860
rect 18095 25857 18107 25891
rect 18049 25851 18107 25857
rect 18141 25891 18199 25897
rect 18141 25857 18153 25891
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 29825 25891 29883 25897
rect 29825 25857 29837 25891
rect 29871 25857 29883 25891
rect 29825 25851 29883 25857
rect 29917 25891 29975 25897
rect 29917 25857 29929 25891
rect 29963 25857 29975 25891
rect 29917 25851 29975 25857
rect 4338 25780 4344 25832
rect 4396 25780 4402 25832
rect 8018 25780 8024 25832
rect 8076 25820 8082 25832
rect 10781 25823 10839 25829
rect 10781 25820 10793 25823
rect 8076 25792 10793 25820
rect 8076 25780 8082 25792
rect 10781 25789 10793 25792
rect 10827 25820 10839 25823
rect 10870 25820 10876 25832
rect 10827 25792 10876 25820
rect 10827 25789 10839 25792
rect 10781 25783 10839 25789
rect 10870 25780 10876 25792
rect 10928 25780 10934 25832
rect 14918 25780 14924 25832
rect 14976 25820 14982 25832
rect 15105 25823 15163 25829
rect 15105 25820 15117 25823
rect 14976 25792 15117 25820
rect 14976 25780 14982 25792
rect 15105 25789 15117 25792
rect 15151 25820 15163 25823
rect 15930 25820 15936 25832
rect 15151 25792 15936 25820
rect 15151 25789 15163 25792
rect 15105 25783 15163 25789
rect 15930 25780 15936 25792
rect 15988 25780 15994 25832
rect 17770 25780 17776 25832
rect 17828 25820 17834 25832
rect 18156 25820 18184 25851
rect 17828 25792 18184 25820
rect 17828 25780 17834 25792
rect 28994 25780 29000 25832
rect 29052 25820 29058 25832
rect 29932 25820 29960 25851
rect 30098 25848 30104 25900
rect 30156 25848 30162 25900
rect 30190 25848 30196 25900
rect 30248 25888 30254 25900
rect 30248 25860 31754 25888
rect 30248 25848 30254 25860
rect 29052 25792 29960 25820
rect 29052 25780 29058 25792
rect 4614 25752 4620 25764
rect 2823 25724 4016 25752
rect 4080 25724 4620 25752
rect 2823 25721 2835 25724
rect 2777 25715 2835 25721
rect 3789 25687 3847 25693
rect 3789 25653 3801 25687
rect 3835 25684 3847 25687
rect 3878 25684 3884 25696
rect 3835 25656 3884 25684
rect 3835 25653 3847 25656
rect 3789 25647 3847 25653
rect 3878 25644 3884 25656
rect 3936 25644 3942 25696
rect 3988 25684 4016 25724
rect 4614 25712 4620 25724
rect 4672 25712 4678 25764
rect 19334 25712 19340 25764
rect 19392 25752 19398 25764
rect 30834 25752 30840 25764
rect 19392 25724 30840 25752
rect 19392 25712 19398 25724
rect 30834 25712 30840 25724
rect 30892 25712 30898 25764
rect 31726 25752 31754 25860
rect 32122 25848 32128 25900
rect 32180 25888 32186 25900
rect 32309 25891 32367 25897
rect 32309 25888 32321 25891
rect 32180 25860 32321 25888
rect 32180 25848 32186 25860
rect 32309 25857 32321 25860
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 32490 25848 32496 25900
rect 32548 25848 32554 25900
rect 33502 25848 33508 25900
rect 33560 25888 33566 25900
rect 33597 25891 33655 25897
rect 33597 25888 33609 25891
rect 33560 25860 33609 25888
rect 33560 25848 33566 25860
rect 33597 25857 33609 25860
rect 33643 25857 33655 25891
rect 33597 25851 33655 25857
rect 33686 25848 33692 25900
rect 33744 25848 33750 25900
rect 35176 25897 35204 25928
rect 37366 25916 37372 25928
rect 37424 25916 37430 25968
rect 38838 25916 38844 25968
rect 38896 25916 38902 25968
rect 39868 25965 39896 25996
rect 40126 25984 40132 26036
rect 40184 26024 40190 26036
rect 41417 26027 41475 26033
rect 41417 26024 41429 26027
rect 40184 25996 41429 26024
rect 40184 25984 40190 25996
rect 41417 25993 41429 25996
rect 41463 26024 41475 26027
rect 42705 26027 42763 26033
rect 42705 26024 42717 26027
rect 41463 25996 42717 26024
rect 41463 25993 41475 25996
rect 41417 25987 41475 25993
rect 42705 25993 42717 25996
rect 42751 25993 42763 26027
rect 42705 25987 42763 25993
rect 39853 25959 39911 25965
rect 39853 25925 39865 25959
rect 39899 25956 39911 25959
rect 40218 25956 40224 25968
rect 39899 25928 40224 25956
rect 39899 25925 39911 25928
rect 39853 25919 39911 25925
rect 40218 25916 40224 25928
rect 40276 25916 40282 25968
rect 34977 25891 35035 25897
rect 34977 25857 34989 25891
rect 35023 25857 35035 25891
rect 34977 25851 35035 25857
rect 35161 25891 35219 25897
rect 35161 25857 35173 25891
rect 35207 25857 35219 25891
rect 35161 25851 35219 25857
rect 34992 25820 35020 25851
rect 35250 25848 35256 25900
rect 35308 25888 35314 25900
rect 35989 25891 36047 25897
rect 35989 25888 36001 25891
rect 35308 25860 36001 25888
rect 35308 25848 35314 25860
rect 35989 25857 36001 25860
rect 36035 25888 36047 25891
rect 36035 25860 36124 25888
rect 36035 25857 36047 25860
rect 35989 25851 36047 25857
rect 35894 25820 35900 25832
rect 33888 25792 35900 25820
rect 33888 25752 33916 25792
rect 35894 25780 35900 25792
rect 35952 25780 35958 25832
rect 31726 25724 33916 25752
rect 6730 25684 6736 25696
rect 3988 25656 6736 25684
rect 6730 25644 6736 25656
rect 6788 25644 6794 25696
rect 10226 25644 10232 25696
rect 10284 25644 10290 25696
rect 14921 25687 14979 25693
rect 14921 25653 14933 25687
rect 14967 25684 14979 25687
rect 15010 25684 15016 25696
rect 14967 25656 15016 25684
rect 14967 25653 14979 25656
rect 14921 25647 14979 25653
rect 15010 25644 15016 25656
rect 15068 25644 15074 25696
rect 18325 25687 18383 25693
rect 18325 25653 18337 25687
rect 18371 25684 18383 25687
rect 19610 25684 19616 25696
rect 18371 25656 19616 25684
rect 18371 25653 18383 25656
rect 18325 25647 18383 25653
rect 19610 25644 19616 25656
rect 19668 25644 19674 25696
rect 29641 25687 29699 25693
rect 29641 25653 29653 25687
rect 29687 25684 29699 25687
rect 29914 25684 29920 25696
rect 29687 25656 29920 25684
rect 29687 25653 29699 25656
rect 29641 25647 29699 25653
rect 29914 25644 29920 25656
rect 29972 25644 29978 25696
rect 33781 25687 33839 25693
rect 33781 25653 33793 25687
rect 33827 25684 33839 25687
rect 33888 25684 33916 25724
rect 33965 25755 34023 25761
rect 33965 25721 33977 25755
rect 34011 25752 34023 25755
rect 35250 25752 35256 25764
rect 34011 25724 35256 25752
rect 34011 25721 34023 25724
rect 33965 25715 34023 25721
rect 35250 25712 35256 25724
rect 35308 25712 35314 25764
rect 36096 25752 36124 25860
rect 36170 25848 36176 25900
rect 36228 25848 36234 25900
rect 38746 25848 38752 25900
rect 38804 25848 38810 25900
rect 38933 25891 38991 25897
rect 38933 25857 38945 25891
rect 38979 25857 38991 25891
rect 38933 25851 38991 25857
rect 37642 25780 37648 25832
rect 37700 25820 37706 25832
rect 38948 25820 38976 25851
rect 39206 25848 39212 25900
rect 39264 25848 39270 25900
rect 40034 25848 40040 25900
rect 40092 25848 40098 25900
rect 40129 25891 40187 25897
rect 40129 25857 40141 25891
rect 40175 25888 40187 25891
rect 40310 25888 40316 25900
rect 40175 25860 40316 25888
rect 40175 25857 40187 25860
rect 40129 25851 40187 25857
rect 40310 25848 40316 25860
rect 40368 25848 40374 25900
rect 41509 25891 41567 25897
rect 41509 25857 41521 25891
rect 41555 25857 41567 25891
rect 41509 25851 41567 25857
rect 40402 25820 40408 25832
rect 37700 25792 38976 25820
rect 39040 25792 40408 25820
rect 37700 25780 37706 25792
rect 39040 25752 39068 25792
rect 40402 25780 40408 25792
rect 40460 25780 40466 25832
rect 41046 25780 41052 25832
rect 41104 25780 41110 25832
rect 41524 25752 41552 25851
rect 42610 25848 42616 25900
rect 42668 25848 42674 25900
rect 36096 25724 39068 25752
rect 40144 25724 41552 25752
rect 40144 25696 40172 25724
rect 33827 25656 33916 25684
rect 33827 25653 33839 25656
rect 33781 25647 33839 25653
rect 36078 25644 36084 25696
rect 36136 25644 36142 25696
rect 40126 25644 40132 25696
rect 40184 25644 40190 25696
rect 41230 25644 41236 25696
rect 41288 25644 41294 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 6362 25440 6368 25492
rect 6420 25480 6426 25492
rect 6733 25483 6791 25489
rect 6733 25480 6745 25483
rect 6420 25452 6745 25480
rect 6420 25440 6426 25452
rect 6733 25449 6745 25452
rect 6779 25480 6791 25483
rect 7190 25480 7196 25492
rect 6779 25452 7196 25480
rect 6779 25449 6791 25452
rect 6733 25443 6791 25449
rect 7190 25440 7196 25452
rect 7248 25440 7254 25492
rect 15657 25483 15715 25489
rect 15657 25449 15669 25483
rect 15703 25480 15715 25483
rect 15838 25480 15844 25492
rect 15703 25452 15844 25480
rect 15703 25449 15715 25452
rect 15657 25443 15715 25449
rect 15838 25440 15844 25452
rect 15896 25440 15902 25492
rect 22278 25440 22284 25492
rect 22336 25440 22342 25492
rect 25958 25440 25964 25492
rect 26016 25440 26022 25492
rect 34606 25440 34612 25492
rect 34664 25480 34670 25492
rect 36909 25483 36967 25489
rect 36909 25480 36921 25483
rect 34664 25452 36921 25480
rect 34664 25440 34670 25452
rect 36909 25449 36921 25452
rect 36955 25480 36967 25483
rect 39942 25480 39948 25492
rect 36955 25452 39948 25480
rect 36955 25449 36967 25452
rect 36909 25443 36967 25449
rect 39942 25440 39948 25452
rect 40000 25480 40006 25492
rect 41046 25480 41052 25492
rect 40000 25452 41052 25480
rect 40000 25440 40006 25452
rect 41046 25440 41052 25452
rect 41104 25440 41110 25492
rect 36538 25372 36544 25424
rect 36596 25372 36602 25424
rect 10778 25304 10784 25356
rect 10836 25304 10842 25356
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 28902 25304 28908 25356
rect 28960 25344 28966 25356
rect 29733 25347 29791 25353
rect 29733 25344 29745 25347
rect 28960 25316 29745 25344
rect 28960 25304 28966 25316
rect 29733 25313 29745 25316
rect 29779 25344 29791 25347
rect 32950 25344 32956 25356
rect 29779 25316 32956 25344
rect 29779 25313 29791 25316
rect 29733 25307 29791 25313
rect 32950 25304 32956 25316
rect 33008 25304 33014 25356
rect 36078 25304 36084 25356
rect 36136 25344 36142 25356
rect 36814 25344 36820 25356
rect 36136 25316 36820 25344
rect 36136 25304 36142 25316
rect 36814 25304 36820 25316
rect 36872 25344 36878 25356
rect 36872 25316 38056 25344
rect 36872 25304 36878 25316
rect 2038 25236 2044 25288
rect 2096 25236 2102 25288
rect 2314 25285 2320 25288
rect 2308 25239 2320 25285
rect 2314 25236 2320 25239
rect 2372 25236 2378 25288
rect 3602 25236 3608 25288
rect 3660 25276 3666 25288
rect 5353 25279 5411 25285
rect 5353 25276 5365 25279
rect 3660 25248 5365 25276
rect 3660 25236 3666 25248
rect 5353 25245 5365 25248
rect 5399 25276 5411 25279
rect 6546 25276 6552 25288
rect 5399 25248 6552 25276
rect 5399 25245 5411 25248
rect 5353 25239 5411 25245
rect 6546 25236 6552 25248
rect 6604 25276 6610 25288
rect 7466 25285 7472 25288
rect 7193 25279 7251 25285
rect 7193 25276 7205 25279
rect 6604 25248 7205 25276
rect 6604 25236 6610 25248
rect 7193 25245 7205 25248
rect 7239 25245 7251 25279
rect 7193 25239 7251 25245
rect 7460 25239 7472 25285
rect 7466 25236 7472 25239
rect 7524 25236 7530 25288
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 15010 25276 15016 25288
rect 14323 25248 15016 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 19426 25236 19432 25288
rect 19484 25236 19490 25288
rect 19610 25236 19616 25288
rect 19668 25236 19674 25288
rect 20898 25236 20904 25288
rect 20956 25236 20962 25288
rect 21168 25279 21226 25285
rect 21168 25245 21180 25279
rect 21214 25276 21226 25279
rect 21542 25276 21548 25288
rect 21214 25248 21548 25276
rect 21214 25245 21226 25248
rect 21168 25239 21226 25245
rect 21542 25236 21548 25248
rect 21600 25236 21606 25288
rect 24578 25236 24584 25288
rect 24636 25236 24642 25288
rect 24854 25285 24860 25288
rect 24848 25276 24860 25285
rect 24815 25248 24860 25276
rect 24848 25239 24860 25248
rect 24854 25236 24860 25239
rect 24912 25236 24918 25288
rect 30006 25236 30012 25288
rect 30064 25236 30070 25288
rect 37642 25236 37648 25288
rect 37700 25276 37706 25288
rect 38028 25285 38056 25316
rect 37737 25279 37795 25285
rect 37737 25276 37749 25279
rect 37700 25248 37749 25276
rect 37700 25236 37706 25248
rect 37737 25245 37749 25248
rect 37783 25245 37795 25279
rect 37737 25239 37795 25245
rect 38013 25279 38071 25285
rect 38013 25245 38025 25279
rect 38059 25276 38071 25279
rect 38746 25276 38752 25288
rect 38059 25248 38752 25276
rect 38059 25245 38071 25248
rect 38013 25239 38071 25245
rect 38746 25236 38752 25248
rect 38804 25236 38810 25288
rect 5620 25211 5678 25217
rect 5620 25177 5632 25211
rect 5666 25208 5678 25211
rect 5994 25208 6000 25220
rect 5666 25180 6000 25208
rect 5666 25177 5678 25180
rect 5620 25171 5678 25177
rect 5994 25168 6000 25180
rect 6052 25168 6058 25220
rect 14544 25211 14602 25217
rect 14544 25177 14556 25211
rect 14590 25208 14602 25211
rect 15378 25208 15384 25220
rect 14590 25180 15384 25208
rect 14590 25177 14602 25180
rect 14544 25171 14602 25177
rect 15378 25168 15384 25180
rect 15436 25168 15442 25220
rect 36909 25211 36967 25217
rect 36909 25177 36921 25211
rect 36955 25208 36967 25211
rect 37553 25211 37611 25217
rect 37553 25208 37565 25211
rect 36955 25180 37565 25208
rect 36955 25177 36967 25180
rect 36909 25171 36967 25177
rect 37553 25177 37565 25180
rect 37599 25177 37611 25211
rect 37553 25171 37611 25177
rect 3418 25100 3424 25152
rect 3476 25100 3482 25152
rect 7650 25100 7656 25152
rect 7708 25140 7714 25152
rect 8573 25143 8631 25149
rect 8573 25140 8585 25143
rect 7708 25112 8585 25140
rect 7708 25100 7714 25112
rect 8573 25109 8585 25112
rect 8619 25109 8631 25143
rect 8573 25103 8631 25109
rect 10318 25100 10324 25152
rect 10376 25100 10382 25152
rect 10689 25143 10747 25149
rect 10689 25109 10701 25143
rect 10735 25140 10747 25143
rect 10778 25140 10784 25152
rect 10735 25112 10784 25140
rect 10735 25109 10747 25112
rect 10689 25103 10747 25109
rect 10778 25100 10784 25112
rect 10836 25100 10842 25152
rect 19334 25100 19340 25152
rect 19392 25140 19398 25152
rect 19521 25143 19579 25149
rect 19521 25140 19533 25143
rect 19392 25112 19533 25140
rect 19392 25100 19398 25112
rect 19521 25109 19533 25112
rect 19567 25109 19579 25143
rect 19521 25103 19579 25109
rect 30374 25100 30380 25152
rect 30432 25140 30438 25152
rect 31113 25143 31171 25149
rect 31113 25140 31125 25143
rect 30432 25112 31125 25140
rect 30432 25100 30438 25112
rect 31113 25109 31125 25112
rect 31159 25109 31171 25143
rect 31113 25103 31171 25109
rect 37093 25143 37151 25149
rect 37093 25109 37105 25143
rect 37139 25140 37151 25143
rect 37274 25140 37280 25152
rect 37139 25112 37280 25140
rect 37139 25109 37151 25112
rect 37093 25103 37151 25109
rect 37274 25100 37280 25112
rect 37332 25100 37338 25152
rect 37918 25100 37924 25152
rect 37976 25100 37982 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 4982 24896 4988 24948
rect 5040 24896 5046 24948
rect 20165 24939 20223 24945
rect 20165 24905 20177 24939
rect 20211 24936 20223 24939
rect 20438 24936 20444 24948
rect 20211 24908 20444 24936
rect 20211 24905 20223 24908
rect 20165 24899 20223 24905
rect 20438 24896 20444 24908
rect 20496 24896 20502 24948
rect 29733 24939 29791 24945
rect 29733 24905 29745 24939
rect 29779 24936 29791 24939
rect 30006 24936 30012 24948
rect 29779 24908 30012 24936
rect 29779 24905 29791 24908
rect 29733 24899 29791 24905
rect 30006 24896 30012 24908
rect 30064 24896 30070 24948
rect 37642 24896 37648 24948
rect 37700 24936 37706 24948
rect 38378 24936 38384 24948
rect 37700 24908 38384 24936
rect 37700 24896 37706 24908
rect 38378 24896 38384 24908
rect 38436 24936 38442 24948
rect 38473 24939 38531 24945
rect 38473 24936 38485 24939
rect 38436 24908 38485 24936
rect 38436 24896 38442 24908
rect 38473 24905 38485 24908
rect 38519 24905 38531 24939
rect 38657 24939 38715 24945
rect 38657 24936 38669 24939
rect 38473 24899 38531 24905
rect 38580 24908 38669 24936
rect 10036 24871 10094 24877
rect 10036 24837 10048 24871
rect 10082 24868 10094 24871
rect 10226 24868 10232 24880
rect 10082 24840 10232 24868
rect 10082 24837 10094 24840
rect 10036 24831 10094 24837
rect 10226 24828 10232 24840
rect 10284 24828 10290 24880
rect 15010 24868 15016 24880
rect 13556 24840 15016 24868
rect 934 24760 940 24812
rect 992 24800 998 24812
rect 3878 24809 3884 24812
rect 1673 24803 1731 24809
rect 1673 24800 1685 24803
rect 992 24772 1685 24800
rect 992 24760 998 24772
rect 1673 24769 1685 24772
rect 1719 24769 1731 24803
rect 2593 24803 2651 24809
rect 2593 24800 2605 24803
rect 1673 24763 1731 24769
rect 1780 24772 2605 24800
rect 1026 24692 1032 24744
rect 1084 24732 1090 24744
rect 1780 24732 1808 24772
rect 2593 24769 2605 24772
rect 2639 24769 2651 24803
rect 3872 24800 3884 24809
rect 3839 24772 3884 24800
rect 2593 24763 2651 24769
rect 3872 24763 3884 24772
rect 3878 24760 3884 24763
rect 3936 24760 3942 24812
rect 13357 24803 13415 24809
rect 13357 24769 13369 24803
rect 13403 24800 13415 24803
rect 13556 24800 13584 24840
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 24578 24868 24584 24880
rect 24228 24840 24584 24868
rect 13630 24809 13636 24812
rect 13403 24772 13584 24800
rect 13403 24769 13415 24772
rect 13357 24763 13415 24769
rect 13624 24763 13636 24809
rect 13688 24800 13694 24812
rect 13688 24772 13724 24800
rect 13630 24760 13636 24763
rect 13688 24760 13694 24772
rect 16114 24760 16120 24812
rect 16172 24800 16178 24812
rect 19058 24809 19064 24812
rect 17109 24803 17167 24809
rect 17109 24800 17121 24803
rect 16172 24772 17121 24800
rect 16172 24760 16178 24772
rect 17109 24769 17121 24772
rect 17155 24769 17167 24803
rect 19052 24800 19064 24809
rect 19019 24772 19064 24800
rect 17109 24763 17167 24769
rect 19052 24763 19064 24772
rect 19058 24760 19064 24763
rect 19116 24760 19122 24812
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 20622 24800 20628 24812
rect 19668 24772 20628 24800
rect 19668 24760 19674 24772
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 24228 24809 24256 24840
rect 24578 24828 24584 24840
rect 24636 24828 24642 24880
rect 30098 24828 30104 24880
rect 30156 24868 30162 24880
rect 32309 24871 32367 24877
rect 32309 24868 32321 24871
rect 30156 24840 32321 24868
rect 30156 24828 30162 24840
rect 32309 24837 32321 24840
rect 32355 24868 32367 24871
rect 33502 24868 33508 24880
rect 32355 24840 33508 24868
rect 32355 24837 32367 24840
rect 32309 24831 32367 24837
rect 33502 24828 33508 24840
rect 33560 24828 33566 24880
rect 34606 24828 34612 24880
rect 34664 24828 34670 24880
rect 38580 24868 38608 24908
rect 38657 24905 38669 24908
rect 38703 24936 38715 24939
rect 39206 24936 39212 24948
rect 38703 24908 39212 24936
rect 38703 24905 38715 24908
rect 38657 24899 38715 24905
rect 39206 24896 39212 24908
rect 39264 24896 39270 24948
rect 37936 24840 38608 24868
rect 38672 24840 38884 24868
rect 37936 24812 37964 24840
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 24480 24803 24538 24809
rect 24480 24769 24492 24803
rect 24526 24800 24538 24803
rect 24762 24800 24768 24812
rect 24526 24772 24768 24800
rect 24526 24769 24538 24772
rect 24480 24763 24538 24769
rect 24762 24760 24768 24772
rect 24820 24760 24826 24812
rect 27341 24803 27399 24809
rect 27341 24769 27353 24803
rect 27387 24800 27399 24803
rect 27706 24800 27712 24812
rect 27387 24772 27712 24800
rect 27387 24769 27399 24772
rect 27341 24763 27399 24769
rect 27706 24760 27712 24772
rect 27764 24800 27770 24812
rect 28902 24800 28908 24812
rect 27764 24772 28908 24800
rect 27764 24760 27770 24772
rect 28902 24760 28908 24772
rect 28960 24760 28966 24812
rect 29914 24760 29920 24812
rect 29972 24760 29978 24812
rect 30193 24803 30251 24809
rect 30193 24769 30205 24803
rect 30239 24800 30251 24803
rect 30282 24800 30288 24812
rect 30239 24772 30288 24800
rect 30239 24769 30251 24772
rect 30193 24763 30251 24769
rect 30282 24760 30288 24772
rect 30340 24760 30346 24812
rect 30374 24760 30380 24812
rect 30432 24760 30438 24812
rect 32490 24760 32496 24812
rect 32548 24760 32554 24812
rect 32582 24760 32588 24812
rect 32640 24760 32646 24812
rect 33042 24760 33048 24812
rect 33100 24800 33106 24812
rect 34241 24803 34299 24809
rect 34241 24800 34253 24803
rect 33100 24772 34253 24800
rect 33100 24760 33106 24772
rect 34241 24769 34253 24772
rect 34287 24769 34299 24803
rect 34241 24763 34299 24769
rect 34422 24760 34428 24812
rect 34480 24760 34486 24812
rect 36354 24760 36360 24812
rect 36412 24800 36418 24812
rect 37918 24800 37924 24812
rect 36412 24772 37924 24800
rect 36412 24760 36418 24772
rect 37918 24760 37924 24772
rect 37976 24760 37982 24812
rect 38289 24803 38347 24809
rect 38289 24769 38301 24803
rect 38335 24800 38347 24803
rect 38672 24800 38700 24840
rect 38335 24772 38700 24800
rect 38335 24769 38347 24772
rect 38289 24763 38347 24769
rect 38746 24760 38752 24812
rect 38804 24760 38810 24812
rect 38856 24800 38884 24840
rect 40310 24800 40316 24812
rect 38856 24772 40316 24800
rect 40310 24760 40316 24772
rect 40368 24760 40374 24812
rect 40862 24809 40868 24812
rect 40856 24800 40868 24809
rect 40823 24772 40868 24800
rect 40856 24763 40868 24772
rect 40862 24760 40868 24763
rect 40920 24760 40926 24812
rect 1084 24704 1808 24732
rect 1084 24692 1090 24704
rect 2038 24692 2044 24744
rect 2096 24732 2102 24744
rect 3602 24732 3608 24744
rect 2096 24704 3608 24732
rect 2096 24692 2102 24704
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 9674 24692 9680 24744
rect 9732 24732 9738 24744
rect 9769 24735 9827 24741
rect 9769 24732 9781 24735
rect 9732 24704 9781 24732
rect 9732 24692 9738 24704
rect 9769 24701 9781 24704
rect 9815 24701 9827 24735
rect 9769 24695 9827 24701
rect 16853 24735 16911 24741
rect 16853 24701 16865 24735
rect 16899 24701 16911 24735
rect 16853 24695 16911 24701
rect 18785 24735 18843 24741
rect 18785 24701 18797 24735
rect 18831 24701 18843 24735
rect 18785 24695 18843 24701
rect 27617 24735 27675 24741
rect 27617 24701 27629 24735
rect 27663 24732 27675 24735
rect 27663 24704 28764 24732
rect 27663 24701 27675 24704
rect 27617 24695 27675 24701
rect 1949 24667 2007 24673
rect 1949 24633 1961 24667
rect 1995 24664 2007 24667
rect 3510 24664 3516 24676
rect 1995 24636 3516 24664
rect 1995 24633 2007 24636
rect 1949 24627 2007 24633
rect 3510 24624 3516 24636
rect 3568 24624 3574 24676
rect 2222 24556 2228 24608
rect 2280 24596 2286 24608
rect 2590 24596 2596 24608
rect 2280 24568 2596 24596
rect 2280 24556 2286 24568
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 2685 24599 2743 24605
rect 2685 24565 2697 24599
rect 2731 24596 2743 24599
rect 4890 24596 4896 24608
rect 2731 24568 4896 24596
rect 2731 24565 2743 24568
rect 2685 24559 2743 24565
rect 4890 24556 4896 24568
rect 4948 24556 4954 24608
rect 10686 24556 10692 24608
rect 10744 24596 10750 24608
rect 11149 24599 11207 24605
rect 11149 24596 11161 24599
rect 10744 24568 11161 24596
rect 10744 24556 10750 24568
rect 11149 24565 11161 24568
rect 11195 24565 11207 24599
rect 11149 24559 11207 24565
rect 14734 24556 14740 24608
rect 14792 24556 14798 24608
rect 15010 24556 15016 24608
rect 15068 24596 15074 24608
rect 16868 24596 16896 24695
rect 18800 24664 18828 24695
rect 20898 24664 20904 24676
rect 17788 24636 18828 24664
rect 17788 24596 17816 24636
rect 18800 24608 18828 24636
rect 19720 24636 20904 24664
rect 15068 24568 17816 24596
rect 15068 24556 15074 24568
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 17920 24568 18245 24596
rect 17920 24556 17926 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18233 24559 18291 24565
rect 18782 24556 18788 24608
rect 18840 24596 18846 24608
rect 19720 24596 19748 24636
rect 20898 24624 20904 24636
rect 20956 24624 20962 24676
rect 28736 24664 28764 24704
rect 28810 24692 28816 24744
rect 28868 24732 28874 24744
rect 30392 24732 30420 24760
rect 28868 24704 30420 24732
rect 38381 24735 38439 24741
rect 28868 24692 28874 24704
rect 38381 24701 38393 24735
rect 38427 24701 38439 24735
rect 38381 24695 38439 24701
rect 29730 24664 29736 24676
rect 25516 24636 27384 24664
rect 28736 24636 29736 24664
rect 18840 24568 19748 24596
rect 18840 24556 18846 24568
rect 20346 24556 20352 24608
rect 20404 24596 20410 24608
rect 25516 24596 25544 24636
rect 20404 24568 25544 24596
rect 20404 24556 20410 24568
rect 25590 24556 25596 24608
rect 25648 24556 25654 24608
rect 27356 24596 27384 24636
rect 29730 24624 29736 24636
rect 29788 24624 29794 24676
rect 33778 24624 33784 24676
rect 33836 24664 33842 24676
rect 35710 24664 35716 24676
rect 33836 24636 35716 24664
rect 33836 24624 33842 24636
rect 35710 24624 35716 24636
rect 35768 24624 35774 24676
rect 38396 24664 38424 24695
rect 40586 24692 40592 24744
rect 40644 24692 40650 24744
rect 38396 24636 40080 24664
rect 40052 24608 40080 24636
rect 28810 24596 28816 24608
rect 27356 24568 28816 24596
rect 28810 24556 28816 24568
rect 28868 24556 28874 24608
rect 28905 24599 28963 24605
rect 28905 24565 28917 24599
rect 28951 24596 28963 24599
rect 29362 24596 29368 24608
rect 28951 24568 29368 24596
rect 28951 24565 28963 24568
rect 28905 24559 28963 24565
rect 29362 24556 29368 24568
rect 29420 24596 29426 24608
rect 32214 24596 32220 24608
rect 29420 24568 32220 24596
rect 29420 24556 29426 24568
rect 32214 24556 32220 24568
rect 32272 24556 32278 24608
rect 32309 24599 32367 24605
rect 32309 24565 32321 24599
rect 32355 24596 32367 24599
rect 33134 24596 33140 24608
rect 32355 24568 33140 24596
rect 32355 24565 32367 24568
rect 32309 24559 32367 24565
rect 33134 24556 33140 24568
rect 33192 24556 33198 24608
rect 38105 24599 38163 24605
rect 38105 24565 38117 24599
rect 38151 24596 38163 24599
rect 39114 24596 39120 24608
rect 38151 24568 39120 24596
rect 38151 24565 38163 24568
rect 38105 24559 38163 24565
rect 39114 24556 39120 24568
rect 39172 24556 39178 24608
rect 40034 24556 40040 24608
rect 40092 24596 40098 24608
rect 41969 24599 42027 24605
rect 41969 24596 41981 24599
rect 40092 24568 41981 24596
rect 40092 24556 40098 24568
rect 41969 24565 41981 24568
rect 42015 24565 42027 24599
rect 41969 24559 42027 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1946 24352 1952 24404
rect 2004 24392 2010 24404
rect 2004 24364 11744 24392
rect 2004 24352 2010 24364
rect 11716 24324 11744 24364
rect 15930 24352 15936 24404
rect 15988 24352 15994 24404
rect 16114 24352 16120 24404
rect 16172 24352 16178 24404
rect 16500 24364 24716 24392
rect 16500 24324 16528 24364
rect 11716 24296 16528 24324
rect 19426 24284 19432 24336
rect 19484 24324 19490 24336
rect 19981 24327 20039 24333
rect 19981 24324 19993 24327
rect 19484 24296 19993 24324
rect 19484 24284 19490 24296
rect 19981 24293 19993 24296
rect 20027 24293 20039 24327
rect 24688 24324 24716 24364
rect 24762 24352 24768 24404
rect 24820 24352 24826 24404
rect 27617 24395 27675 24401
rect 24872 24364 27200 24392
rect 24872 24324 24900 24364
rect 24688 24296 24900 24324
rect 27172 24324 27200 24364
rect 27617 24361 27629 24395
rect 27663 24392 27675 24395
rect 28994 24392 29000 24404
rect 27663 24364 29000 24392
rect 27663 24361 27675 24364
rect 27617 24355 27675 24361
rect 28994 24352 29000 24364
rect 29052 24352 29058 24404
rect 36265 24395 36323 24401
rect 36265 24361 36277 24395
rect 36311 24392 36323 24395
rect 36354 24392 36360 24404
rect 36311 24364 36360 24392
rect 36311 24361 36323 24364
rect 36265 24355 36323 24361
rect 36354 24352 36360 24364
rect 36412 24352 36418 24404
rect 38378 24352 38384 24404
rect 38436 24352 38442 24404
rect 42337 24395 42395 24401
rect 42337 24361 42349 24395
rect 42383 24392 42395 24395
rect 42610 24392 42616 24404
rect 42383 24364 42616 24392
rect 42383 24361 42395 24364
rect 42337 24355 42395 24361
rect 42610 24352 42616 24364
rect 42668 24352 42674 24404
rect 29454 24324 29460 24336
rect 27172 24296 29460 24324
rect 19981 24287 20039 24293
rect 29454 24284 29460 24296
rect 29512 24284 29518 24336
rect 32309 24327 32367 24333
rect 32309 24293 32321 24327
rect 32355 24324 32367 24327
rect 32398 24324 32404 24336
rect 32355 24296 32404 24324
rect 32355 24293 32367 24296
rect 32309 24287 32367 24293
rect 32398 24284 32404 24296
rect 32456 24284 32462 24336
rect 14734 24216 14740 24268
rect 14792 24256 14798 24268
rect 19702 24256 19708 24268
rect 14792 24228 19708 24256
rect 14792 24216 14798 24228
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 20956 24228 21373 24256
rect 20956 24216 20962 24228
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 21361 24219 21419 24225
rect 24578 24216 24584 24268
rect 24636 24256 24642 24268
rect 24636 24228 26280 24256
rect 24636 24216 24642 24228
rect 1670 24148 1676 24200
rect 1728 24188 1734 24200
rect 2038 24188 2044 24200
rect 1728 24160 2044 24188
rect 1728 24148 1734 24160
rect 2038 24148 2044 24160
rect 2096 24148 2102 24200
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 4672 24160 6914 24188
rect 4672 24148 4678 24160
rect 2308 24123 2366 24129
rect 2308 24089 2320 24123
rect 2354 24120 2366 24123
rect 2498 24120 2504 24132
rect 2354 24092 2504 24120
rect 2354 24089 2366 24092
rect 2308 24083 2366 24089
rect 2498 24080 2504 24092
rect 2556 24080 2562 24132
rect 6886 24120 6914 24160
rect 9674 24148 9680 24200
rect 9732 24188 9738 24200
rect 10229 24191 10287 24197
rect 10229 24188 10241 24191
rect 9732 24160 10241 24188
rect 9732 24148 9738 24160
rect 10229 24157 10241 24160
rect 10275 24157 10287 24191
rect 10229 24151 10287 24157
rect 10318 24148 10324 24200
rect 10376 24188 10382 24200
rect 10485 24191 10543 24197
rect 10485 24188 10497 24191
rect 10376 24160 10497 24188
rect 10376 24148 10382 24160
rect 10485 24157 10497 24160
rect 10531 24157 10543 24191
rect 10485 24151 10543 24157
rect 15562 24148 15568 24200
rect 15620 24148 15626 24200
rect 17862 24148 17868 24200
rect 17920 24188 17926 24200
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 17920 24160 19809 24188
rect 17920 24148 17926 24160
rect 19797 24157 19809 24160
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 25222 24148 25228 24200
rect 25280 24148 25286 24200
rect 26252 24197 26280 24228
rect 31754 24216 31760 24268
rect 31812 24256 31818 24268
rect 31941 24259 31999 24265
rect 31941 24256 31953 24259
rect 31812 24228 31953 24256
rect 31812 24216 31818 24228
rect 31941 24225 31953 24228
rect 31987 24256 31999 24259
rect 32582 24256 32588 24268
rect 31987 24228 32588 24256
rect 31987 24225 31999 24228
rect 31941 24219 31999 24225
rect 32582 24216 32588 24228
rect 32640 24216 32646 24268
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24188 26295 24191
rect 27706 24188 27712 24200
rect 26283 24160 27712 24188
rect 26283 24157 26295 24160
rect 26237 24151 26295 24157
rect 27706 24148 27712 24160
rect 27764 24148 27770 24200
rect 32861 24191 32919 24197
rect 32861 24157 32873 24191
rect 32907 24188 32919 24191
rect 32950 24188 32956 24200
rect 32907 24160 32956 24188
rect 32907 24157 32919 24160
rect 32861 24151 32919 24157
rect 32950 24148 32956 24160
rect 33008 24148 33014 24200
rect 33134 24197 33140 24200
rect 33128 24188 33140 24197
rect 33095 24160 33140 24188
rect 33128 24151 33140 24160
rect 33134 24148 33140 24151
rect 33192 24148 33198 24200
rect 34885 24191 34943 24197
rect 34885 24157 34897 24191
rect 34931 24188 34943 24191
rect 36538 24188 36544 24200
rect 34931 24160 36544 24188
rect 34931 24157 34943 24160
rect 34885 24151 34943 24157
rect 36538 24148 36544 24160
rect 36596 24188 36602 24200
rect 37274 24197 37280 24200
rect 37001 24191 37059 24197
rect 37001 24188 37013 24191
rect 36596 24160 37013 24188
rect 36596 24148 36602 24160
rect 37001 24157 37013 24160
rect 37047 24157 37059 24191
rect 37268 24188 37280 24197
rect 37235 24160 37280 24188
rect 37001 24151 37059 24157
rect 37268 24151 37280 24160
rect 37274 24148 37280 24151
rect 37332 24148 37338 24200
rect 39114 24148 39120 24200
rect 39172 24148 39178 24200
rect 39209 24191 39267 24197
rect 39209 24157 39221 24191
rect 39255 24188 39267 24191
rect 40126 24188 40132 24200
rect 39255 24160 40132 24188
rect 39255 24157 39267 24160
rect 39209 24151 39267 24157
rect 40126 24148 40132 24160
rect 40184 24148 40190 24200
rect 40218 24148 40224 24200
rect 40276 24188 40282 24200
rect 40586 24188 40592 24200
rect 40276 24160 40592 24188
rect 40276 24148 40282 24160
rect 40586 24148 40592 24160
rect 40644 24188 40650 24200
rect 41230 24197 41236 24200
rect 40957 24191 41015 24197
rect 40957 24188 40969 24191
rect 40644 24160 40969 24188
rect 40644 24148 40650 24160
rect 40957 24157 40969 24160
rect 41003 24157 41015 24191
rect 41224 24188 41236 24197
rect 41191 24160 41236 24188
rect 40957 24151 41015 24157
rect 41224 24151 41236 24160
rect 41230 24148 41236 24151
rect 41288 24148 41294 24200
rect 11330 24120 11336 24132
rect 6886 24092 11336 24120
rect 11330 24080 11336 24092
rect 11388 24080 11394 24132
rect 15933 24123 15991 24129
rect 15933 24089 15945 24123
rect 15979 24120 15991 24123
rect 16574 24120 16580 24132
rect 15979 24092 16580 24120
rect 15979 24089 15991 24092
rect 15933 24083 15991 24089
rect 16574 24080 16580 24092
rect 16632 24080 16638 24132
rect 19429 24123 19487 24129
rect 19429 24089 19441 24123
rect 19475 24120 19487 24123
rect 19475 24092 20484 24120
rect 19475 24089 19487 24092
rect 19429 24083 19487 24089
rect 3421 24055 3479 24061
rect 3421 24021 3433 24055
rect 3467 24052 3479 24055
rect 4798 24052 4804 24064
rect 3467 24024 4804 24052
rect 3467 24021 3479 24024
rect 3421 24015 3479 24021
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 10778 24012 10784 24064
rect 10836 24052 10842 24064
rect 11609 24055 11667 24061
rect 11609 24052 11621 24055
rect 10836 24024 11621 24052
rect 10836 24012 10842 24024
rect 11609 24021 11621 24024
rect 11655 24021 11667 24055
rect 11609 24015 11667 24021
rect 19610 24012 19616 24064
rect 19668 24012 19674 24064
rect 19702 24012 19708 24064
rect 19760 24012 19766 24064
rect 20456 24052 20484 24092
rect 20530 24080 20536 24132
rect 20588 24120 20594 24132
rect 21606 24123 21664 24129
rect 21606 24120 21618 24123
rect 20588 24092 21618 24120
rect 20588 24080 20594 24092
rect 21606 24089 21618 24092
rect 21652 24089 21664 24123
rect 21606 24083 21664 24089
rect 25133 24123 25191 24129
rect 25133 24089 25145 24123
rect 25179 24120 25191 24123
rect 25590 24120 25596 24132
rect 25179 24092 25596 24120
rect 25179 24089 25191 24092
rect 25133 24083 25191 24089
rect 25590 24080 25596 24092
rect 25648 24080 25654 24132
rect 26142 24080 26148 24132
rect 26200 24120 26206 24132
rect 26482 24123 26540 24129
rect 26482 24120 26494 24123
rect 26200 24092 26494 24120
rect 26200 24080 26206 24092
rect 26482 24089 26494 24092
rect 26528 24089 26540 24123
rect 26482 24083 26540 24089
rect 34790 24080 34796 24132
rect 34848 24120 34854 24132
rect 35130 24123 35188 24129
rect 35130 24120 35142 24123
rect 34848 24092 35142 24120
rect 34848 24080 34854 24092
rect 35130 24089 35142 24092
rect 35176 24089 35188 24123
rect 35130 24083 35188 24089
rect 36170 24080 36176 24132
rect 36228 24120 36234 24132
rect 38841 24123 38899 24129
rect 38841 24120 38853 24123
rect 36228 24092 38853 24120
rect 36228 24080 36234 24092
rect 38841 24089 38853 24092
rect 38887 24089 38899 24123
rect 38841 24083 38899 24089
rect 20990 24052 20996 24064
rect 20456 24024 20996 24052
rect 20990 24012 20996 24024
rect 21048 24052 21054 24064
rect 22741 24055 22799 24061
rect 22741 24052 22753 24055
rect 21048 24024 22753 24052
rect 21048 24012 21054 24024
rect 22741 24021 22753 24024
rect 22787 24021 22799 24055
rect 22741 24015 22799 24021
rect 30558 24012 30564 24064
rect 30616 24052 30622 24064
rect 32401 24055 32459 24061
rect 32401 24052 32413 24055
rect 30616 24024 32413 24052
rect 30616 24012 30622 24024
rect 32401 24021 32413 24024
rect 32447 24021 32459 24055
rect 32401 24015 32459 24021
rect 34241 24055 34299 24061
rect 34241 24021 34253 24055
rect 34287 24052 34299 24055
rect 34606 24052 34612 24064
rect 34287 24024 34612 24052
rect 34287 24021 34299 24024
rect 34241 24015 34299 24021
rect 34606 24012 34612 24024
rect 34664 24012 34670 24064
rect 38930 24012 38936 24064
rect 38988 24052 38994 24064
rect 39025 24055 39083 24061
rect 39025 24052 39037 24055
rect 38988 24024 39037 24052
rect 38988 24012 38994 24024
rect 39025 24021 39037 24024
rect 39071 24021 39083 24055
rect 39025 24015 39083 24021
rect 39390 24012 39396 24064
rect 39448 24012 39454 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1946 23808 1952 23860
rect 2004 23808 2010 23860
rect 2498 23808 2504 23860
rect 2556 23808 2562 23860
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 2961 23851 3019 23857
rect 2961 23848 2973 23851
rect 2832 23820 2973 23848
rect 2832 23808 2838 23820
rect 2961 23817 2973 23820
rect 3007 23817 3019 23851
rect 2961 23811 3019 23817
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 3568 23820 22094 23848
rect 3568 23808 3574 23820
rect 4893 23783 4951 23789
rect 4893 23749 4905 23783
rect 4939 23780 4951 23783
rect 4982 23780 4988 23792
rect 4939 23752 4988 23780
rect 4939 23749 4951 23752
rect 4893 23743 4951 23749
rect 4982 23740 4988 23752
rect 5040 23740 5046 23792
rect 16945 23783 17003 23789
rect 16945 23749 16957 23783
rect 16991 23749 17003 23783
rect 16945 23743 17003 23749
rect 934 23672 940 23724
rect 992 23712 998 23724
rect 1673 23715 1731 23721
rect 1673 23712 1685 23715
rect 992 23684 1685 23712
rect 992 23672 998 23684
rect 1673 23681 1685 23684
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 2869 23715 2927 23721
rect 2869 23681 2881 23715
rect 2915 23712 2927 23715
rect 2915 23684 4844 23712
rect 2915 23681 2927 23684
rect 2869 23675 2927 23681
rect 4816 23656 4844 23684
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 6546 23672 6552 23724
rect 6604 23672 6610 23724
rect 6638 23672 6644 23724
rect 6696 23712 6702 23724
rect 6805 23715 6863 23721
rect 6805 23712 6817 23715
rect 6696 23684 6817 23712
rect 6696 23672 6702 23684
rect 6805 23681 6817 23684
rect 6851 23681 6863 23715
rect 16960 23712 16988 23743
rect 17034 23740 17040 23792
rect 17092 23780 17098 23792
rect 17145 23783 17203 23789
rect 17145 23780 17157 23783
rect 17092 23752 17157 23780
rect 17092 23740 17098 23752
rect 17145 23749 17157 23752
rect 17191 23749 17203 23783
rect 17145 23743 17203 23749
rect 20070 23740 20076 23792
rect 20128 23740 20134 23792
rect 20530 23740 20536 23792
rect 20588 23740 20594 23792
rect 22066 23780 22094 23820
rect 26142 23808 26148 23860
rect 26200 23808 26206 23860
rect 26252 23820 31708 23848
rect 26252 23780 26280 23820
rect 22066 23752 26280 23780
rect 28721 23783 28779 23789
rect 28721 23749 28733 23783
rect 28767 23749 28779 23783
rect 28721 23743 28779 23749
rect 17862 23712 17868 23724
rect 16960 23684 17868 23712
rect 6805 23675 6863 23681
rect 17144 23656 17172 23684
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 20257 23715 20315 23721
rect 20257 23681 20269 23715
rect 20303 23712 20315 23715
rect 20303 23684 20668 23712
rect 20303 23681 20315 23684
rect 20257 23675 20315 23681
rect 2958 23604 2964 23656
rect 3016 23644 3022 23656
rect 3053 23647 3111 23653
rect 3053 23644 3065 23647
rect 3016 23616 3065 23644
rect 3016 23604 3022 23616
rect 3053 23613 3065 23616
rect 3099 23613 3111 23647
rect 3053 23607 3111 23613
rect 4798 23604 4804 23656
rect 4856 23644 4862 23656
rect 4985 23647 5043 23653
rect 4985 23644 4997 23647
rect 4856 23616 4997 23644
rect 4856 23604 4862 23616
rect 4985 23613 4997 23616
rect 5031 23613 5043 23647
rect 4985 23607 5043 23613
rect 17126 23604 17132 23656
rect 17184 23604 17190 23656
rect 20438 23604 20444 23656
rect 20496 23604 20502 23656
rect 20640 23644 20668 23684
rect 20990 23672 20996 23724
rect 21048 23672 21054 23724
rect 26326 23672 26332 23724
rect 26384 23672 26390 23724
rect 28736 23712 28764 23743
rect 29362 23740 29368 23792
rect 29420 23740 29426 23792
rect 31680 23780 31708 23820
rect 31754 23808 31760 23860
rect 31812 23808 31818 23860
rect 32490 23808 32496 23860
rect 32548 23808 32554 23860
rect 40310 23808 40316 23860
rect 40368 23848 40374 23860
rect 41785 23851 41843 23857
rect 41785 23848 41797 23851
rect 40368 23820 41797 23848
rect 40368 23808 40374 23820
rect 41785 23817 41797 23820
rect 41831 23817 41843 23851
rect 41785 23811 41843 23817
rect 36722 23780 36728 23792
rect 31680 23752 36728 23780
rect 36722 23740 36728 23752
rect 36780 23740 36786 23792
rect 39390 23740 39396 23792
rect 39448 23780 39454 23792
rect 40650 23783 40708 23789
rect 40650 23780 40662 23783
rect 39448 23752 40662 23780
rect 39448 23740 39454 23752
rect 40650 23749 40662 23752
rect 40696 23749 40708 23783
rect 40650 23743 40708 23749
rect 28736 23684 29316 23712
rect 21085 23647 21143 23653
rect 21085 23644 21097 23647
rect 20640 23616 21097 23644
rect 21085 23613 21097 23616
rect 21131 23613 21143 23647
rect 21085 23607 21143 23613
rect 26605 23647 26663 23653
rect 26605 23613 26617 23647
rect 26651 23644 26663 23647
rect 26651 23616 28948 23644
rect 26651 23613 26663 23616
rect 26605 23607 26663 23613
rect 5000 23548 6592 23576
rect 5000 23517 5028 23548
rect 6564 23520 6592 23548
rect 7742 23536 7748 23588
rect 7800 23576 7806 23588
rect 9858 23576 9864 23588
rect 7800 23548 9864 23576
rect 7800 23536 7806 23548
rect 9858 23536 9864 23548
rect 9916 23536 9922 23588
rect 15562 23536 15568 23588
rect 15620 23576 15626 23588
rect 17313 23579 17371 23585
rect 17313 23576 17325 23579
rect 15620 23548 17325 23576
rect 15620 23536 15626 23548
rect 17313 23545 17325 23548
rect 17359 23545 17371 23579
rect 17313 23539 17371 23545
rect 28258 23536 28264 23588
rect 28316 23576 28322 23588
rect 28920 23585 28948 23616
rect 28353 23579 28411 23585
rect 28353 23576 28365 23579
rect 28316 23548 28365 23576
rect 28316 23536 28322 23548
rect 28353 23545 28365 23548
rect 28399 23545 28411 23579
rect 28353 23539 28411 23545
rect 28905 23579 28963 23585
rect 28905 23545 28917 23579
rect 28951 23545 28963 23579
rect 29288 23576 29316 23684
rect 30190 23672 30196 23724
rect 30248 23672 30254 23724
rect 30466 23672 30472 23724
rect 30524 23712 30530 23724
rect 31389 23715 31447 23721
rect 31389 23712 31401 23715
rect 30524 23684 31401 23712
rect 30524 23672 30530 23684
rect 31389 23681 31401 23684
rect 31435 23681 31447 23715
rect 31389 23675 31447 23681
rect 32306 23672 32312 23724
rect 32364 23672 32370 23724
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 33045 23715 33103 23721
rect 33045 23681 33057 23715
rect 33091 23712 33103 23715
rect 34606 23712 34612 23724
rect 33091 23684 34612 23712
rect 33091 23681 33103 23684
rect 33045 23675 33103 23681
rect 31481 23647 31539 23653
rect 31481 23613 31493 23647
rect 31527 23644 31539 23647
rect 31754 23644 31760 23656
rect 31527 23616 31760 23644
rect 31527 23613 31539 23616
rect 31481 23607 31539 23613
rect 31754 23604 31760 23616
rect 31812 23644 31818 23656
rect 32508 23644 32536 23675
rect 34606 23672 34612 23684
rect 34664 23672 34670 23724
rect 31812 23616 33088 23644
rect 31812 23604 31818 23616
rect 33060 23588 33088 23616
rect 33318 23604 33324 23656
rect 33376 23604 33382 23656
rect 40218 23604 40224 23656
rect 40276 23644 40282 23656
rect 40405 23647 40463 23653
rect 40405 23644 40417 23647
rect 40276 23616 40417 23644
rect 40276 23604 40282 23616
rect 40405 23613 40417 23616
rect 40451 23613 40463 23647
rect 40405 23607 40463 23613
rect 31202 23576 31208 23588
rect 29288 23548 31208 23576
rect 28905 23539 28963 23545
rect 31202 23536 31208 23548
rect 31260 23536 31266 23588
rect 33042 23536 33048 23588
rect 33100 23536 33106 23588
rect 4985 23511 5043 23517
rect 4985 23477 4997 23511
rect 5031 23477 5043 23511
rect 4985 23471 5043 23477
rect 5074 23468 5080 23520
rect 5132 23508 5138 23520
rect 5353 23511 5411 23517
rect 5353 23508 5365 23511
rect 5132 23480 5365 23508
rect 5132 23468 5138 23480
rect 5353 23477 5365 23480
rect 5399 23477 5411 23511
rect 5353 23471 5411 23477
rect 6546 23468 6552 23520
rect 6604 23508 6610 23520
rect 7929 23511 7987 23517
rect 7929 23508 7941 23511
rect 6604 23480 7941 23508
rect 6604 23468 6610 23480
rect 7929 23477 7941 23480
rect 7975 23477 7987 23511
rect 7929 23471 7987 23477
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 13446 23508 13452 23520
rect 11756 23480 13452 23508
rect 11756 23468 11762 23480
rect 13446 23468 13452 23480
rect 13504 23468 13510 23520
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 17129 23511 17187 23517
rect 17129 23508 17141 23511
rect 16908 23480 17141 23508
rect 16908 23468 16914 23480
rect 17129 23477 17141 23480
rect 17175 23508 17187 23511
rect 17770 23508 17776 23520
rect 17175 23480 17776 23508
rect 17175 23477 17187 23480
rect 17129 23471 17187 23477
rect 17770 23468 17776 23480
rect 17828 23468 17834 23520
rect 18874 23468 18880 23520
rect 18932 23508 18938 23520
rect 20349 23511 20407 23517
rect 20349 23508 20361 23511
rect 18932 23480 20361 23508
rect 18932 23468 18938 23480
rect 20349 23477 20361 23480
rect 20395 23477 20407 23511
rect 20349 23471 20407 23477
rect 26510 23468 26516 23520
rect 26568 23468 26574 23520
rect 28721 23511 28779 23517
rect 28721 23477 28733 23511
rect 28767 23508 28779 23511
rect 28994 23508 29000 23520
rect 28767 23480 29000 23508
rect 28767 23477 28779 23480
rect 28721 23471 28779 23477
rect 28994 23468 29000 23480
rect 29052 23468 29058 23520
rect 31573 23511 31631 23517
rect 31573 23477 31585 23511
rect 31619 23508 31631 23511
rect 32306 23508 32312 23520
rect 31619 23480 32312 23508
rect 31619 23477 31631 23480
rect 31573 23471 31631 23477
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 6273 23307 6331 23313
rect 6273 23273 6285 23307
rect 6319 23304 6331 23307
rect 6638 23304 6644 23316
rect 6319 23276 6644 23304
rect 6319 23273 6331 23276
rect 6273 23267 6331 23273
rect 6638 23264 6644 23276
rect 6696 23264 6702 23316
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 7469 23307 7527 23313
rect 7469 23304 7481 23307
rect 7248 23276 7481 23304
rect 7248 23264 7254 23276
rect 7469 23273 7481 23276
rect 7515 23273 7527 23307
rect 7469 23267 7527 23273
rect 13538 23264 13544 23316
rect 13596 23264 13602 23316
rect 16574 23264 16580 23316
rect 16632 23264 16638 23316
rect 26053 23307 26111 23313
rect 26053 23273 26065 23307
rect 26099 23273 26111 23307
rect 26053 23267 26111 23273
rect 26237 23307 26295 23313
rect 26237 23273 26249 23307
rect 26283 23304 26295 23307
rect 26510 23304 26516 23316
rect 26283 23276 26516 23304
rect 26283 23273 26295 23276
rect 26237 23267 26295 23273
rect 3418 23196 3424 23248
rect 3476 23236 3482 23248
rect 3476 23208 7512 23236
rect 3476 23196 3482 23208
rect 1026 23128 1032 23180
rect 1084 23168 1090 23180
rect 1765 23171 1823 23177
rect 1765 23168 1777 23171
rect 1084 23140 1777 23168
rect 1084 23128 1090 23140
rect 1765 23137 1777 23140
rect 1811 23137 1823 23171
rect 1765 23131 1823 23137
rect 2958 23128 2964 23180
rect 3016 23168 3022 23180
rect 4985 23171 5043 23177
rect 4985 23168 4997 23171
rect 3016 23140 4997 23168
rect 3016 23128 3022 23140
rect 4985 23137 4997 23140
rect 5031 23168 5043 23171
rect 6825 23171 6883 23177
rect 6825 23168 6837 23171
rect 5031 23140 6837 23168
rect 5031 23137 5043 23140
rect 4985 23131 5043 23137
rect 6825 23137 6837 23140
rect 6871 23168 6883 23171
rect 7282 23168 7288 23180
rect 6871 23140 7288 23168
rect 6871 23137 6883 23140
rect 6825 23131 6883 23137
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 7484 23109 7512 23208
rect 16942 23196 16948 23248
rect 17000 23196 17006 23248
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17681 23239 17739 23245
rect 17681 23236 17693 23239
rect 17092 23208 17693 23236
rect 17092 23196 17098 23208
rect 17681 23205 17693 23208
rect 17727 23205 17739 23239
rect 26068 23236 26096 23267
rect 26510 23264 26516 23276
rect 26568 23264 26574 23316
rect 29730 23264 29736 23316
rect 29788 23264 29794 23316
rect 32953 23307 33011 23313
rect 32953 23273 32965 23307
rect 32999 23304 33011 23307
rect 33042 23304 33048 23316
rect 32999 23276 33048 23304
rect 32999 23273 33011 23276
rect 32953 23267 33011 23273
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 42150 23264 42156 23316
rect 42208 23264 42214 23316
rect 28718 23236 28724 23248
rect 26068 23208 28724 23236
rect 17681 23199 17739 23205
rect 28718 23196 28724 23208
rect 28776 23196 28782 23248
rect 30101 23239 30159 23245
rect 30101 23205 30113 23239
rect 30147 23236 30159 23239
rect 30558 23236 30564 23248
rect 30147 23208 30564 23236
rect 30147 23205 30159 23208
rect 30101 23199 30159 23205
rect 30558 23196 30564 23208
rect 30616 23196 30622 23248
rect 7650 23128 7656 23180
rect 7708 23128 7714 23180
rect 16960 23168 16988 23196
rect 28077 23171 28135 23177
rect 16960 23140 18000 23168
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 7469 23103 7527 23109
rect 1627 23072 6914 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 2593 23035 2651 23041
rect 2593 23032 2605 23035
rect 1964 23004 2605 23032
rect 934 22924 940 22976
rect 992 22964 998 22976
rect 1964 22964 1992 23004
rect 2593 23001 2605 23004
rect 2639 23001 2651 23035
rect 2593 22995 2651 23001
rect 4801 23035 4859 23041
rect 4801 23001 4813 23035
rect 4847 23032 4859 23035
rect 5166 23032 5172 23044
rect 4847 23004 5172 23032
rect 4847 23001 4859 23004
rect 4801 22995 4859 23001
rect 5166 22992 5172 23004
rect 5224 22992 5230 23044
rect 6730 22992 6736 23044
rect 6788 22992 6794 23044
rect 6886 23032 6914 23072
rect 7469 23069 7481 23103
rect 7515 23069 7527 23103
rect 7469 23063 7527 23069
rect 7742 23060 7748 23112
rect 7800 23060 7806 23112
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23100 12219 23103
rect 12894 23100 12900 23112
rect 12207 23072 12900 23100
rect 12207 23069 12219 23072
rect 12161 23063 12219 23069
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 16758 23060 16764 23112
rect 16816 23060 16822 23112
rect 16850 23060 16856 23112
rect 16908 23060 16914 23112
rect 16945 23103 17003 23109
rect 16945 23069 16957 23103
rect 16991 23069 17003 23103
rect 16945 23063 17003 23069
rect 17037 23103 17095 23109
rect 17037 23069 17049 23103
rect 17083 23100 17095 23103
rect 17126 23100 17132 23112
rect 17083 23072 17132 23100
rect 17083 23069 17095 23072
rect 17037 23063 17095 23069
rect 12428 23035 12486 23041
rect 6886 23004 12388 23032
rect 992 22936 1992 22964
rect 992 22924 998 22936
rect 2406 22924 2412 22976
rect 2464 22964 2470 22976
rect 2685 22967 2743 22973
rect 2685 22964 2697 22967
rect 2464 22936 2697 22964
rect 2464 22924 2470 22936
rect 2685 22933 2697 22936
rect 2731 22933 2743 22967
rect 2685 22927 2743 22933
rect 4430 22924 4436 22976
rect 4488 22924 4494 22976
rect 4890 22924 4896 22976
rect 4948 22924 4954 22976
rect 6638 22924 6644 22976
rect 6696 22924 6702 22976
rect 7929 22967 7987 22973
rect 7929 22933 7941 22967
rect 7975 22964 7987 22967
rect 8202 22964 8208 22976
rect 7975 22936 8208 22964
rect 7975 22933 7987 22936
rect 7929 22927 7987 22933
rect 8202 22924 8208 22936
rect 8260 22924 8266 22976
rect 12360 22964 12388 23004
rect 12428 23001 12440 23035
rect 12474 23032 12486 23035
rect 12802 23032 12808 23044
rect 12474 23004 12808 23032
rect 12474 23001 12486 23004
rect 12428 22995 12486 23001
rect 12802 22992 12808 23004
rect 12860 22992 12866 23044
rect 14642 23032 14648 23044
rect 13464 23004 14648 23032
rect 13464 22964 13492 23004
rect 14642 22992 14648 23004
rect 14700 22992 14706 23044
rect 12360 22936 13492 22964
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 16960 22964 16988 23063
rect 17126 23060 17132 23072
rect 17184 23060 17190 23112
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 17972 23109 18000 23140
rect 28077 23137 28089 23171
rect 28123 23168 28135 23171
rect 28258 23168 28264 23180
rect 28123 23140 28264 23168
rect 28123 23137 28135 23140
rect 28077 23131 28135 23137
rect 28258 23128 28264 23140
rect 28316 23168 28322 23180
rect 28316 23140 29960 23168
rect 28316 23128 28322 23140
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 17828 23072 17877 23100
rect 17828 23060 17834 23072
rect 17865 23069 17877 23072
rect 17911 23069 17923 23103
rect 17865 23063 17923 23069
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 20864 23072 21189 23100
rect 20864 23060 20870 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 22186 23060 22192 23112
rect 22244 23100 22250 23112
rect 22244 23072 25912 23100
rect 22244 23060 22250 23072
rect 17681 23035 17739 23041
rect 17681 23001 17693 23035
rect 17727 23032 17739 23035
rect 20254 23032 20260 23044
rect 17727 23004 20260 23032
rect 17727 23001 17739 23004
rect 17681 22995 17739 23001
rect 20254 22992 20260 23004
rect 20312 23032 20318 23044
rect 20438 23032 20444 23044
rect 20312 23004 20444 23032
rect 20312 22992 20318 23004
rect 20438 22992 20444 23004
rect 20496 22992 20502 23044
rect 21358 22992 21364 23044
rect 21416 23032 21422 23044
rect 25884 23041 25912 23072
rect 28350 23060 28356 23112
rect 28408 23060 28414 23112
rect 28442 23060 28448 23112
rect 28500 23060 28506 23112
rect 28537 23103 28595 23109
rect 28537 23069 28549 23103
rect 28583 23069 28595 23103
rect 28537 23063 28595 23069
rect 25869 23035 25927 23041
rect 21416 23004 22232 23032
rect 21416 22992 21422 23004
rect 16908 22936 16988 22964
rect 21269 22967 21327 22973
rect 16908 22924 16914 22936
rect 21269 22933 21281 22967
rect 21315 22964 21327 22967
rect 22094 22964 22100 22976
rect 21315 22936 22100 22964
rect 21315 22933 21327 22936
rect 21269 22927 21327 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22204 22964 22232 23004
rect 25869 23001 25881 23035
rect 25915 23032 25927 23035
rect 28552 23032 28580 23063
rect 28718 23060 28724 23112
rect 28776 23060 28782 23112
rect 29932 23109 29960 23140
rect 35894 23128 35900 23180
rect 35952 23168 35958 23180
rect 36262 23168 36268 23180
rect 35952 23140 36268 23168
rect 35952 23128 35958 23140
rect 36262 23128 36268 23140
rect 36320 23168 36326 23180
rect 36320 23140 36584 23168
rect 36320 23128 36326 23140
rect 29917 23103 29975 23109
rect 29917 23069 29929 23103
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 30006 23060 30012 23112
rect 30064 23060 30070 23112
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23100 30251 23103
rect 30650 23100 30656 23112
rect 30239 23072 30656 23100
rect 30239 23069 30251 23072
rect 30193 23063 30251 23069
rect 30650 23060 30656 23072
rect 30708 23060 30714 23112
rect 32122 23100 32128 23112
rect 31726 23072 32128 23100
rect 25915 23004 28580 23032
rect 25915 23001 25927 23004
rect 25869 22995 25927 23001
rect 29178 22992 29184 23044
rect 29236 23032 29242 23044
rect 31386 23032 31392 23044
rect 29236 23004 31392 23032
rect 29236 22992 29242 23004
rect 31386 22992 31392 23004
rect 31444 23032 31450 23044
rect 31726 23032 31754 23072
rect 32122 23060 32128 23072
rect 32180 23100 32186 23112
rect 32861 23103 32919 23109
rect 32861 23100 32873 23103
rect 32180 23072 32873 23100
rect 32180 23060 32186 23072
rect 32861 23069 32873 23072
rect 32907 23100 32919 23103
rect 33318 23100 33324 23112
rect 32907 23072 33324 23100
rect 32907 23069 32919 23072
rect 32861 23063 32919 23069
rect 33318 23060 33324 23072
rect 33376 23100 33382 23112
rect 35434 23100 35440 23112
rect 33376 23072 35440 23100
rect 33376 23060 33382 23072
rect 35434 23060 35440 23072
rect 35492 23100 35498 23112
rect 36170 23100 36176 23112
rect 35492 23072 36176 23100
rect 35492 23060 35498 23072
rect 36170 23060 36176 23072
rect 36228 23100 36234 23112
rect 36556 23109 36584 23140
rect 37366 23128 37372 23180
rect 37424 23168 37430 23180
rect 38565 23171 38623 23177
rect 38565 23168 38577 23171
rect 37424 23140 38577 23168
rect 37424 23128 37430 23140
rect 38565 23137 38577 23140
rect 38611 23137 38623 23171
rect 38565 23131 38623 23137
rect 36449 23103 36507 23109
rect 36449 23100 36461 23103
rect 36228 23072 36461 23100
rect 36228 23060 36234 23072
rect 36449 23069 36461 23072
rect 36495 23069 36507 23103
rect 36449 23063 36507 23069
rect 36541 23103 36599 23109
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 36633 23103 36691 23109
rect 36633 23069 36645 23103
rect 36679 23069 36691 23103
rect 36633 23063 36691 23069
rect 31444 23004 31754 23032
rect 31444 22992 31450 23004
rect 34514 22992 34520 23044
rect 34572 23032 34578 23044
rect 36648 23032 36676 23063
rect 36814 23060 36820 23112
rect 36872 23060 36878 23112
rect 38749 23103 38807 23109
rect 38749 23069 38761 23103
rect 38795 23069 38807 23103
rect 38749 23063 38807 23069
rect 38764 23032 38792 23063
rect 40218 23060 40224 23112
rect 40276 23100 40282 23112
rect 40773 23103 40831 23109
rect 40773 23100 40785 23103
rect 40276 23072 40785 23100
rect 40276 23060 40282 23072
rect 40773 23069 40785 23072
rect 40819 23069 40831 23103
rect 40773 23063 40831 23069
rect 38838 23032 38844 23044
rect 34572 23004 38844 23032
rect 34572 22992 34578 23004
rect 38838 22992 38844 23004
rect 38896 22992 38902 23044
rect 38933 23035 38991 23041
rect 38933 23001 38945 23035
rect 38979 23032 38991 23035
rect 41018 23035 41076 23041
rect 41018 23032 41030 23035
rect 38979 23004 41030 23032
rect 38979 23001 38991 23004
rect 38933 22995 38991 23001
rect 41018 23001 41030 23004
rect 41064 23001 41076 23035
rect 41018 22995 41076 23001
rect 26069 22967 26127 22973
rect 26069 22964 26081 22967
rect 22204 22936 26081 22964
rect 26069 22933 26081 22936
rect 26115 22933 26127 22967
rect 26069 22927 26127 22933
rect 28350 22924 28356 22976
rect 28408 22964 28414 22976
rect 29086 22964 29092 22976
rect 28408 22936 29092 22964
rect 28408 22924 28414 22936
rect 29086 22924 29092 22936
rect 29144 22924 29150 22976
rect 36173 22967 36231 22973
rect 36173 22933 36185 22967
rect 36219 22964 36231 22967
rect 36814 22964 36820 22976
rect 36219 22936 36820 22964
rect 36219 22933 36231 22936
rect 36173 22927 36231 22933
rect 36814 22924 36820 22936
rect 36872 22924 36878 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 2406 22720 2412 22772
rect 2464 22720 2470 22772
rect 5166 22720 5172 22772
rect 5224 22760 5230 22772
rect 5445 22763 5503 22769
rect 5445 22760 5457 22763
rect 5224 22732 5457 22760
rect 5224 22720 5230 22732
rect 5445 22729 5457 22732
rect 5491 22729 5503 22763
rect 5445 22723 5503 22729
rect 12802 22720 12808 22772
rect 12860 22720 12866 22772
rect 13173 22763 13231 22769
rect 13173 22729 13185 22763
rect 13219 22760 13231 22763
rect 13538 22760 13544 22772
rect 13219 22732 13544 22760
rect 13219 22729 13231 22732
rect 13173 22723 13231 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 18414 22720 18420 22772
rect 18472 22760 18478 22772
rect 18785 22763 18843 22769
rect 18785 22760 18797 22763
rect 18472 22732 18797 22760
rect 18472 22720 18478 22732
rect 18785 22729 18797 22732
rect 18831 22760 18843 22763
rect 18874 22760 18880 22772
rect 18831 22732 18880 22760
rect 18831 22729 18843 22732
rect 18785 22723 18843 22729
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 23750 22720 23756 22772
rect 23808 22720 23814 22772
rect 26050 22720 26056 22772
rect 26108 22760 26114 22772
rect 26145 22763 26203 22769
rect 26145 22760 26157 22763
rect 26108 22732 26157 22760
rect 26108 22720 26114 22732
rect 26145 22729 26157 22732
rect 26191 22729 26203 22763
rect 26145 22723 26203 22729
rect 28442 22720 28448 22772
rect 28500 22760 28506 22772
rect 29549 22763 29607 22769
rect 28500 22732 29500 22760
rect 28500 22720 28506 22732
rect 4332 22695 4390 22701
rect 4332 22661 4344 22695
rect 4378 22692 4390 22695
rect 4430 22692 4436 22704
rect 4378 22664 4436 22692
rect 4378 22661 4390 22664
rect 4332 22655 4390 22661
rect 4430 22652 4436 22664
rect 4488 22652 4494 22704
rect 10778 22692 10784 22704
rect 8036 22664 10784 22692
rect 2317 22627 2375 22633
rect 2317 22593 2329 22627
rect 2363 22624 2375 22627
rect 3050 22624 3056 22636
rect 2363 22596 3056 22624
rect 2363 22593 2375 22596
rect 2317 22587 2375 22593
rect 3050 22584 3056 22596
rect 3108 22584 3114 22636
rect 3234 22584 3240 22636
rect 3292 22584 3298 22636
rect 3602 22584 3608 22636
rect 3660 22624 3666 22636
rect 8036 22633 8064 22664
rect 10778 22652 10784 22664
rect 10836 22652 10842 22704
rect 14366 22652 14372 22704
rect 14424 22692 14430 22704
rect 22186 22692 22192 22704
rect 14424 22664 22192 22692
rect 14424 22652 14430 22664
rect 22186 22652 22192 22664
rect 22244 22652 22250 22704
rect 22388 22664 24624 22692
rect 4065 22627 4123 22633
rect 4065 22624 4077 22627
rect 3660 22596 4077 22624
rect 3660 22584 3666 22596
rect 4065 22593 4077 22596
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 8202 22584 8208 22636
rect 8260 22584 8266 22636
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22624 8355 22627
rect 9030 22624 9036 22636
rect 8343 22596 9036 22624
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 9674 22633 9680 22636
rect 9668 22587 9680 22633
rect 9674 22584 9680 22587
rect 9732 22584 9738 22636
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22624 13047 22627
rect 13078 22624 13084 22636
rect 13035 22596 13084 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 13262 22584 13268 22636
rect 13320 22584 13326 22636
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22624 14979 22627
rect 15010 22624 15016 22636
rect 14967 22596 15016 22624
rect 14967 22593 14979 22596
rect 14921 22587 14979 22593
rect 2590 22516 2596 22568
rect 2648 22556 2654 22568
rect 2958 22556 2964 22568
rect 2648 22528 2964 22556
rect 2648 22516 2654 22528
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 9398 22516 9404 22568
rect 9456 22516 9462 22568
rect 12894 22516 12900 22568
rect 12952 22556 12958 22568
rect 14936 22556 14964 22587
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15188 22627 15246 22633
rect 15188 22593 15200 22627
rect 15234 22624 15246 22627
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 15234 22596 16865 22624
rect 15234 22593 15246 22596
rect 15188 22587 15246 22593
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 17034 22584 17040 22636
rect 17092 22584 17098 22636
rect 17313 22627 17371 22633
rect 17313 22593 17325 22627
rect 17359 22624 17371 22627
rect 17770 22624 17776 22636
rect 17359 22596 17776 22624
rect 17359 22593 17371 22596
rect 17313 22587 17371 22593
rect 17328 22556 17356 22587
rect 17770 22584 17776 22596
rect 17828 22584 17834 22636
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 12952 22528 14964 22556
rect 16316 22528 17356 22556
rect 18708 22556 18736 22587
rect 18874 22584 18880 22636
rect 18932 22584 18938 22636
rect 22278 22584 22284 22636
rect 22336 22624 22342 22636
rect 22388 22633 22416 22664
rect 24596 22636 24624 22664
rect 29178 22652 29184 22704
rect 29236 22652 29242 22704
rect 29381 22695 29439 22701
rect 29381 22692 29393 22695
rect 29288 22664 29393 22692
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 22336 22596 22385 22624
rect 22336 22584 22342 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 22640 22627 22698 22633
rect 22640 22593 22652 22627
rect 22686 22624 22698 22627
rect 23382 22624 23388 22636
rect 22686 22596 23388 22624
rect 22686 22593 22698 22596
rect 22640 22587 22698 22593
rect 23382 22584 23388 22596
rect 23440 22584 23446 22636
rect 24578 22584 24584 22636
rect 24636 22624 24642 22636
rect 25038 22633 25044 22636
rect 24765 22627 24823 22633
rect 24765 22624 24777 22627
rect 24636 22596 24777 22624
rect 24636 22584 24642 22596
rect 24765 22593 24777 22596
rect 24811 22593 24823 22627
rect 24765 22587 24823 22593
rect 25032 22587 25044 22633
rect 25038 22584 25044 22587
rect 25096 22584 25102 22636
rect 19334 22556 19340 22568
rect 18708 22528 19340 22556
rect 12952 22516 12958 22528
rect 8113 22491 8171 22497
rect 8113 22457 8125 22491
rect 8159 22457 8171 22491
rect 8113 22451 8171 22457
rect 1946 22380 1952 22432
rect 2004 22380 2010 22432
rect 3326 22380 3332 22432
rect 3384 22380 3390 22432
rect 6730 22380 6736 22432
rect 6788 22420 6794 22432
rect 7837 22423 7895 22429
rect 7837 22420 7849 22423
rect 6788 22392 7849 22420
rect 6788 22380 6794 22392
rect 7837 22389 7849 22392
rect 7883 22389 7895 22423
rect 8128 22420 8156 22451
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 16316 22497 16344 22528
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 10781 22491 10839 22497
rect 10781 22488 10793 22491
rect 10468 22460 10793 22488
rect 10468 22448 10474 22460
rect 10781 22457 10793 22460
rect 10827 22457 10839 22491
rect 10781 22451 10839 22457
rect 16301 22491 16359 22497
rect 16301 22457 16313 22491
rect 16347 22457 16359 22491
rect 16301 22451 16359 22457
rect 16850 22448 16856 22500
rect 16908 22488 16914 22500
rect 20346 22488 20352 22500
rect 16908 22460 20352 22488
rect 16908 22448 16914 22460
rect 20346 22448 20352 22460
rect 20404 22448 20410 22500
rect 29288 22488 29316 22664
rect 29381 22661 29393 22664
rect 29427 22661 29439 22695
rect 29381 22655 29439 22661
rect 29472 22624 29500 22732
rect 29549 22729 29561 22763
rect 29595 22760 29607 22763
rect 30006 22760 30012 22772
rect 29595 22732 30012 22760
rect 29595 22729 29607 22732
rect 29549 22723 29607 22729
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 31754 22760 31760 22772
rect 31312 22732 31760 22760
rect 31312 22701 31340 22732
rect 31754 22720 31760 22732
rect 31812 22720 31818 22772
rect 31297 22695 31355 22701
rect 31297 22661 31309 22695
rect 31343 22661 31355 22695
rect 31297 22655 31355 22661
rect 31481 22695 31539 22701
rect 31481 22661 31493 22695
rect 31527 22692 31539 22695
rect 35802 22692 35808 22704
rect 31527 22664 35808 22692
rect 31527 22661 31539 22664
rect 31481 22655 31539 22661
rect 31496 22624 31524 22655
rect 35802 22652 35808 22664
rect 35860 22652 35866 22704
rect 29472 22596 31524 22624
rect 28966 22460 29316 22488
rect 10686 22420 10692 22432
rect 8128 22392 10692 22420
rect 7837 22383 7895 22389
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 17221 22423 17279 22429
rect 17221 22420 17233 22423
rect 17000 22392 17233 22420
rect 17000 22380 17006 22392
rect 17221 22389 17233 22392
rect 17267 22389 17279 22423
rect 17221 22383 17279 22389
rect 19702 22380 19708 22432
rect 19760 22420 19766 22432
rect 28966 22420 28994 22460
rect 19760 22392 28994 22420
rect 29365 22423 29423 22429
rect 19760 22380 19766 22392
rect 29365 22389 29377 22423
rect 29411 22420 29423 22423
rect 30190 22420 30196 22432
rect 29411 22392 30196 22420
rect 29411 22389 29423 22392
rect 29365 22383 29423 22389
rect 30190 22380 30196 22392
rect 30248 22420 30254 22432
rect 30558 22420 30564 22432
rect 30248 22392 30564 22420
rect 30248 22380 30254 22392
rect 30558 22380 30564 22392
rect 30616 22420 30622 22432
rect 31481 22423 31539 22429
rect 31481 22420 31493 22423
rect 30616 22392 31493 22420
rect 30616 22380 30622 22392
rect 31481 22389 31493 22392
rect 31527 22389 31539 22423
rect 31481 22383 31539 22389
rect 31665 22423 31723 22429
rect 31665 22389 31677 22423
rect 31711 22420 31723 22423
rect 32306 22420 32312 22432
rect 31711 22392 32312 22420
rect 31711 22389 31723 22392
rect 31665 22383 31723 22389
rect 32306 22380 32312 22392
rect 32364 22380 32370 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 3050 22176 3056 22228
rect 3108 22176 3114 22228
rect 5166 22176 5172 22228
rect 5224 22176 5230 22228
rect 9674 22176 9680 22228
rect 9732 22216 9738 22228
rect 9861 22219 9919 22225
rect 9861 22216 9873 22219
rect 9732 22188 9873 22216
rect 9732 22176 9738 22188
rect 9861 22185 9873 22188
rect 9907 22185 9919 22219
rect 9861 22179 9919 22185
rect 19334 22176 19340 22228
rect 19392 22216 19398 22228
rect 19797 22219 19855 22225
rect 19797 22216 19809 22219
rect 19392 22188 19809 22216
rect 19392 22176 19398 22188
rect 19797 22185 19809 22188
rect 19843 22185 19855 22219
rect 19797 22179 19855 22185
rect 23382 22176 23388 22228
rect 23440 22176 23446 22228
rect 25038 22176 25044 22228
rect 25096 22216 25102 22228
rect 25133 22219 25191 22225
rect 25133 22216 25145 22219
rect 25096 22188 25145 22216
rect 25096 22176 25102 22188
rect 25133 22185 25145 22188
rect 25179 22185 25191 22219
rect 25133 22179 25191 22185
rect 27522 22176 27528 22228
rect 27580 22176 27586 22228
rect 29178 22176 29184 22228
rect 29236 22216 29242 22228
rect 30282 22216 30288 22228
rect 29236 22188 30288 22216
rect 29236 22176 29242 22188
rect 30282 22176 30288 22188
rect 30340 22176 30346 22228
rect 30834 22176 30840 22228
rect 30892 22216 30898 22228
rect 31478 22216 31484 22228
rect 30892 22188 31484 22216
rect 30892 22176 30898 22188
rect 31478 22176 31484 22188
rect 31536 22176 31542 22228
rect 37458 22176 37464 22228
rect 37516 22216 37522 22228
rect 37921 22219 37979 22225
rect 37921 22216 37933 22219
rect 37516 22188 37933 22216
rect 37516 22176 37522 22188
rect 37921 22185 37933 22188
rect 37967 22185 37979 22219
rect 37921 22179 37979 22185
rect 3068 22080 3096 22176
rect 4724 22120 5120 22148
rect 4724 22080 4752 22120
rect 3068 22052 4752 22080
rect 4798 22040 4804 22092
rect 4856 22080 4862 22092
rect 4985 22083 5043 22089
rect 4985 22080 4997 22083
rect 4856 22052 4997 22080
rect 4856 22040 4862 22052
rect 4985 22049 4997 22052
rect 5031 22049 5043 22083
rect 5092 22080 5120 22120
rect 16758 22108 16764 22160
rect 16816 22148 16822 22160
rect 19702 22148 19708 22160
rect 16816 22120 19708 22148
rect 16816 22108 16822 22120
rect 19702 22108 19708 22120
rect 19760 22108 19766 22160
rect 19981 22151 20039 22157
rect 19981 22117 19993 22151
rect 20027 22148 20039 22151
rect 20070 22148 20076 22160
rect 20027 22120 20076 22148
rect 20027 22117 20039 22120
rect 19981 22111 20039 22117
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 27540 22148 27568 22176
rect 30650 22148 30656 22160
rect 27540 22120 30656 22148
rect 30650 22108 30656 22120
rect 30708 22108 30714 22160
rect 13170 22080 13176 22092
rect 5092 22052 5212 22080
rect 4985 22043 5043 22049
rect 5184 22024 5212 22052
rect 6886 22052 13176 22080
rect 1670 21972 1676 22024
rect 1728 21972 1734 22024
rect 1946 22021 1952 22024
rect 1940 22012 1952 22021
rect 1907 21984 1952 22012
rect 1940 21975 1952 21984
rect 1946 21972 1952 21975
rect 2004 21972 2010 22024
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4295 21984 5120 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 934 21904 940 21956
rect 992 21944 998 21956
rect 4065 21947 4123 21953
rect 4065 21944 4077 21947
rect 992 21916 4077 21944
rect 992 21904 998 21916
rect 4065 21913 4077 21916
rect 4111 21913 4123 21947
rect 4065 21907 4123 21913
rect 4893 21947 4951 21953
rect 4893 21913 4905 21947
rect 4939 21944 4951 21947
rect 4982 21944 4988 21956
rect 4939 21916 4988 21944
rect 4939 21913 4951 21916
rect 4893 21907 4951 21913
rect 4982 21904 4988 21916
rect 5040 21904 5046 21956
rect 5092 21944 5120 21984
rect 5166 21972 5172 22024
rect 5224 21972 5230 22024
rect 5258 21972 5264 22024
rect 5316 22012 5322 22024
rect 6886 22012 6914 22052
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 13262 22040 13268 22092
rect 13320 22080 13326 22092
rect 18785 22083 18843 22089
rect 13320 22052 14780 22080
rect 13320 22040 13326 22052
rect 5316 21984 6914 22012
rect 5316 21972 5322 21984
rect 10042 21972 10048 22024
rect 10100 21972 10106 22024
rect 10318 21972 10324 22024
rect 10376 21972 10382 22024
rect 14752 22021 14780 22052
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 19889 22083 19947 22089
rect 19889 22080 19901 22083
rect 18831 22052 19901 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 19889 22049 19901 22052
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 25240 22052 25636 22080
rect 25240 22024 25268 22052
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 14737 22015 14795 22021
rect 14737 21981 14749 22015
rect 14783 21981 14795 22015
rect 14737 21975 14795 21981
rect 11882 21944 11888 21956
rect 5092 21916 11888 21944
rect 11882 21904 11888 21916
rect 11940 21904 11946 21956
rect 14090 21904 14096 21956
rect 14148 21944 14154 21956
rect 14476 21944 14504 21975
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 18693 22015 18751 22021
rect 18693 22012 18705 22015
rect 17736 21984 18705 22012
rect 17736 21972 17742 21984
rect 18693 21981 18705 21984
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 19702 21972 19708 22024
rect 19760 21972 19766 22024
rect 20162 21972 20168 22024
rect 20220 21972 20226 22024
rect 21453 22015 21511 22021
rect 21453 21981 21465 22015
rect 21499 22012 21511 22015
rect 22278 22012 22284 22024
rect 21499 21984 22284 22012
rect 21499 21981 21511 21984
rect 21453 21975 21511 21981
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 23474 21972 23480 22024
rect 23532 22012 23538 22024
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 23532 21984 23581 22012
rect 23532 21972 23538 21984
rect 23569 21981 23581 21984
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 23750 21972 23756 22024
rect 23808 21972 23814 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 22012 23903 22015
rect 25222 22012 25228 22024
rect 23891 21984 25228 22012
rect 23891 21981 23903 21984
rect 23845 21975 23903 21981
rect 21720 21947 21778 21953
rect 14148 21916 14412 21944
rect 14476 21916 19564 21944
rect 14148 21904 14154 21916
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 5258 21876 5264 21888
rect 2280 21848 5264 21876
rect 2280 21836 2286 21848
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 5353 21879 5411 21885
rect 5353 21845 5365 21879
rect 5399 21876 5411 21879
rect 6454 21876 6460 21888
rect 5399 21848 6460 21876
rect 5399 21845 5411 21848
rect 5353 21839 5411 21845
rect 6454 21836 6460 21848
rect 6512 21836 6518 21888
rect 10229 21879 10287 21885
rect 10229 21845 10241 21879
rect 10275 21876 10287 21879
rect 10410 21876 10416 21888
rect 10275 21848 10416 21876
rect 10275 21845 10287 21848
rect 10229 21839 10287 21845
rect 10410 21836 10416 21848
rect 10468 21836 10474 21888
rect 14274 21836 14280 21888
rect 14332 21836 14338 21888
rect 14384 21876 14412 21916
rect 14645 21879 14703 21885
rect 14645 21876 14657 21879
rect 14384 21848 14657 21876
rect 14645 21845 14657 21848
rect 14691 21845 14703 21879
rect 14645 21839 14703 21845
rect 18046 21836 18052 21888
rect 18104 21876 18110 21888
rect 19429 21879 19487 21885
rect 19429 21876 19441 21879
rect 18104 21848 19441 21876
rect 18104 21836 18110 21848
rect 19429 21845 19441 21848
rect 19475 21845 19487 21879
rect 19536 21876 19564 21916
rect 21720 21913 21732 21947
rect 21766 21944 21778 21947
rect 22186 21944 22192 21956
rect 21766 21916 22192 21944
rect 21766 21913 21778 21916
rect 21720 21907 21778 21913
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 23860 21944 23888 21975
rect 25222 21972 25228 21984
rect 25280 21972 25286 22024
rect 25314 21972 25320 22024
rect 25372 21972 25378 22024
rect 25608 22021 25636 22052
rect 26326 22040 26332 22092
rect 26384 22080 26390 22092
rect 27522 22080 27528 22092
rect 26384 22052 27528 22080
rect 26384 22040 26390 22052
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 35345 22083 35403 22089
rect 29932 22052 30972 22080
rect 29932 22021 29960 22052
rect 25593 22015 25651 22021
rect 25593 21981 25605 22015
rect 25639 21981 25651 22015
rect 25593 21975 25651 21981
rect 29917 22015 29975 22021
rect 29917 21981 29929 22015
rect 29963 21981 29975 22015
rect 29917 21975 29975 21981
rect 30190 21972 30196 22024
rect 30248 21972 30254 22024
rect 22296 21916 23888 21944
rect 25501 21947 25559 21953
rect 22296 21888 22324 21916
rect 25501 21913 25513 21947
rect 25547 21944 25559 21947
rect 26050 21944 26056 21956
rect 25547 21916 26056 21944
rect 25547 21913 25559 21916
rect 25501 21907 25559 21913
rect 26050 21904 26056 21916
rect 26108 21904 26114 21956
rect 30653 21947 30711 21953
rect 30653 21913 30665 21947
rect 30699 21944 30711 21947
rect 30742 21944 30748 21956
rect 30699 21916 30748 21944
rect 30699 21913 30711 21916
rect 30653 21907 30711 21913
rect 30742 21904 30748 21916
rect 30800 21904 30806 21956
rect 20714 21876 20720 21888
rect 19536 21848 20720 21876
rect 19429 21839 19487 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 22278 21836 22284 21888
rect 22336 21836 22342 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 22830 21876 22836 21888
rect 22612 21848 22836 21876
rect 22612 21836 22618 21848
rect 22830 21836 22836 21848
rect 22888 21836 22894 21888
rect 29730 21836 29736 21888
rect 29788 21836 29794 21888
rect 30098 21836 30104 21888
rect 30156 21836 30162 21888
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 30853 21879 30911 21885
rect 30853 21876 30865 21879
rect 30524 21848 30865 21876
rect 30524 21836 30530 21848
rect 30853 21845 30865 21848
rect 30899 21845 30911 21879
rect 30944 21876 30972 22052
rect 35345 22049 35357 22083
rect 35391 22080 35403 22083
rect 35802 22080 35808 22092
rect 35391 22052 35808 22080
rect 35391 22049 35403 22052
rect 35345 22043 35403 22049
rect 35802 22040 35808 22052
rect 35860 22040 35866 22092
rect 36538 22040 36544 22092
rect 36596 22040 36602 22092
rect 36814 22040 36820 22092
rect 36872 22040 36878 22092
rect 32950 21972 32956 22024
rect 33008 21972 33014 22024
rect 40218 21972 40224 22024
rect 40276 21972 40282 22024
rect 33220 21947 33278 21953
rect 33220 21913 33232 21947
rect 33266 21944 33278 21947
rect 33318 21944 33324 21956
rect 33266 21916 33324 21944
rect 33266 21913 33278 21916
rect 33220 21907 33278 21913
rect 33318 21904 33324 21916
rect 33376 21904 33382 21956
rect 34977 21947 35035 21953
rect 34977 21944 34989 21947
rect 34348 21916 34989 21944
rect 34348 21888 34376 21916
rect 34977 21913 34989 21916
rect 35023 21913 35035 21947
rect 34977 21907 35035 21913
rect 35161 21947 35219 21953
rect 35161 21913 35173 21947
rect 35207 21913 35219 21947
rect 35161 21907 35219 21913
rect 40488 21947 40546 21953
rect 40488 21913 40500 21947
rect 40534 21944 40546 21947
rect 40586 21944 40592 21956
rect 40534 21916 40592 21944
rect 40534 21913 40546 21916
rect 40488 21907 40546 21913
rect 31021 21879 31079 21885
rect 31021 21876 31033 21879
rect 30944 21848 31033 21876
rect 30853 21839 30911 21845
rect 31021 21845 31033 21848
rect 31067 21876 31079 21879
rect 33594 21876 33600 21888
rect 31067 21848 33600 21876
rect 31067 21845 31079 21848
rect 31021 21839 31079 21845
rect 33594 21836 33600 21848
rect 33652 21836 33658 21888
rect 34330 21836 34336 21888
rect 34388 21836 34394 21888
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 35176 21876 35204 21907
rect 40586 21904 40592 21916
rect 40644 21904 40650 21956
rect 34848 21848 35204 21876
rect 34848 21836 34854 21848
rect 40954 21836 40960 21888
rect 41012 21876 41018 21888
rect 41601 21879 41659 21885
rect 41601 21876 41613 21879
rect 41012 21848 41613 21876
rect 41012 21836 41018 21848
rect 41601 21845 41613 21848
rect 41647 21845 41659 21879
rect 41601 21839 41659 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 934 21632 940 21684
rect 992 21672 998 21684
rect 3234 21672 3240 21684
rect 992 21644 3240 21672
rect 992 21632 998 21644
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 9493 21675 9551 21681
rect 9493 21672 9505 21675
rect 4028 21644 9505 21672
rect 4028 21632 4034 21644
rect 9493 21641 9505 21644
rect 9539 21672 9551 21675
rect 9674 21672 9680 21684
rect 9539 21644 9680 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 32858 21672 32864 21684
rect 11440 21644 32864 21672
rect 8478 21604 8484 21616
rect 1596 21576 8484 21604
rect 1596 21545 1624 21576
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 1581 21539 1639 21545
rect 1581 21505 1593 21539
rect 1627 21505 1639 21539
rect 1581 21499 1639 21505
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 4062 21536 4068 21548
rect 2547 21508 4068 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 4062 21496 4068 21508
rect 4120 21496 4126 21548
rect 5074 21496 5080 21548
rect 5132 21496 5138 21548
rect 5534 21496 5540 21548
rect 5592 21536 5598 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 5592 21508 6561 21536
rect 5592 21496 5598 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 7009 21539 7067 21545
rect 7009 21536 7021 21539
rect 6549 21499 6607 21505
rect 6656 21508 7021 21536
rect 1026 21428 1032 21480
rect 1084 21468 1090 21480
rect 1765 21471 1823 21477
rect 1765 21468 1777 21471
rect 1084 21440 1777 21468
rect 1084 21428 1090 21440
rect 1765 21437 1777 21440
rect 1811 21437 1823 21471
rect 1765 21431 1823 21437
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 934 21360 940 21412
rect 992 21400 998 21412
rect 2700 21400 2728 21431
rect 3418 21428 3424 21480
rect 3476 21468 3482 21480
rect 5169 21471 5227 21477
rect 5169 21468 5181 21471
rect 3476 21440 5181 21468
rect 3476 21428 3482 21440
rect 5169 21437 5181 21440
rect 5215 21468 5227 21471
rect 6656 21468 6684 21508
rect 7009 21505 7021 21508
rect 7055 21505 7067 21539
rect 7009 21499 7067 21505
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21536 9367 21539
rect 9490 21536 9496 21548
rect 9355 21508 9496 21536
rect 9355 21505 9367 21508
rect 9309 21499 9367 21505
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 9582 21496 9588 21548
rect 9640 21496 9646 21548
rect 5215 21440 6684 21468
rect 6917 21471 6975 21477
rect 5215 21437 5227 21440
rect 5169 21431 5227 21437
rect 6917 21437 6929 21471
rect 6963 21468 6975 21471
rect 7190 21468 7196 21480
rect 6963 21440 7196 21468
rect 6963 21437 6975 21440
rect 6917 21431 6975 21437
rect 7190 21428 7196 21440
rect 7248 21428 7254 21480
rect 11440 21400 11468 21644
rect 32858 21632 32864 21644
rect 32916 21632 32922 21684
rect 33318 21632 33324 21684
rect 33376 21632 33382 21684
rect 33689 21675 33747 21681
rect 33689 21641 33701 21675
rect 33735 21672 33747 21675
rect 34330 21672 34336 21684
rect 33735 21644 34336 21672
rect 33735 21641 33747 21644
rect 33689 21635 33747 21641
rect 34330 21632 34336 21644
rect 34388 21672 34394 21684
rect 34698 21672 34704 21684
rect 34388 21644 34704 21672
rect 34388 21632 34394 21644
rect 34698 21632 34704 21644
rect 34756 21632 34762 21684
rect 37829 21675 37887 21681
rect 37829 21641 37841 21675
rect 37875 21641 37887 21675
rect 37829 21635 37887 21641
rect 11882 21564 11888 21616
rect 11940 21564 11946 21616
rect 13164 21607 13222 21613
rect 13164 21573 13176 21607
rect 13210 21604 13222 21607
rect 14274 21604 14280 21616
rect 13210 21576 14280 21604
rect 13210 21573 13222 21576
rect 13164 21567 13222 21573
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 15930 21564 15936 21616
rect 15988 21604 15994 21616
rect 17405 21607 17463 21613
rect 17405 21604 17417 21607
rect 15988 21576 17417 21604
rect 15988 21564 15994 21576
rect 17405 21573 17417 21576
rect 17451 21573 17463 21607
rect 17405 21567 17463 21573
rect 17621 21607 17679 21613
rect 17621 21573 17633 21607
rect 17667 21604 17679 21607
rect 17954 21604 17960 21616
rect 17667 21576 17960 21604
rect 17667 21573 17679 21576
rect 17621 21567 17679 21573
rect 11514 21496 11520 21548
rect 11572 21536 11578 21548
rect 11977 21539 12035 21545
rect 11977 21536 11989 21539
rect 11572 21508 11989 21536
rect 11572 21496 11578 21508
rect 11977 21505 11989 21508
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21536 12955 21539
rect 12986 21536 12992 21548
rect 12943 21508 12992 21536
rect 12943 21505 12955 21508
rect 12897 21499 12955 21505
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 17420 21468 17448 21567
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 19429 21607 19487 21613
rect 19429 21573 19441 21607
rect 19475 21604 19487 21607
rect 20162 21604 20168 21616
rect 19475 21576 20168 21604
rect 19475 21573 19487 21576
rect 19429 21567 19487 21573
rect 20162 21564 20168 21576
rect 20220 21564 20226 21616
rect 22094 21564 22100 21616
rect 22152 21564 22158 21616
rect 22465 21607 22523 21613
rect 22465 21573 22477 21607
rect 22511 21604 22523 21607
rect 26326 21604 26332 21616
rect 22511 21576 26332 21604
rect 22511 21573 22523 21576
rect 22465 21567 22523 21573
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 20346 21536 20352 21548
rect 19383 21508 20352 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 22480 21536 22508 21567
rect 26326 21564 26332 21576
rect 26384 21564 26390 21616
rect 28896 21607 28954 21613
rect 28896 21573 28908 21607
rect 28942 21604 28954 21607
rect 29730 21604 29736 21616
rect 28942 21576 29736 21604
rect 28942 21573 28954 21576
rect 28896 21567 28954 21573
rect 29730 21564 29736 21576
rect 29788 21564 29794 21616
rect 30834 21564 30840 21616
rect 30892 21604 30898 21616
rect 34514 21604 34520 21616
rect 30892 21576 34520 21604
rect 30892 21564 30898 21576
rect 34514 21564 34520 21576
rect 34572 21564 34578 21616
rect 37461 21607 37519 21613
rect 37461 21573 37473 21607
rect 37507 21573 37519 21607
rect 37461 21567 37519 21573
rect 21131 21508 22508 21536
rect 25961 21539 26019 21545
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 19978 21468 19984 21480
rect 17420 21440 19984 21468
rect 19978 21428 19984 21440
rect 20036 21468 20042 21480
rect 20438 21468 20444 21480
rect 20036 21440 20444 21468
rect 20036 21428 20042 21440
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 992 21372 2728 21400
rect 2792 21372 11468 21400
rect 11532 21372 12204 21400
rect 992 21360 998 21372
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 2792 21332 2820 21372
rect 1912 21304 2820 21332
rect 1912 21292 1918 21304
rect 5166 21292 5172 21344
rect 5224 21292 5230 21344
rect 5442 21292 5448 21344
rect 5500 21292 5506 21344
rect 6638 21292 6644 21344
rect 6696 21292 6702 21344
rect 7190 21292 7196 21344
rect 7248 21292 7254 21344
rect 8570 21292 8576 21344
rect 8628 21332 8634 21344
rect 9125 21335 9183 21341
rect 9125 21332 9137 21335
rect 8628 21304 9137 21332
rect 8628 21292 8634 21304
rect 9125 21301 9137 21304
rect 9171 21301 9183 21335
rect 9125 21295 9183 21301
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11532 21332 11560 21372
rect 11112 21304 11560 21332
rect 11112 21292 11118 21304
rect 11698 21292 11704 21344
rect 11756 21292 11762 21344
rect 12176 21341 12204 21372
rect 14090 21360 14096 21412
rect 14148 21400 14154 21412
rect 14277 21403 14335 21409
rect 14277 21400 14289 21403
rect 14148 21372 14289 21400
rect 14148 21360 14154 21372
rect 14277 21369 14289 21372
rect 14323 21369 14335 21403
rect 18506 21400 18512 21412
rect 14277 21363 14335 21369
rect 17604 21372 18512 21400
rect 17604 21341 17632 21372
rect 18506 21360 18512 21372
rect 18564 21360 18570 21412
rect 12161 21335 12219 21341
rect 12161 21301 12173 21335
rect 12207 21301 12219 21335
rect 12161 21295 12219 21301
rect 17589 21335 17647 21341
rect 17589 21301 17601 21335
rect 17635 21301 17647 21335
rect 17589 21295 17647 21301
rect 17770 21292 17776 21344
rect 17828 21292 17834 21344
rect 20990 21292 20996 21344
rect 21048 21332 21054 21344
rect 21177 21335 21235 21341
rect 21177 21332 21189 21335
rect 21048 21304 21189 21332
rect 21048 21292 21054 21304
rect 21177 21301 21189 21304
rect 21223 21301 21235 21335
rect 21177 21295 21235 21301
rect 21634 21292 21640 21344
rect 21692 21332 21698 21344
rect 22066 21332 22094 21508
rect 25961 21505 25973 21539
rect 26007 21536 26019 21539
rect 27154 21536 27160 21548
rect 26007 21508 27160 21536
rect 26007 21505 26019 21508
rect 25961 21499 26019 21505
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 30650 21496 30656 21548
rect 30708 21496 30714 21548
rect 33502 21496 33508 21548
rect 33560 21496 33566 21548
rect 33778 21542 33784 21548
rect 33612 21514 33784 21542
rect 25866 21428 25872 21480
rect 25924 21468 25930 21480
rect 26053 21471 26111 21477
rect 26053 21468 26065 21471
rect 25924 21440 26065 21468
rect 25924 21428 25930 21440
rect 26053 21437 26065 21440
rect 26099 21437 26111 21471
rect 26053 21431 26111 21437
rect 26142 21428 26148 21480
rect 26200 21428 26206 21480
rect 26234 21428 26240 21480
rect 26292 21428 26298 21480
rect 27338 21428 27344 21480
rect 27396 21428 27402 21480
rect 27433 21471 27491 21477
rect 27433 21437 27445 21471
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 27062 21360 27068 21412
rect 27120 21400 27126 21412
rect 27448 21400 27476 21431
rect 27522 21428 27528 21480
rect 27580 21428 27586 21480
rect 27614 21428 27620 21480
rect 27672 21428 27678 21480
rect 28626 21428 28632 21480
rect 28684 21428 28690 21480
rect 27120 21372 27476 21400
rect 30668 21400 30696 21496
rect 30834 21428 30840 21480
rect 30892 21428 30898 21480
rect 31202 21428 31208 21480
rect 31260 21468 31266 21480
rect 33612 21468 33640 21514
rect 33778 21496 33784 21514
rect 33836 21496 33842 21548
rect 33870 21496 33876 21548
rect 33928 21536 33934 21548
rect 34241 21539 34299 21545
rect 34241 21536 34253 21539
rect 33928 21508 34253 21536
rect 33928 21496 33934 21508
rect 34241 21505 34253 21508
rect 34287 21505 34299 21539
rect 34241 21499 34299 21505
rect 34422 21496 34428 21548
rect 34480 21536 34486 21548
rect 37366 21536 37372 21548
rect 34480 21508 37372 21536
rect 34480 21496 34486 21508
rect 37366 21496 37372 21508
rect 37424 21496 37430 21548
rect 31260 21440 33640 21468
rect 31260 21428 31266 21440
rect 34330 21428 34336 21480
rect 34388 21428 34394 21480
rect 37476 21400 37504 21567
rect 37550 21564 37556 21616
rect 37608 21604 37614 21616
rect 37661 21607 37719 21613
rect 37661 21604 37673 21607
rect 37608 21576 37673 21604
rect 37608 21564 37614 21576
rect 37661 21573 37673 21576
rect 37707 21573 37719 21607
rect 37661 21567 37719 21573
rect 37844 21536 37872 21635
rect 40586 21632 40592 21684
rect 40644 21632 40650 21684
rect 40954 21632 40960 21684
rect 41012 21632 41018 21684
rect 41693 21607 41751 21613
rect 41693 21604 41705 21607
rect 40788 21576 41705 21604
rect 40788 21545 40816 21576
rect 41693 21573 41705 21576
rect 41739 21573 41751 21607
rect 41693 21567 41751 21573
rect 40773 21539 40831 21545
rect 40773 21536 40785 21539
rect 37844 21508 40785 21536
rect 40773 21505 40785 21508
rect 40819 21505 40831 21539
rect 41049 21539 41107 21545
rect 41049 21536 41061 21539
rect 40773 21499 40831 21505
rect 41033 21505 41061 21536
rect 41095 21536 41107 21539
rect 41509 21539 41567 21545
rect 41095 21508 41460 21536
rect 41095 21505 41107 21508
rect 41033 21499 41107 21505
rect 40402 21428 40408 21480
rect 40460 21468 40466 21480
rect 41033 21468 41061 21499
rect 40460 21440 41061 21468
rect 41432 21468 41460 21508
rect 41509 21505 41521 21539
rect 41555 21536 41567 21539
rect 45186 21536 45192 21548
rect 41555 21508 45192 21536
rect 41555 21505 41567 21508
rect 41509 21499 41567 21505
rect 45186 21496 45192 21508
rect 45244 21496 45250 21548
rect 45830 21468 45836 21480
rect 41432 21440 45836 21468
rect 40460 21428 40466 21440
rect 45830 21428 45836 21440
rect 45888 21428 45894 21480
rect 30668 21372 37504 21400
rect 27120 21360 27126 21372
rect 21692 21304 22094 21332
rect 21692 21292 21698 21304
rect 25774 21292 25780 21344
rect 25832 21292 25838 21344
rect 25958 21292 25964 21344
rect 26016 21332 26022 21344
rect 27157 21335 27215 21341
rect 27157 21332 27169 21335
rect 26016 21304 27169 21332
rect 26016 21292 26022 21304
rect 27157 21301 27169 21304
rect 27203 21301 27215 21335
rect 27157 21295 27215 21301
rect 28534 21292 28540 21344
rect 28592 21332 28598 21344
rect 30009 21335 30067 21341
rect 30009 21332 30021 21335
rect 28592 21304 30021 21332
rect 28592 21292 28598 21304
rect 30009 21301 30021 21304
rect 30055 21332 30067 21335
rect 30098 21332 30104 21344
rect 30055 21304 30104 21332
rect 30055 21301 30067 21304
rect 30009 21295 30067 21301
rect 30098 21292 30104 21304
rect 30156 21292 30162 21344
rect 32858 21292 32864 21344
rect 32916 21332 32922 21344
rect 37645 21335 37703 21341
rect 37645 21332 37657 21335
rect 32916 21304 37657 21332
rect 32916 21292 32922 21304
rect 37645 21301 37657 21304
rect 37691 21332 37703 21335
rect 38105 21335 38163 21341
rect 38105 21332 38117 21335
rect 37691 21304 38117 21332
rect 37691 21301 37703 21304
rect 37645 21295 37703 21301
rect 38105 21301 38117 21304
rect 38151 21301 38163 21335
rect 38105 21295 38163 21301
rect 41230 21292 41236 21344
rect 41288 21332 41294 21344
rect 41877 21335 41935 21341
rect 41877 21332 41889 21335
rect 41288 21304 41889 21332
rect 41288 21292 41294 21304
rect 41877 21301 41889 21304
rect 41923 21301 41935 21335
rect 41877 21295 41935 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 7742 21088 7748 21140
rect 7800 21088 7806 21140
rect 10042 21088 10048 21140
rect 10100 21128 10106 21140
rect 10100 21100 11560 21128
rect 10100 21088 10106 21100
rect 11532 21060 11560 21100
rect 11974 21088 11980 21140
rect 12032 21088 12038 21140
rect 17954 21088 17960 21140
rect 18012 21088 18018 21140
rect 18506 21088 18512 21140
rect 18564 21088 18570 21140
rect 22186 21088 22192 21140
rect 22244 21088 22250 21140
rect 23474 21088 23480 21140
rect 23532 21088 23538 21140
rect 27522 21088 27528 21140
rect 27580 21128 27586 21140
rect 34333 21131 34391 21137
rect 27580 21100 34284 21128
rect 27580 21088 27586 21100
rect 25774 21060 25780 21072
rect 11532 21032 25780 21060
rect 25774 21020 25780 21032
rect 25832 21020 25838 21072
rect 27246 21020 27252 21072
rect 27304 21060 27310 21072
rect 30193 21063 30251 21069
rect 30193 21060 30205 21063
rect 27304 21032 30205 21060
rect 27304 21020 27310 21032
rect 30193 21029 30205 21032
rect 30239 21029 30251 21063
rect 30193 21023 30251 21029
rect 30558 21020 30564 21072
rect 30616 21020 30622 21072
rect 31202 21020 31208 21072
rect 31260 21020 31266 21072
rect 34256 21060 34284 21100
rect 34333 21097 34345 21131
rect 34379 21128 34391 21131
rect 34790 21128 34796 21140
rect 34379 21100 34796 21128
rect 34379 21097 34391 21100
rect 34333 21091 34391 21097
rect 34790 21088 34796 21100
rect 34848 21088 34854 21140
rect 40954 21128 40960 21140
rect 36648 21100 40960 21128
rect 36648 21060 36676 21100
rect 40954 21088 40960 21100
rect 41012 21088 41018 21140
rect 44545 21131 44603 21137
rect 44545 21097 44557 21131
rect 44591 21128 44603 21131
rect 44591 21100 45140 21128
rect 44591 21097 44603 21100
rect 44545 21091 44603 21097
rect 34256 21032 36676 21060
rect 42337 21063 42395 21069
rect 42337 21029 42349 21063
rect 42383 21060 42395 21063
rect 43438 21060 43444 21072
rect 42383 21032 43444 21060
rect 42383 21029 42395 21032
rect 42337 21023 42395 21029
rect 43438 21020 43444 21032
rect 43496 21060 43502 21072
rect 43496 21032 44680 21060
rect 43496 21020 43502 21032
rect 2590 20952 2596 21004
rect 2648 20952 2654 21004
rect 21729 20995 21787 21001
rect 16040 20964 21220 20992
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 1728 20896 6377 20924
rect 1728 20884 1734 20896
rect 6365 20893 6377 20896
rect 6411 20924 6423 20927
rect 9398 20924 9404 20936
rect 6411 20896 9404 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 9398 20884 9404 20896
rect 9456 20924 9462 20936
rect 9861 20927 9919 20933
rect 9861 20924 9873 20927
rect 9456 20896 9873 20924
rect 9456 20884 9462 20896
rect 9861 20893 9873 20896
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 10597 20927 10655 20933
rect 10597 20893 10609 20927
rect 10643 20924 10655 20927
rect 12986 20924 12992 20936
rect 10643 20896 12992 20924
rect 10643 20893 10655 20896
rect 10597 20887 10655 20893
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 13170 20884 13176 20936
rect 13228 20924 13234 20936
rect 16040 20924 16068 20964
rect 13228 20896 16068 20924
rect 17589 20927 17647 20933
rect 13228 20884 13234 20896
rect 17589 20893 17601 20927
rect 17635 20924 17647 20927
rect 18414 20924 18420 20936
rect 17635 20896 18420 20924
rect 17635 20893 17647 20896
rect 17589 20887 17647 20893
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20893 18659 20927
rect 18601 20887 18659 20893
rect 2409 20859 2467 20865
rect 2409 20825 2421 20859
rect 2455 20856 2467 20859
rect 3326 20856 3332 20868
rect 2455 20828 3332 20856
rect 2455 20825 2467 20828
rect 2409 20819 2467 20825
rect 3326 20816 3332 20828
rect 3384 20816 3390 20868
rect 6638 20865 6644 20868
rect 6632 20819 6644 20865
rect 6638 20816 6644 20819
rect 6696 20816 6702 20868
rect 9122 20816 9128 20868
rect 9180 20816 9186 20868
rect 10864 20859 10922 20865
rect 10864 20825 10876 20859
rect 10910 20856 10922 20859
rect 12342 20856 12348 20868
rect 10910 20828 12348 20856
rect 10910 20825 10922 20828
rect 10864 20819 10922 20825
rect 12342 20816 12348 20828
rect 12400 20816 12406 20868
rect 15102 20816 15108 20868
rect 15160 20856 15166 20868
rect 15197 20859 15255 20865
rect 15197 20856 15209 20859
rect 15160 20828 15209 20856
rect 15160 20816 15166 20828
rect 15197 20825 15209 20828
rect 15243 20825 15255 20859
rect 15197 20819 15255 20825
rect 15286 20816 15292 20868
rect 15344 20856 15350 20868
rect 15933 20859 15991 20865
rect 15933 20856 15945 20859
rect 15344 20828 15945 20856
rect 15344 20816 15350 20828
rect 15933 20825 15945 20828
rect 15979 20825 15991 20859
rect 15933 20819 15991 20825
rect 17678 20816 17684 20868
rect 17736 20856 17742 20868
rect 17773 20859 17831 20865
rect 17773 20856 17785 20859
rect 17736 20828 17785 20856
rect 17736 20816 17742 20828
rect 17773 20825 17785 20828
rect 17819 20856 17831 20859
rect 18616 20856 18644 20887
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 20990 20924 20996 20936
rect 19300 20896 20996 20924
rect 19300 20884 19306 20896
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21192 20933 21220 20964
rect 21729 20961 21741 20995
rect 21775 20992 21787 20995
rect 21775 20964 23152 20992
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 21269 20927 21327 20933
rect 21269 20893 21281 20927
rect 21315 20924 21327 20927
rect 21358 20924 21364 20936
rect 21315 20896 21364 20924
rect 21315 20893 21327 20896
rect 21269 20887 21327 20893
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 22554 20884 22560 20936
rect 22612 20884 22618 20936
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 22664 20856 22692 20887
rect 17819 20828 18644 20856
rect 22066 20828 22692 20856
rect 17819 20825 17831 20828
rect 17773 20819 17831 20825
rect 1949 20791 2007 20797
rect 1949 20757 1961 20791
rect 1995 20788 2007 20791
rect 2222 20788 2228 20800
rect 1995 20760 2228 20788
rect 1995 20757 2007 20760
rect 1949 20751 2007 20757
rect 2222 20748 2228 20760
rect 2280 20748 2286 20800
rect 2317 20791 2375 20797
rect 2317 20757 2329 20791
rect 2363 20788 2375 20791
rect 3418 20788 3424 20800
rect 2363 20760 3424 20788
rect 2363 20757 2375 20760
rect 2317 20751 2375 20757
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 9582 20748 9588 20800
rect 9640 20788 9646 20800
rect 12434 20788 12440 20800
rect 9640 20760 12440 20788
rect 9640 20748 9646 20760
rect 12434 20748 12440 20760
rect 12492 20788 12498 20800
rect 13262 20788 13268 20800
rect 12492 20760 13268 20788
rect 12492 20748 12498 20760
rect 13262 20748 13268 20760
rect 13320 20748 13326 20800
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 22066 20788 22094 20828
rect 18656 20760 22094 20788
rect 23124 20788 23152 20964
rect 23198 20952 23204 21004
rect 23256 20992 23262 21004
rect 23845 20995 23903 21001
rect 23845 20992 23857 20995
rect 23256 20964 23857 20992
rect 23256 20952 23262 20964
rect 23845 20961 23857 20964
rect 23891 20961 23903 20995
rect 23845 20955 23903 20961
rect 25958 20952 25964 21004
rect 26016 20952 26022 21004
rect 27157 20995 27215 21001
rect 27157 20961 27169 20995
rect 27203 20992 27215 20995
rect 28534 20992 28540 21004
rect 27203 20964 28540 20992
rect 27203 20961 27215 20964
rect 27157 20955 27215 20961
rect 28534 20952 28540 20964
rect 28592 20952 28598 21004
rect 28626 20952 28632 21004
rect 28684 20992 28690 21004
rect 30926 20992 30932 21004
rect 28684 20964 30932 20992
rect 28684 20952 28690 20964
rect 30926 20952 30932 20964
rect 30984 20992 30990 21004
rect 32950 20992 32956 21004
rect 30984 20964 32956 20992
rect 30984 20952 30990 20964
rect 32950 20952 32956 20964
rect 33008 20952 33014 21004
rect 40218 20952 40224 21004
rect 40276 20992 40282 21004
rect 40957 20995 41015 21001
rect 40957 20992 40969 20995
rect 40276 20964 40969 20992
rect 40276 20952 40282 20964
rect 40957 20961 40969 20964
rect 41003 20961 41015 20995
rect 40957 20955 41015 20961
rect 23658 20884 23664 20936
rect 23716 20884 23722 20936
rect 23750 20884 23756 20936
rect 23808 20884 23814 20936
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20893 23995 20927
rect 23937 20887 23995 20893
rect 23566 20816 23572 20868
rect 23624 20856 23630 20868
rect 23952 20856 23980 20887
rect 26050 20884 26056 20936
rect 26108 20884 26114 20936
rect 26142 20884 26148 20936
rect 26200 20884 26206 20936
rect 26234 20884 26240 20936
rect 26292 20884 26298 20936
rect 26970 20884 26976 20936
rect 27028 20884 27034 20936
rect 27062 20884 27068 20936
rect 27120 20884 27126 20936
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20924 27307 20927
rect 27614 20924 27620 20936
rect 27295 20896 27620 20924
rect 27295 20893 27307 20896
rect 27249 20887 27307 20893
rect 27614 20884 27620 20896
rect 27672 20884 27678 20936
rect 30377 20927 30435 20933
rect 30377 20893 30389 20927
rect 30423 20924 30435 20927
rect 30466 20924 30472 20936
rect 30423 20896 30472 20924
rect 30423 20893 30435 20896
rect 30377 20887 30435 20893
rect 30466 20884 30472 20896
rect 30524 20884 30530 20936
rect 30653 20927 30711 20933
rect 30653 20893 30665 20927
rect 30699 20924 30711 20927
rect 31018 20924 31024 20936
rect 30699 20896 31024 20924
rect 30699 20893 30711 20896
rect 30653 20887 30711 20893
rect 31018 20884 31024 20896
rect 31076 20884 31082 20936
rect 31205 20927 31263 20933
rect 31205 20893 31217 20927
rect 31251 20893 31263 20927
rect 31205 20887 31263 20893
rect 28718 20856 28724 20868
rect 23624 20828 23980 20856
rect 25240 20828 28724 20856
rect 23624 20816 23630 20828
rect 25240 20788 25268 20828
rect 28718 20816 28724 20828
rect 28776 20816 28782 20868
rect 30558 20816 30564 20868
rect 30616 20856 30622 20868
rect 31220 20856 31248 20887
rect 31386 20884 31392 20936
rect 31444 20884 31450 20936
rect 33220 20927 33278 20933
rect 33220 20893 33232 20927
rect 33266 20924 33278 20927
rect 34330 20924 34336 20936
rect 33266 20896 34336 20924
rect 33266 20893 33278 20896
rect 33220 20887 33278 20893
rect 34330 20884 34336 20896
rect 34388 20884 34394 20936
rect 34790 20884 34796 20936
rect 34848 20924 34854 20936
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 34848 20896 34897 20924
rect 34848 20884 34854 20896
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 36630 20884 36636 20936
rect 36688 20884 36694 20936
rect 41230 20933 41236 20936
rect 36900 20927 36958 20933
rect 36900 20893 36912 20927
rect 36946 20924 36958 20927
rect 38933 20927 38991 20933
rect 38933 20924 38945 20927
rect 36946 20896 38945 20924
rect 36946 20893 36958 20896
rect 36900 20887 36958 20893
rect 38933 20893 38945 20896
rect 38979 20893 38991 20927
rect 38933 20887 38991 20893
rect 41224 20887 41236 20933
rect 41230 20884 41236 20887
rect 41288 20884 41294 20936
rect 44652 20933 44680 21032
rect 45112 20992 45140 21100
rect 45186 21088 45192 21140
rect 45244 21088 45250 21140
rect 45112 20964 45692 20992
rect 45664 20933 45692 20964
rect 44453 20927 44511 20933
rect 44453 20893 44465 20927
rect 44499 20893 44511 20927
rect 44453 20887 44511 20893
rect 44637 20927 44695 20933
rect 44637 20893 44649 20927
rect 44683 20924 44695 20927
rect 45465 20927 45523 20933
rect 45465 20924 45477 20927
rect 44683 20896 45477 20924
rect 44683 20893 44695 20896
rect 44637 20887 44695 20893
rect 45465 20893 45477 20896
rect 45511 20893 45523 20927
rect 45465 20887 45523 20893
rect 45557 20927 45615 20933
rect 45557 20893 45569 20927
rect 45603 20893 45615 20927
rect 45557 20887 45615 20893
rect 45649 20927 45707 20933
rect 45649 20893 45661 20927
rect 45695 20893 45707 20927
rect 45649 20887 45707 20893
rect 30616 20828 31248 20856
rect 30616 20816 30622 20828
rect 33594 20816 33600 20868
rect 33652 20856 33658 20868
rect 38565 20859 38623 20865
rect 33652 20828 38148 20856
rect 33652 20816 33658 20828
rect 23124 20760 25268 20788
rect 18656 20748 18662 20760
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25777 20791 25835 20797
rect 25777 20788 25789 20791
rect 25372 20760 25789 20788
rect 25372 20748 25378 20760
rect 25777 20757 25789 20760
rect 25823 20757 25835 20791
rect 25777 20751 25835 20757
rect 26786 20748 26792 20800
rect 26844 20748 26850 20800
rect 34974 20748 34980 20800
rect 35032 20748 35038 20800
rect 38010 20748 38016 20800
rect 38068 20748 38074 20800
rect 38120 20788 38148 20828
rect 38565 20825 38577 20859
rect 38611 20856 38623 20859
rect 38654 20856 38660 20868
rect 38611 20828 38660 20856
rect 38611 20825 38623 20828
rect 38565 20819 38623 20825
rect 38654 20816 38660 20828
rect 38712 20816 38718 20868
rect 38749 20859 38807 20865
rect 38749 20825 38761 20859
rect 38795 20825 38807 20859
rect 44468 20856 44496 20887
rect 45572 20856 45600 20887
rect 45830 20884 45836 20936
rect 45888 20884 45894 20936
rect 45922 20856 45928 20868
rect 44468 20828 45928 20856
rect 38749 20819 38807 20825
rect 38764 20788 38792 20819
rect 45922 20816 45928 20828
rect 45980 20816 45986 20868
rect 38120 20760 38792 20788
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 2130 20544 2136 20596
rect 2188 20584 2194 20596
rect 2958 20584 2964 20596
rect 2188 20556 2964 20584
rect 2188 20544 2194 20556
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3329 20587 3387 20593
rect 3329 20553 3341 20587
rect 3375 20584 3387 20587
rect 3418 20584 3424 20596
rect 3375 20556 3424 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 6638 20544 6644 20596
rect 6696 20544 6702 20596
rect 7009 20587 7067 20593
rect 7009 20553 7021 20587
rect 7055 20584 7067 20587
rect 7742 20584 7748 20596
rect 7055 20556 7748 20584
rect 7055 20553 7067 20556
rect 7009 20547 7067 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 8404 20556 8708 20584
rect 2222 20525 2228 20528
rect 2216 20516 2228 20525
rect 2183 20488 2228 20516
rect 2216 20479 2228 20488
rect 2222 20476 2228 20479
rect 2280 20476 2286 20528
rect 2498 20476 2504 20528
rect 2556 20516 2562 20528
rect 8404 20516 8432 20556
rect 8570 20525 8576 20528
rect 8564 20516 8576 20525
rect 2556 20488 8432 20516
rect 8531 20488 8576 20516
rect 2556 20476 2562 20488
rect 8564 20479 8576 20488
rect 8570 20476 8576 20479
rect 8628 20476 8634 20528
rect 8680 20516 8708 20556
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 11974 20544 11980 20596
rect 12032 20544 12038 20596
rect 12342 20544 12348 20596
rect 12400 20544 12406 20596
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 14369 20587 14427 20593
rect 14369 20584 14381 20587
rect 13504 20556 14381 20584
rect 13504 20544 13510 20556
rect 14369 20553 14381 20556
rect 14415 20553 14427 20587
rect 26694 20584 26700 20596
rect 14369 20547 14427 20553
rect 14936 20556 26700 20584
rect 11422 20516 11428 20528
rect 8680 20488 11428 20516
rect 11422 20476 11428 20488
rect 11480 20476 11486 20528
rect 11992 20516 12020 20544
rect 12069 20519 12127 20525
rect 12069 20516 12081 20519
rect 11992 20488 12081 20516
rect 12069 20485 12081 20488
rect 12115 20485 12127 20519
rect 14826 20516 14832 20528
rect 12069 20479 12127 20485
rect 13188 20488 14832 20516
rect 1670 20408 1676 20460
rect 1728 20448 1734 20460
rect 1949 20451 2007 20457
rect 1949 20448 1961 20451
rect 1728 20420 1961 20448
rect 1728 20408 1734 20420
rect 1949 20417 1961 20420
rect 1995 20417 2007 20451
rect 3881 20451 3939 20457
rect 3881 20448 3893 20451
rect 1949 20411 2007 20417
rect 2056 20420 3893 20448
rect 934 20340 940 20392
rect 992 20380 998 20392
rect 2056 20380 2084 20420
rect 3881 20417 3893 20420
rect 3927 20417 3939 20451
rect 6822 20448 6828 20460
rect 3881 20411 3939 20417
rect 3988 20420 6828 20448
rect 992 20352 2084 20380
rect 992 20340 998 20352
rect 2958 20340 2964 20392
rect 3016 20380 3022 20392
rect 3988 20380 4016 20420
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 8128 20420 9352 20448
rect 3016 20352 4016 20380
rect 3016 20340 3022 20352
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 7101 20383 7159 20389
rect 7101 20380 7113 20383
rect 4764 20352 7113 20380
rect 4764 20340 4770 20352
rect 7101 20349 7113 20352
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 7282 20340 7288 20392
rect 7340 20340 7346 20392
rect 8128 20312 8156 20420
rect 8202 20340 8208 20392
rect 8260 20380 8266 20392
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 8260 20352 8309 20380
rect 8260 20340 8266 20352
rect 8297 20349 8309 20352
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 2884 20284 8156 20312
rect 9324 20312 9352 20420
rect 10410 20408 10416 20460
rect 10468 20448 10474 20460
rect 11606 20448 11612 20460
rect 10468 20420 11612 20448
rect 10468 20408 10474 20420
rect 11606 20408 11612 20420
rect 11664 20448 11670 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 11664 20420 11713 20448
rect 11664 20408 11670 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11790 20408 11796 20460
rect 11848 20408 11854 20460
rect 12250 20457 12256 20460
rect 11977 20451 12035 20457
rect 11977 20417 11989 20451
rect 12023 20448 12035 20451
rect 12207 20451 12256 20457
rect 12023 20420 12112 20448
rect 12023 20417 12035 20420
rect 11977 20411 12035 20417
rect 12084 20380 12112 20420
rect 12207 20417 12219 20451
rect 12253 20417 12256 20451
rect 12207 20411 12256 20417
rect 12250 20408 12256 20411
rect 12308 20408 12314 20460
rect 12986 20408 12992 20460
rect 13044 20448 13050 20460
rect 13188 20448 13216 20488
rect 14826 20476 14832 20488
rect 14884 20476 14890 20528
rect 13044 20420 13216 20448
rect 13256 20451 13314 20457
rect 13044 20408 13050 20420
rect 13256 20417 13268 20451
rect 13302 20448 13314 20451
rect 13722 20448 13728 20460
rect 13302 20420 13728 20448
rect 13302 20417 13314 20420
rect 13256 20411 13314 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 14936 20448 14964 20556
rect 26694 20544 26700 20556
rect 26752 20544 26758 20596
rect 27154 20544 27160 20596
rect 27212 20544 27218 20596
rect 28902 20544 28908 20596
rect 28960 20584 28966 20596
rect 30101 20587 30159 20593
rect 30101 20584 30113 20587
rect 28960 20556 30113 20584
rect 28960 20544 28966 20556
rect 30101 20553 30113 20556
rect 30147 20553 30159 20587
rect 30101 20547 30159 20553
rect 33689 20587 33747 20593
rect 33689 20553 33701 20587
rect 33735 20584 33747 20587
rect 33870 20584 33876 20596
rect 33735 20556 33876 20584
rect 33735 20553 33747 20556
rect 33689 20547 33747 20553
rect 33870 20544 33876 20556
rect 33928 20544 33934 20596
rect 37642 20544 37648 20596
rect 37700 20584 37706 20596
rect 38010 20584 38016 20596
rect 37700 20556 38016 20584
rect 37700 20544 37706 20556
rect 38010 20544 38016 20556
rect 38068 20584 38074 20596
rect 44450 20584 44456 20596
rect 38068 20556 44456 20584
rect 38068 20544 38074 20556
rect 44450 20544 44456 20556
rect 44508 20544 44514 20596
rect 15188 20519 15246 20525
rect 15188 20485 15200 20519
rect 15234 20516 15246 20519
rect 17770 20516 17776 20528
rect 15234 20488 17776 20516
rect 15234 20485 15246 20488
rect 15188 20479 15246 20485
rect 17770 20476 17776 20488
rect 17828 20476 17834 20528
rect 20162 20516 20168 20528
rect 18248 20488 20168 20516
rect 18248 20457 18276 20488
rect 20162 20476 20168 20488
rect 20220 20476 20226 20528
rect 34149 20519 34207 20525
rect 25884 20488 29776 20516
rect 14844 20420 14964 20448
rect 18233 20451 18291 20457
rect 12342 20380 12348 20392
rect 12084 20352 12348 20380
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 9324 20284 13032 20312
rect 2314 20204 2320 20256
rect 2372 20244 2378 20256
rect 2884 20244 2912 20284
rect 2372 20216 2912 20244
rect 2372 20204 2378 20216
rect 3970 20204 3976 20256
rect 4028 20204 4034 20256
rect 6178 20204 6184 20256
rect 6236 20244 6242 20256
rect 6638 20244 6644 20256
rect 6236 20216 6644 20244
rect 6236 20204 6242 20216
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 6822 20204 6828 20256
rect 6880 20244 6886 20256
rect 8662 20244 8668 20256
rect 6880 20216 8668 20244
rect 6880 20204 6886 20216
rect 8662 20204 8668 20216
rect 8720 20204 8726 20256
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 11698 20244 11704 20256
rect 10560 20216 11704 20244
rect 10560 20204 10566 20216
rect 11698 20204 11704 20216
rect 11756 20244 11762 20256
rect 12894 20244 12900 20256
rect 11756 20216 12900 20244
rect 11756 20204 11762 20216
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 13004 20244 13032 20284
rect 14844 20244 14872 20420
rect 18233 20417 18245 20451
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 19334 20457 19340 20460
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 18840 20420 19073 20448
rect 18840 20408 18846 20420
rect 19061 20417 19073 20420
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 19328 20411 19340 20457
rect 19334 20408 19340 20411
rect 19392 20408 19398 20460
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20349 14979 20383
rect 14921 20343 14979 20349
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20380 18383 20383
rect 18506 20380 18512 20392
rect 18371 20352 18512 20380
rect 18371 20349 18383 20352
rect 18325 20343 18383 20349
rect 13004 20216 14872 20244
rect 14936 20244 14964 20343
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 25777 20383 25835 20389
rect 25777 20380 25789 20383
rect 20772 20352 25789 20380
rect 20772 20340 20778 20352
rect 25777 20349 25789 20352
rect 25823 20349 25835 20383
rect 25884 20380 25912 20488
rect 25961 20451 26019 20457
rect 25961 20417 25973 20451
rect 26007 20448 26019 20451
rect 26786 20448 26792 20460
rect 26007 20420 26792 20448
rect 26007 20417 26019 20420
rect 25961 20411 26019 20417
rect 26786 20408 26792 20420
rect 26844 20408 26850 20460
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27120 20420 27476 20448
rect 27120 20408 27126 20420
rect 27448 20392 27476 20420
rect 28810 20408 28816 20460
rect 28868 20448 28874 20460
rect 28977 20451 29035 20457
rect 28977 20448 28989 20451
rect 28868 20420 28989 20448
rect 28868 20408 28874 20420
rect 28977 20417 28989 20420
rect 29023 20417 29035 20451
rect 28977 20411 29035 20417
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 25884 20352 26065 20380
rect 25777 20343 25835 20349
rect 26053 20349 26065 20352
rect 26099 20349 26111 20383
rect 26053 20343 26111 20349
rect 26142 20340 26148 20392
rect 26200 20340 26206 20392
rect 26234 20340 26240 20392
rect 26292 20380 26298 20392
rect 26878 20380 26884 20392
rect 26292 20352 26884 20380
rect 26292 20340 26298 20352
rect 26878 20340 26884 20352
rect 26936 20340 26942 20392
rect 27154 20340 27160 20392
rect 27212 20380 27218 20392
rect 27338 20380 27344 20392
rect 27212 20352 27344 20380
rect 27212 20340 27218 20352
rect 27338 20340 27344 20352
rect 27396 20340 27402 20392
rect 27430 20340 27436 20392
rect 27488 20340 27494 20392
rect 27522 20340 27528 20392
rect 27580 20340 27586 20392
rect 27614 20340 27620 20392
rect 27672 20340 27678 20392
rect 28721 20383 28779 20389
rect 28721 20349 28733 20383
rect 28767 20349 28779 20383
rect 28721 20343 28779 20349
rect 16301 20315 16359 20321
rect 16301 20281 16313 20315
rect 16347 20312 16359 20315
rect 17678 20312 17684 20324
rect 16347 20284 17684 20312
rect 16347 20281 16359 20284
rect 16301 20275 16359 20281
rect 17678 20272 17684 20284
rect 17736 20272 17742 20324
rect 20162 20272 20168 20324
rect 20220 20312 20226 20324
rect 20441 20315 20499 20321
rect 20441 20312 20453 20315
rect 20220 20284 20453 20312
rect 20220 20272 20226 20284
rect 20441 20281 20453 20284
rect 20487 20281 20499 20315
rect 26160 20312 26188 20340
rect 26326 20312 26332 20324
rect 26160 20284 26332 20312
rect 20441 20275 20499 20281
rect 26326 20272 26332 20284
rect 26384 20272 26390 20324
rect 15286 20244 15292 20256
rect 14936 20216 15292 20244
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 18601 20247 18659 20253
rect 18601 20213 18613 20247
rect 18647 20244 18659 20247
rect 19426 20244 19432 20256
rect 18647 20216 19432 20244
rect 18647 20213 18659 20216
rect 18601 20207 18659 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 28736 20244 28764 20343
rect 29748 20312 29776 20488
rect 34149 20485 34161 20519
rect 34195 20516 34207 20519
rect 34514 20516 34520 20528
rect 34195 20488 34520 20516
rect 34195 20485 34207 20488
rect 34149 20479 34207 20485
rect 34514 20476 34520 20488
rect 34572 20516 34578 20528
rect 40218 20516 40224 20528
rect 34572 20488 35020 20516
rect 34572 20476 34578 20488
rect 34992 20460 35020 20488
rect 37476 20488 40224 20516
rect 30006 20408 30012 20460
rect 30064 20448 30070 20460
rect 30561 20451 30619 20457
rect 30561 20448 30573 20451
rect 30064 20420 30573 20448
rect 30064 20408 30070 20420
rect 30561 20417 30573 20420
rect 30607 20417 30619 20451
rect 30561 20411 30619 20417
rect 34057 20451 34115 20457
rect 34057 20417 34069 20451
rect 34103 20448 34115 20451
rect 34698 20448 34704 20460
rect 34103 20420 34704 20448
rect 34103 20417 34115 20420
rect 34057 20411 34115 20417
rect 34698 20408 34704 20420
rect 34756 20408 34762 20460
rect 34790 20408 34796 20460
rect 34848 20448 34854 20460
rect 34885 20451 34943 20457
rect 34885 20448 34897 20451
rect 34848 20420 34897 20448
rect 34848 20408 34854 20420
rect 34885 20417 34897 20420
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 34974 20408 34980 20460
rect 35032 20448 35038 20460
rect 35069 20451 35127 20457
rect 35069 20448 35081 20451
rect 35032 20420 35081 20448
rect 35032 20408 35038 20420
rect 35069 20417 35081 20420
rect 35115 20417 35127 20451
rect 35069 20411 35127 20417
rect 36538 20408 36544 20460
rect 36596 20448 36602 20460
rect 37090 20448 37096 20460
rect 36596 20420 37096 20448
rect 36596 20408 36602 20420
rect 37090 20408 37096 20420
rect 37148 20448 37154 20460
rect 37476 20457 37504 20488
rect 40218 20476 40224 20488
rect 40276 20476 40282 20528
rect 37734 20457 37740 20460
rect 37461 20451 37519 20457
rect 37461 20448 37473 20451
rect 37148 20420 37473 20448
rect 37148 20408 37154 20420
rect 37461 20417 37473 20420
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 37728 20411 37740 20457
rect 37734 20408 37740 20411
rect 37792 20408 37798 20460
rect 40236 20448 40264 20476
rect 40681 20451 40739 20457
rect 40681 20448 40693 20451
rect 40236 20420 40693 20448
rect 40681 20417 40693 20420
rect 40727 20417 40739 20451
rect 40681 20411 40739 20417
rect 40948 20451 41006 20457
rect 40948 20417 40960 20451
rect 40994 20448 41006 20451
rect 41414 20448 41420 20460
rect 40994 20420 41420 20448
rect 40994 20417 41006 20420
rect 40948 20411 41006 20417
rect 41414 20408 41420 20420
rect 41472 20408 41478 20460
rect 29914 20340 29920 20392
rect 29972 20380 29978 20392
rect 30190 20380 30196 20392
rect 29972 20352 30196 20380
rect 29972 20340 29978 20352
rect 30190 20340 30196 20352
rect 30248 20380 30254 20392
rect 30837 20383 30895 20389
rect 30837 20380 30849 20383
rect 30248 20352 30849 20380
rect 30248 20340 30254 20352
rect 30837 20349 30849 20352
rect 30883 20380 30895 20383
rect 32030 20380 32036 20392
rect 30883 20352 32036 20380
rect 30883 20349 30895 20352
rect 30837 20343 30895 20349
rect 32030 20340 32036 20352
rect 32088 20340 32094 20392
rect 33778 20340 33784 20392
rect 33836 20380 33842 20392
rect 34241 20383 34299 20389
rect 34241 20380 34253 20383
rect 33836 20352 34253 20380
rect 33836 20340 33842 20352
rect 34241 20349 34253 20352
rect 34287 20349 34299 20383
rect 34241 20343 34299 20349
rect 29748 20284 37504 20312
rect 29822 20244 29828 20256
rect 28736 20216 29828 20244
rect 29822 20204 29828 20216
rect 29880 20204 29886 20256
rect 30006 20204 30012 20256
rect 30064 20244 30070 20256
rect 34422 20244 34428 20256
rect 30064 20216 34428 20244
rect 30064 20204 30070 20216
rect 34422 20204 34428 20216
rect 34480 20204 34486 20256
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 34977 20247 35035 20253
rect 34977 20244 34989 20247
rect 34756 20216 34989 20244
rect 34756 20204 34762 20216
rect 34977 20213 34989 20216
rect 35023 20213 35035 20247
rect 37476 20244 37504 20284
rect 38102 20244 38108 20256
rect 37476 20216 38108 20244
rect 34977 20207 35035 20213
rect 38102 20204 38108 20216
rect 38160 20204 38166 20256
rect 38838 20204 38844 20256
rect 38896 20204 38902 20256
rect 42058 20204 42064 20256
rect 42116 20204 42122 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 6546 20000 6552 20052
rect 6604 20040 6610 20052
rect 10410 20040 10416 20052
rect 6604 20012 10416 20040
rect 6604 20000 6610 20012
rect 10410 20000 10416 20012
rect 10468 20000 10474 20052
rect 10502 20000 10508 20052
rect 10560 20000 10566 20052
rect 11790 20040 11796 20052
rect 11164 20012 11796 20040
rect 5445 19975 5503 19981
rect 5445 19941 5457 19975
rect 5491 19972 5503 19975
rect 7466 19972 7472 19984
rect 5491 19944 7472 19972
rect 5491 19941 5503 19944
rect 5445 19935 5503 19941
rect 7466 19932 7472 19944
rect 7524 19932 7530 19984
rect 934 19864 940 19916
rect 992 19904 998 19916
rect 2777 19907 2835 19913
rect 2777 19904 2789 19907
rect 992 19876 2789 19904
rect 992 19864 998 19876
rect 2777 19873 2789 19876
rect 2823 19873 2835 19907
rect 5316 19907 5374 19913
rect 5316 19904 5328 19907
rect 2777 19867 2835 19873
rect 5092 19876 5328 19904
rect 1026 19796 1032 19848
rect 1084 19836 1090 19848
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1084 19808 1685 19836
rect 1084 19796 1090 19808
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 2498 19796 2504 19848
rect 2556 19796 2562 19848
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 4065 19771 4123 19777
rect 4065 19768 4077 19771
rect 992 19740 4077 19768
rect 992 19728 998 19740
rect 4065 19737 4077 19740
rect 4111 19737 4123 19771
rect 4065 19731 4123 19737
rect 4433 19771 4491 19777
rect 4433 19737 4445 19771
rect 4479 19768 4491 19771
rect 4614 19768 4620 19780
rect 4479 19740 4620 19768
rect 4479 19737 4491 19740
rect 4433 19731 4491 19737
rect 4614 19728 4620 19740
rect 4672 19728 4678 19780
rect 5092 19768 5120 19876
rect 5316 19873 5328 19876
rect 5362 19873 5374 19907
rect 5316 19867 5374 19873
rect 5534 19864 5540 19916
rect 5592 19864 5598 19916
rect 6454 19864 6460 19916
rect 6512 19864 6518 19916
rect 8662 19864 8668 19916
rect 8720 19904 8726 19916
rect 8720 19876 10732 19904
rect 8720 19864 8726 19876
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19836 5227 19839
rect 5442 19836 5448 19848
rect 5215 19808 5448 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 5994 19796 6000 19848
rect 6052 19836 6058 19848
rect 6365 19839 6423 19845
rect 6365 19836 6377 19839
rect 6052 19808 6377 19836
rect 6052 19796 6058 19808
rect 6365 19805 6377 19808
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 6730 19836 6736 19848
rect 6687 19808 6736 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 6656 19768 6684 19799
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 8202 19796 8208 19848
rect 8260 19836 8266 19848
rect 10704 19845 10732 19876
rect 9861 19839 9919 19845
rect 9861 19836 9873 19839
rect 8260 19808 9873 19836
rect 8260 19796 8266 19808
rect 9861 19805 9873 19808
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19836 10839 19839
rect 11164 19836 11192 20012
rect 11790 20000 11796 20012
rect 11848 20040 11854 20052
rect 12802 20040 12808 20052
rect 11848 20012 12808 20040
rect 11848 20000 11854 20012
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 13630 20040 13636 20052
rect 12952 20012 13636 20040
rect 12952 20000 12958 20012
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 13722 20000 13728 20052
rect 13780 20000 13786 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16172 20012 16865 20040
rect 16172 20000 16178 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19429 20043 19487 20049
rect 19429 20040 19441 20043
rect 19392 20012 19441 20040
rect 19392 20000 19398 20012
rect 19429 20009 19441 20012
rect 19475 20009 19487 20043
rect 19429 20003 19487 20009
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 24581 20043 24639 20049
rect 24581 20040 24593 20043
rect 23716 20012 24593 20040
rect 23716 20000 23722 20012
rect 24581 20009 24593 20012
rect 24627 20009 24639 20043
rect 24581 20003 24639 20009
rect 24946 20000 24952 20052
rect 25004 20040 25010 20052
rect 25961 20043 26019 20049
rect 25961 20040 25973 20043
rect 25004 20012 25973 20040
rect 25004 20000 25010 20012
rect 25961 20009 25973 20012
rect 26007 20009 26019 20043
rect 25961 20003 26019 20009
rect 28721 20043 28779 20049
rect 28721 20009 28733 20043
rect 28767 20040 28779 20043
rect 28810 20040 28816 20052
rect 28767 20012 28816 20040
rect 28767 20009 28779 20012
rect 28721 20003 28779 20009
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 37734 20000 37740 20052
rect 37792 20000 37798 20052
rect 41414 20000 41420 20052
rect 41472 20000 41478 20052
rect 25130 19972 25136 19984
rect 11256 19944 18184 19972
rect 11256 19913 11284 19944
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19873 11299 19907
rect 11241 19867 11299 19873
rect 11422 19864 11428 19916
rect 11480 19904 11486 19916
rect 11882 19904 11888 19916
rect 11480 19876 11888 19904
rect 11480 19864 11486 19876
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13262 19864 13268 19916
rect 13320 19904 13326 19916
rect 13320 19876 13584 19904
rect 13320 19864 13326 19876
rect 10827 19808 11192 19836
rect 10827 19805 10839 19808
rect 10781 19799 10839 19805
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 13081 19839 13139 19845
rect 13081 19836 13093 19839
rect 11664 19808 13093 19836
rect 11664 19796 11670 19808
rect 13081 19805 13093 19808
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 13170 19796 13176 19848
rect 13228 19796 13234 19848
rect 13446 19796 13452 19848
rect 13504 19796 13510 19848
rect 13556 19845 13584 19876
rect 13630 19864 13636 19916
rect 13688 19904 13694 19916
rect 16945 19907 17003 19913
rect 13688 19876 16712 19904
rect 13688 19864 13694 19876
rect 13546 19839 13604 19845
rect 13546 19805 13558 19839
rect 13592 19805 13604 19839
rect 13546 19799 13604 19805
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 16684 19845 16712 19876
rect 16945 19873 16957 19907
rect 16991 19904 17003 19907
rect 18046 19904 18052 19916
rect 16991 19876 18052 19904
rect 16991 19873 17003 19876
rect 16945 19867 17003 19873
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 18156 19904 18184 19944
rect 19260 19944 25136 19972
rect 19260 19904 19288 19944
rect 18156 19876 19288 19904
rect 19352 19876 21220 19904
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 14884 19808 15853 19836
rect 14884 19796 14890 19808
rect 15841 19805 15853 19808
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19836 16727 19839
rect 19242 19836 19248 19848
rect 16715 19808 19248 19836
rect 16715 19805 16727 19808
rect 16669 19799 16727 19805
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 5092 19740 6684 19768
rect 7101 19771 7159 19777
rect 7101 19737 7113 19771
rect 7147 19768 7159 19771
rect 7834 19768 7840 19780
rect 7147 19740 7840 19768
rect 7147 19737 7159 19740
rect 7101 19731 7159 19737
rect 7834 19728 7840 19740
rect 7892 19728 7898 19780
rect 9122 19728 9128 19780
rect 9180 19728 9186 19780
rect 11146 19728 11152 19780
rect 11204 19768 11210 19780
rect 11624 19768 11652 19796
rect 11204 19740 11652 19768
rect 11204 19728 11210 19740
rect 13354 19728 13360 19780
rect 13412 19728 13418 19780
rect 15102 19768 15108 19780
rect 13648 19740 15108 19768
rect 1946 19660 1952 19712
rect 2004 19660 2010 19712
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 5813 19703 5871 19709
rect 5813 19700 5825 19703
rect 5500 19672 5825 19700
rect 5500 19660 5506 19672
rect 5813 19669 5825 19672
rect 5859 19669 5871 19703
rect 5813 19663 5871 19669
rect 6270 19660 6276 19712
rect 6328 19700 6334 19712
rect 7190 19700 7196 19712
rect 6328 19672 7196 19700
rect 6328 19660 6334 19672
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 9140 19700 9168 19728
rect 13648 19700 13676 19740
rect 15102 19728 15108 19740
rect 15160 19728 15166 19780
rect 16114 19728 16120 19780
rect 16172 19768 16178 19780
rect 19352 19768 19380 19876
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 20254 19836 20260 19848
rect 19659 19808 20260 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 19628 19768 19656 19799
rect 20254 19796 20260 19808
rect 20312 19796 20318 19848
rect 20806 19796 20812 19848
rect 20864 19796 20870 19848
rect 21192 19830 21220 19876
rect 21358 19830 21364 19848
rect 21192 19802 21364 19830
rect 21358 19796 21364 19802
rect 21416 19796 21422 19848
rect 23492 19836 23520 19944
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 27522 19932 27528 19984
rect 27580 19972 27586 19984
rect 27580 19944 37044 19972
rect 27580 19932 27586 19944
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 26421 19907 26479 19913
rect 26421 19904 26433 19907
rect 23624 19876 26433 19904
rect 23624 19864 23630 19876
rect 26421 19873 26433 19876
rect 26467 19873 26479 19907
rect 26421 19867 26479 19873
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 29362 19904 29368 19916
rect 26752 19876 29368 19904
rect 26752 19864 26758 19876
rect 29362 19864 29368 19876
rect 29420 19864 29426 19916
rect 30926 19864 30932 19916
rect 30984 19864 30990 19916
rect 33502 19864 33508 19916
rect 33560 19904 33566 19916
rect 33560 19876 34652 19904
rect 33560 19864 33566 19876
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23492 19808 23673 19836
rect 23661 19805 23673 19808
rect 23707 19805 23719 19839
rect 23937 19839 23995 19845
rect 23937 19836 23949 19839
rect 23661 19799 23719 19805
rect 23768 19808 23949 19836
rect 16172 19740 19380 19768
rect 19444 19740 19656 19768
rect 16172 19728 16178 19740
rect 19444 19712 19472 19740
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 23768 19768 23796 19808
rect 23937 19805 23949 19808
rect 23983 19805 23995 19839
rect 23937 19799 23995 19805
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 24854 19796 24860 19848
rect 24912 19796 24918 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 22336 19740 23796 19768
rect 23845 19771 23903 19777
rect 22336 19728 22342 19740
rect 23845 19737 23857 19771
rect 23891 19768 23903 19771
rect 24394 19768 24400 19780
rect 23891 19740 24400 19768
rect 23891 19737 23903 19740
rect 23845 19731 23903 19737
rect 24394 19728 24400 19740
rect 24452 19768 24458 19780
rect 24964 19768 24992 19799
rect 25038 19796 25044 19848
rect 25096 19796 25102 19848
rect 26050 19796 26056 19848
rect 26108 19836 26114 19848
rect 26145 19839 26203 19845
rect 26145 19836 26157 19839
rect 26108 19808 26157 19836
rect 26108 19796 26114 19808
rect 26145 19805 26157 19808
rect 26191 19805 26203 19839
rect 26145 19799 26203 19805
rect 26234 19796 26240 19848
rect 26292 19796 26298 19848
rect 26326 19796 26332 19848
rect 26384 19796 26390 19848
rect 28718 19796 28724 19848
rect 28776 19836 28782 19848
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28776 19808 28917 19836
rect 28776 19796 28782 19808
rect 28905 19805 28917 19808
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 29181 19839 29239 19845
rect 29181 19805 29193 19839
rect 29227 19836 29239 19839
rect 29914 19836 29920 19848
rect 29227 19808 29920 19836
rect 29227 19805 29239 19808
rect 29181 19799 29239 19805
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 34149 19839 34207 19845
rect 34149 19805 34161 19839
rect 34195 19836 34207 19839
rect 34514 19836 34520 19848
rect 34195 19808 34520 19836
rect 34195 19805 34207 19808
rect 34149 19799 34207 19805
rect 34514 19796 34520 19808
rect 34572 19796 34578 19848
rect 34624 19836 34652 19876
rect 37016 19836 37044 19944
rect 37458 19932 37464 19984
rect 37516 19972 37522 19984
rect 38838 19972 38844 19984
rect 37516 19944 38844 19972
rect 37516 19932 37522 19944
rect 37090 19864 37096 19916
rect 37148 19864 37154 19916
rect 38304 19913 38332 19944
rect 38838 19932 38844 19944
rect 38896 19932 38902 19984
rect 38289 19907 38347 19913
rect 38289 19873 38301 19907
rect 38335 19904 38347 19907
rect 38335 19876 38369 19904
rect 38335 19873 38347 19876
rect 38289 19867 38347 19873
rect 38654 19864 38660 19916
rect 38712 19904 38718 19916
rect 45189 19907 45247 19913
rect 45189 19904 45201 19907
rect 38712 19876 45201 19904
rect 38712 19864 38718 19876
rect 45189 19873 45201 19876
rect 45235 19873 45247 19907
rect 45189 19867 45247 19873
rect 37458 19836 37464 19848
rect 34624 19808 36952 19836
rect 37016 19808 37464 19836
rect 30006 19768 30012 19780
rect 24452 19740 24992 19768
rect 28736 19740 30012 19768
rect 24452 19728 24458 19740
rect 9140 19672 13676 19700
rect 16482 19660 16488 19712
rect 16540 19660 16546 19712
rect 19426 19660 19432 19712
rect 19484 19660 19490 19712
rect 20898 19660 20904 19712
rect 20956 19660 20962 19712
rect 23474 19660 23480 19712
rect 23532 19660 23538 19712
rect 24302 19660 24308 19712
rect 24360 19700 24366 19712
rect 28736 19700 28764 19740
rect 30006 19728 30012 19740
rect 30064 19728 30070 19780
rect 30098 19728 30104 19780
rect 30156 19768 30162 19780
rect 30193 19771 30251 19777
rect 30193 19768 30205 19771
rect 30156 19740 30205 19768
rect 30156 19728 30162 19740
rect 30193 19737 30205 19740
rect 30239 19737 30251 19771
rect 30193 19731 30251 19737
rect 33965 19771 34023 19777
rect 33965 19737 33977 19771
rect 34011 19768 34023 19771
rect 34790 19768 34796 19780
rect 34011 19740 34796 19768
rect 34011 19737 34023 19740
rect 33965 19731 34023 19737
rect 34790 19728 34796 19740
rect 34848 19728 34854 19780
rect 36354 19728 36360 19780
rect 36412 19728 36418 19780
rect 36924 19768 36952 19808
rect 37458 19796 37464 19808
rect 37516 19796 37522 19848
rect 37921 19839 37979 19845
rect 37921 19805 37933 19839
rect 37967 19805 37979 19839
rect 37921 19799 37979 19805
rect 37936 19768 37964 19799
rect 38010 19796 38016 19848
rect 38068 19796 38074 19848
rect 38381 19839 38439 19845
rect 38381 19836 38393 19839
rect 38212 19808 38393 19836
rect 36924 19740 37964 19768
rect 24360 19672 28764 19700
rect 24360 19660 24366 19672
rect 28902 19660 28908 19712
rect 28960 19700 28966 19712
rect 29089 19703 29147 19709
rect 29089 19700 29101 19703
rect 28960 19672 29101 19700
rect 28960 19660 28966 19672
rect 29089 19669 29101 19672
rect 29135 19669 29147 19703
rect 29089 19663 29147 19669
rect 29178 19660 29184 19712
rect 29236 19700 29242 19712
rect 30282 19700 30288 19712
rect 29236 19672 30288 19700
rect 29236 19660 29242 19672
rect 30282 19660 30288 19672
rect 30340 19660 30346 19712
rect 34330 19660 34336 19712
rect 34388 19660 34394 19712
rect 34882 19660 34888 19712
rect 34940 19700 34946 19712
rect 38212 19700 38240 19808
rect 38381 19805 38393 19808
rect 38427 19836 38439 19839
rect 40402 19836 40408 19848
rect 38427 19808 40408 19836
rect 38427 19805 38439 19808
rect 38381 19799 38439 19805
rect 40402 19796 40408 19808
rect 40460 19796 40466 19848
rect 41417 19839 41475 19845
rect 41417 19805 41429 19839
rect 41463 19805 41475 19839
rect 41417 19799 41475 19805
rect 41432 19768 41460 19799
rect 41598 19796 41604 19848
rect 41656 19796 41662 19848
rect 42058 19796 42064 19848
rect 42116 19836 42122 19848
rect 44174 19836 44180 19848
rect 42116 19808 44180 19836
rect 42116 19796 42122 19808
rect 44174 19796 44180 19808
rect 44232 19796 44238 19848
rect 44450 19796 44456 19848
rect 44508 19836 44514 19848
rect 45465 19839 45523 19845
rect 45465 19836 45477 19839
rect 44508 19808 45477 19836
rect 44508 19796 44514 19808
rect 45465 19805 45477 19808
rect 45511 19805 45523 19839
rect 45465 19799 45523 19805
rect 45554 19796 45560 19848
rect 45612 19796 45618 19848
rect 45646 19796 45652 19848
rect 45704 19796 45710 19848
rect 45830 19796 45836 19848
rect 45888 19796 45894 19848
rect 42886 19768 42892 19780
rect 41432 19740 42892 19768
rect 42886 19728 42892 19740
rect 42944 19728 42950 19780
rect 34940 19672 38240 19700
rect 34940 19660 34946 19672
rect 38562 19660 38568 19712
rect 38620 19700 38626 19712
rect 43346 19700 43352 19712
rect 38620 19672 43352 19700
rect 38620 19660 38626 19672
rect 43346 19660 43352 19672
rect 43404 19660 43410 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 2685 19499 2743 19505
rect 2685 19465 2697 19499
rect 2731 19496 2743 19499
rect 3970 19496 3976 19508
rect 2731 19468 3976 19496
rect 2731 19465 2743 19468
rect 2685 19459 2743 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 5994 19456 6000 19508
rect 6052 19456 6058 19508
rect 6362 19456 6368 19508
rect 6420 19496 6426 19508
rect 7193 19499 7251 19505
rect 7193 19496 7205 19499
rect 6420 19468 7205 19496
rect 6420 19456 6426 19468
rect 7193 19465 7205 19468
rect 7239 19465 7251 19499
rect 7193 19459 7251 19465
rect 9858 19456 9864 19508
rect 9916 19456 9922 19508
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 16114 19496 16120 19508
rect 12860 19468 16120 19496
rect 12860 19456 12866 19468
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 16758 19496 16764 19508
rect 16255 19468 16764 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 20898 19456 20904 19508
rect 20956 19496 20962 19508
rect 24302 19496 24308 19508
rect 20956 19468 24308 19496
rect 20956 19456 20962 19468
rect 24302 19456 24308 19468
rect 24360 19456 24366 19508
rect 24394 19456 24400 19508
rect 24452 19456 24458 19508
rect 26050 19456 26056 19508
rect 26108 19456 26114 19508
rect 29365 19499 29423 19505
rect 29365 19465 29377 19499
rect 29411 19496 29423 19499
rect 32490 19496 32496 19508
rect 29411 19468 32496 19496
rect 29411 19465 29423 19468
rect 29365 19459 29423 19465
rect 32490 19456 32496 19468
rect 32548 19456 32554 19508
rect 32582 19456 32588 19508
rect 32640 19456 32646 19508
rect 44913 19499 44971 19505
rect 32692 19468 43116 19496
rect 2593 19431 2651 19437
rect 2593 19397 2605 19431
rect 2639 19428 2651 19431
rect 3234 19428 3240 19440
rect 2639 19400 3240 19428
rect 2639 19397 2651 19400
rect 2593 19391 2651 19397
rect 3234 19388 3240 19400
rect 3292 19428 3298 19440
rect 5534 19428 5540 19440
rect 3292 19400 5540 19428
rect 3292 19388 3298 19400
rect 5534 19388 5540 19400
rect 5592 19388 5598 19440
rect 6178 19388 6184 19440
rect 6236 19428 6242 19440
rect 6236 19400 6684 19428
rect 6236 19388 6242 19400
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19329 3571 19363
rect 3513 19323 3571 19329
rect 5629 19363 5687 19369
rect 5629 19329 5641 19363
rect 5675 19360 5687 19363
rect 6270 19360 6276 19372
rect 5675 19332 6276 19360
rect 5675 19329 5687 19332
rect 5629 19323 5687 19329
rect 2682 19252 2688 19304
rect 2740 19292 2746 19304
rect 2777 19295 2835 19301
rect 2777 19292 2789 19295
rect 2740 19264 2789 19292
rect 2740 19252 2746 19264
rect 2777 19261 2789 19264
rect 2823 19261 2835 19295
rect 2777 19255 2835 19261
rect 934 19184 940 19236
rect 992 19224 998 19236
rect 3528 19224 3556 19323
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 6656 19369 6684 19400
rect 6730 19388 6736 19440
rect 6788 19428 6794 19440
rect 6917 19431 6975 19437
rect 6917 19428 6929 19431
rect 6788 19400 6929 19428
rect 6788 19388 6794 19400
rect 6917 19397 6929 19400
rect 6963 19397 6975 19431
rect 9582 19428 9588 19440
rect 6917 19391 6975 19397
rect 8128 19400 9588 19428
rect 6642 19363 6700 19369
rect 6642 19329 6654 19363
rect 6688 19329 6700 19363
rect 6642 19323 6700 19329
rect 6822 19320 6828 19372
rect 6880 19320 6886 19372
rect 7055 19363 7113 19369
rect 7055 19329 7067 19363
rect 7101 19360 7113 19363
rect 8128 19360 8156 19400
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 15096 19431 15154 19437
rect 15096 19397 15108 19431
rect 15142 19428 15154 19431
rect 16482 19428 16488 19440
rect 15142 19400 16488 19428
rect 15142 19397 15154 19400
rect 15096 19391 15154 19397
rect 16482 19388 16488 19400
rect 16540 19388 16546 19440
rect 20990 19388 20996 19440
rect 21048 19428 21054 19440
rect 23284 19431 23342 19437
rect 21048 19400 23244 19428
rect 21048 19388 21054 19400
rect 7101 19332 8156 19360
rect 7101 19329 7113 19332
rect 7055 19323 7113 19329
rect 8202 19320 8208 19372
rect 8260 19360 8266 19372
rect 8481 19363 8539 19369
rect 8481 19360 8493 19363
rect 8260 19332 8493 19360
rect 8260 19320 8266 19332
rect 8481 19329 8493 19332
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 8748 19363 8806 19369
rect 8748 19329 8760 19363
rect 8794 19360 8806 19363
rect 10134 19360 10140 19372
rect 8794 19332 10140 19360
rect 8794 19329 8806 19332
rect 8748 19323 8806 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 14826 19320 14832 19372
rect 14884 19320 14890 19372
rect 23017 19363 23075 19369
rect 23017 19329 23029 19363
rect 23063 19329 23075 19363
rect 23216 19360 23244 19400
rect 23284 19397 23296 19431
rect 23330 19428 23342 19431
rect 23474 19428 23480 19440
rect 23330 19400 23480 19428
rect 23330 19397 23342 19400
rect 23284 19391 23342 19397
rect 23474 19388 23480 19400
rect 23532 19388 23538 19440
rect 25958 19388 25964 19440
rect 26016 19428 26022 19440
rect 27430 19428 27436 19440
rect 26016 19400 27436 19428
rect 26016 19388 26022 19400
rect 27430 19388 27436 19400
rect 27488 19388 27494 19440
rect 30282 19428 30288 19440
rect 30024 19400 30288 19428
rect 27154 19360 27160 19372
rect 23216 19332 27160 19360
rect 23017 19323 23075 19329
rect 3697 19295 3755 19301
rect 3697 19261 3709 19295
rect 3743 19292 3755 19295
rect 4706 19292 4712 19304
rect 3743 19264 4712 19292
rect 3743 19261 3755 19264
rect 3697 19255 3755 19261
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19292 5779 19295
rect 6914 19292 6920 19304
rect 5767 19264 6920 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 22922 19224 22928 19236
rect 992 19196 3556 19224
rect 16132 19196 22928 19224
rect 992 19184 998 19196
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 2188 19128 2237 19156
rect 2188 19116 2194 19128
rect 2225 19125 2237 19128
rect 2271 19125 2283 19159
rect 2225 19119 2283 19125
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5629 19159 5687 19165
rect 5629 19156 5641 19159
rect 5316 19128 5641 19156
rect 5316 19116 5322 19128
rect 5629 19125 5641 19128
rect 5675 19125 5687 19159
rect 5629 19119 5687 19125
rect 9490 19116 9496 19168
rect 9548 19156 9554 19168
rect 16132 19156 16160 19196
rect 22922 19184 22928 19196
rect 22980 19184 22986 19236
rect 9548 19128 16160 19156
rect 23032 19156 23060 19323
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 28902 19360 28908 19372
rect 27264 19332 28908 19360
rect 25590 19252 25596 19304
rect 25648 19292 25654 19304
rect 26237 19295 26295 19301
rect 26237 19292 26249 19295
rect 25648 19264 26249 19292
rect 25648 19252 25654 19264
rect 26237 19261 26249 19264
rect 26283 19261 26295 19295
rect 26237 19255 26295 19261
rect 26329 19295 26387 19301
rect 26329 19261 26341 19295
rect 26375 19261 26387 19295
rect 26329 19255 26387 19261
rect 26421 19295 26479 19301
rect 26421 19261 26433 19295
rect 26467 19261 26479 19295
rect 26421 19255 26479 19261
rect 24854 19184 24860 19236
rect 24912 19224 24918 19236
rect 25958 19224 25964 19236
rect 24912 19196 25964 19224
rect 24912 19184 24918 19196
rect 25958 19184 25964 19196
rect 26016 19224 26022 19236
rect 26344 19224 26372 19255
rect 26016 19196 26372 19224
rect 26436 19224 26464 19255
rect 26510 19252 26516 19304
rect 26568 19252 26574 19304
rect 27264 19292 27292 19332
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29178 19320 29184 19372
rect 29236 19320 29242 19372
rect 29362 19320 29368 19372
rect 29420 19320 29426 19372
rect 29822 19320 29828 19372
rect 29880 19369 29886 19372
rect 29880 19360 29890 19369
rect 30024 19360 30052 19400
rect 30282 19388 30288 19400
rect 30340 19388 30346 19440
rect 30374 19388 30380 19440
rect 30432 19428 30438 19440
rect 30432 19400 31754 19428
rect 30432 19388 30438 19400
rect 29880 19332 30052 19360
rect 30092 19363 30150 19369
rect 29880 19323 29890 19332
rect 30092 19329 30104 19363
rect 30138 19360 30150 19363
rect 31726 19360 31754 19400
rect 31938 19388 31944 19440
rect 31996 19428 32002 19440
rect 31996 19400 32536 19428
rect 31996 19388 32002 19400
rect 32508 19372 32536 19400
rect 32401 19363 32459 19369
rect 32401 19360 32413 19363
rect 30138 19332 31432 19360
rect 31726 19332 32413 19360
rect 30138 19329 30150 19332
rect 30092 19323 30150 19329
rect 29880 19320 29886 19323
rect 31404 19304 31432 19332
rect 32401 19329 32413 19332
rect 32447 19329 32459 19363
rect 32401 19323 32459 19329
rect 27080 19264 27292 19292
rect 27080 19224 27108 19264
rect 27338 19252 27344 19304
rect 27396 19252 27402 19304
rect 27430 19252 27436 19304
rect 27488 19252 27494 19304
rect 27522 19252 27528 19304
rect 27580 19252 27586 19304
rect 27614 19252 27620 19304
rect 27672 19252 27678 19304
rect 31386 19252 31392 19304
rect 31444 19252 31450 19304
rect 32416 19292 32444 19323
rect 32490 19320 32496 19372
rect 32548 19360 32554 19372
rect 32585 19363 32643 19369
rect 32585 19360 32597 19363
rect 32548 19332 32597 19360
rect 32548 19320 32554 19332
rect 32585 19329 32597 19332
rect 32631 19329 32643 19363
rect 32585 19323 32643 19329
rect 32692 19292 32720 19468
rect 34330 19428 34336 19440
rect 33980 19400 34336 19428
rect 32766 19320 32772 19372
rect 32824 19360 32830 19372
rect 33980 19369 34008 19400
rect 34330 19388 34336 19400
rect 34388 19388 34394 19440
rect 34992 19400 36676 19428
rect 33965 19363 34023 19369
rect 32824 19332 33916 19360
rect 32824 19320 32830 19332
rect 32416 19264 32720 19292
rect 26436 19196 27108 19224
rect 26016 19184 26022 19196
rect 27154 19184 27160 19236
rect 27212 19184 27218 19236
rect 27632 19224 27660 19252
rect 27448 19196 27660 19224
rect 23934 19156 23940 19168
rect 23032 19128 23940 19156
rect 9548 19116 9554 19128
rect 23934 19116 23940 19128
rect 23992 19116 23998 19168
rect 26510 19116 26516 19168
rect 26568 19156 26574 19168
rect 27448 19156 27476 19196
rect 31570 19184 31576 19236
rect 31628 19224 31634 19236
rect 33502 19224 33508 19236
rect 31628 19196 33508 19224
rect 31628 19184 31634 19196
rect 33502 19184 33508 19196
rect 33560 19184 33566 19236
rect 33888 19224 33916 19332
rect 33965 19329 33977 19363
rect 34011 19329 34023 19363
rect 33965 19323 34023 19329
rect 34149 19363 34207 19369
rect 34149 19329 34161 19363
rect 34195 19360 34207 19363
rect 34514 19360 34520 19372
rect 34195 19332 34520 19360
rect 34195 19329 34207 19332
rect 34149 19323 34207 19329
rect 34514 19320 34520 19332
rect 34572 19360 34578 19372
rect 34698 19360 34704 19372
rect 34572 19332 34704 19360
rect 34572 19320 34578 19332
rect 34698 19320 34704 19332
rect 34756 19320 34762 19372
rect 34992 19369 35020 19400
rect 34977 19363 35035 19369
rect 34977 19360 34989 19363
rect 34808 19332 34989 19360
rect 34241 19295 34299 19301
rect 34241 19261 34253 19295
rect 34287 19292 34299 19295
rect 34330 19292 34336 19304
rect 34287 19264 34336 19292
rect 34287 19261 34299 19264
rect 34241 19255 34299 19261
rect 34330 19252 34336 19264
rect 34388 19252 34394 19304
rect 34808 19292 34836 19332
rect 34977 19329 34989 19332
rect 35023 19329 35035 19363
rect 34977 19323 35035 19329
rect 35253 19363 35311 19369
rect 35253 19329 35265 19363
rect 35299 19360 35311 19363
rect 35434 19360 35440 19372
rect 35299 19332 35440 19360
rect 35299 19329 35311 19332
rect 35253 19323 35311 19329
rect 35434 19320 35440 19332
rect 35492 19320 35498 19372
rect 36262 19360 36268 19372
rect 35728 19332 36268 19360
rect 34440 19264 34836 19292
rect 35161 19295 35219 19301
rect 34440 19224 34468 19264
rect 35161 19261 35173 19295
rect 35207 19292 35219 19295
rect 35728 19292 35756 19332
rect 36262 19320 36268 19332
rect 36320 19320 36326 19372
rect 36648 19369 36676 19400
rect 37366 19388 37372 19440
rect 37424 19428 37430 19440
rect 37737 19431 37795 19437
rect 37737 19428 37749 19431
rect 37424 19400 37749 19428
rect 37424 19388 37430 19400
rect 37737 19397 37749 19400
rect 37783 19397 37795 19431
rect 37737 19391 37795 19397
rect 37829 19431 37887 19437
rect 37829 19397 37841 19431
rect 37875 19428 37887 19431
rect 38470 19428 38476 19440
rect 37875 19400 38476 19428
rect 37875 19397 37887 19400
rect 37829 19391 37887 19397
rect 38470 19388 38476 19400
rect 38528 19388 38534 19440
rect 42426 19428 42432 19440
rect 40972 19400 42432 19428
rect 36633 19363 36691 19369
rect 36633 19329 36645 19363
rect 36679 19360 36691 19363
rect 37274 19360 37280 19372
rect 36679 19332 37280 19360
rect 36679 19329 36691 19332
rect 36633 19323 36691 19329
rect 37274 19320 37280 19332
rect 37332 19320 37338 19372
rect 37642 19369 37648 19372
rect 37461 19363 37519 19369
rect 37461 19329 37473 19363
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 37609 19363 37648 19369
rect 37609 19329 37621 19363
rect 37609 19323 37648 19329
rect 35207 19264 35756 19292
rect 35805 19295 35863 19301
rect 35207 19261 35219 19264
rect 35161 19255 35219 19261
rect 35805 19261 35817 19295
rect 35851 19261 35863 19295
rect 37476 19292 37504 19323
rect 37642 19320 37648 19323
rect 37700 19320 37706 19372
rect 38010 19369 38016 19372
rect 37967 19363 38016 19369
rect 37967 19329 37979 19363
rect 38013 19329 38016 19363
rect 37967 19323 38016 19329
rect 38010 19320 38016 19323
rect 38068 19320 38074 19372
rect 38102 19320 38108 19372
rect 38160 19320 38166 19372
rect 40972 19369 41000 19400
rect 42426 19388 42432 19400
rect 42484 19388 42490 19440
rect 40957 19363 41015 19369
rect 38212 19332 40908 19360
rect 35805 19255 35863 19261
rect 37292 19264 37504 19292
rect 33888 19196 34468 19224
rect 34606 19184 34612 19236
rect 34664 19224 34670 19236
rect 35820 19224 35848 19255
rect 37292 19236 37320 19264
rect 34664 19196 35848 19224
rect 34664 19184 34670 19196
rect 36170 19184 36176 19236
rect 36228 19224 36234 19236
rect 36541 19227 36599 19233
rect 36541 19224 36553 19227
rect 36228 19196 36553 19224
rect 36228 19184 36234 19196
rect 36541 19193 36553 19196
rect 36587 19193 36599 19227
rect 36541 19187 36599 19193
rect 37274 19184 37280 19236
rect 37332 19184 37338 19236
rect 38120 19233 38148 19320
rect 38105 19227 38163 19233
rect 38105 19193 38117 19227
rect 38151 19193 38163 19227
rect 38105 19187 38163 19193
rect 26568 19128 27476 19156
rect 26568 19116 26574 19128
rect 27522 19116 27528 19168
rect 27580 19156 27586 19168
rect 31202 19156 31208 19168
rect 27580 19128 31208 19156
rect 27580 19116 27586 19128
rect 31202 19116 31208 19128
rect 31260 19116 31266 19168
rect 34793 19159 34851 19165
rect 34793 19125 34805 19159
rect 34839 19156 34851 19159
rect 37090 19156 37096 19168
rect 34839 19128 37096 19156
rect 34839 19125 34851 19128
rect 34793 19119 34851 19125
rect 37090 19116 37096 19128
rect 37148 19116 37154 19168
rect 37458 19116 37464 19168
rect 37516 19156 37522 19168
rect 38212 19156 38240 19332
rect 40880 19292 40908 19332
rect 40957 19329 40969 19363
rect 41003 19329 41015 19363
rect 41141 19363 41199 19369
rect 41141 19360 41153 19363
rect 40957 19323 41015 19329
rect 41064 19332 41153 19360
rect 41064 19292 41092 19332
rect 41141 19329 41153 19332
rect 41187 19360 41199 19363
rect 41598 19360 41604 19372
rect 41187 19332 41604 19360
rect 41187 19329 41199 19332
rect 41141 19323 41199 19329
rect 41598 19320 41604 19332
rect 41656 19320 41662 19372
rect 43088 19369 43116 19468
rect 44913 19465 44925 19499
rect 44959 19496 44971 19499
rect 45646 19496 45652 19508
rect 44959 19468 45652 19496
rect 44959 19465 44971 19468
rect 44913 19459 44971 19465
rect 45646 19456 45652 19468
rect 45704 19456 45710 19508
rect 45554 19428 45560 19440
rect 44744 19400 45560 19428
rect 43073 19363 43131 19369
rect 43073 19329 43085 19363
rect 43119 19329 43131 19363
rect 43073 19323 43131 19329
rect 43346 19320 43352 19372
rect 43404 19320 43410 19372
rect 43898 19320 43904 19372
rect 43956 19320 43962 19372
rect 44085 19363 44143 19369
rect 44085 19329 44097 19363
rect 44131 19360 44143 19363
rect 44174 19360 44180 19372
rect 44131 19332 44180 19360
rect 44131 19329 44143 19332
rect 44085 19323 44143 19329
rect 44174 19320 44180 19332
rect 44232 19320 44238 19372
rect 44744 19369 44772 19400
rect 45554 19388 45560 19400
rect 45612 19388 45618 19440
rect 44729 19363 44787 19369
rect 44729 19329 44741 19363
rect 44775 19329 44787 19363
rect 44729 19323 44787 19329
rect 44913 19363 44971 19369
rect 44913 19329 44925 19363
rect 44959 19329 44971 19363
rect 44913 19323 44971 19329
rect 40880 19264 41092 19292
rect 42886 19252 42892 19304
rect 42944 19252 42950 19304
rect 43165 19295 43223 19301
rect 43165 19261 43177 19295
rect 43211 19292 43223 19295
rect 43993 19295 44051 19301
rect 43993 19292 44005 19295
rect 43211 19264 44005 19292
rect 43211 19261 43223 19264
rect 43165 19255 43223 19261
rect 43993 19261 44005 19264
rect 44039 19261 44051 19295
rect 43993 19255 44051 19261
rect 44450 19252 44456 19304
rect 44508 19292 44514 19304
rect 44928 19292 44956 19323
rect 44508 19264 44956 19292
rect 44508 19252 44514 19264
rect 43257 19227 43315 19233
rect 43257 19193 43269 19227
rect 43303 19224 43315 19227
rect 45922 19224 45928 19236
rect 43303 19196 45928 19224
rect 43303 19193 43315 19196
rect 43257 19187 43315 19193
rect 45922 19184 45928 19196
rect 45980 19184 45986 19236
rect 37516 19128 38240 19156
rect 37516 19116 37522 19128
rect 40954 19116 40960 19168
rect 41012 19116 41018 19168
rect 42794 19116 42800 19168
rect 42852 19156 42858 19168
rect 43898 19156 43904 19168
rect 42852 19128 43904 19156
rect 42852 19116 42858 19128
rect 43898 19116 43904 19128
rect 43956 19116 43962 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 3234 18912 3240 18964
rect 3292 18912 3298 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 6549 18955 6607 18961
rect 4120 18924 6500 18952
rect 4120 18912 4126 18924
rect 6472 18884 6500 18924
rect 6549 18921 6561 18955
rect 6595 18952 6607 18955
rect 6730 18952 6736 18964
rect 6595 18924 6736 18952
rect 6595 18921 6607 18924
rect 6549 18915 6607 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 9582 18912 9588 18964
rect 9640 18952 9646 18964
rect 9950 18952 9956 18964
rect 9640 18924 9956 18952
rect 9640 18912 9646 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10134 18912 10140 18964
rect 10192 18912 10198 18964
rect 11517 18955 11575 18961
rect 11517 18921 11529 18955
rect 11563 18952 11575 18955
rect 11698 18952 11704 18964
rect 11563 18924 11704 18952
rect 11563 18921 11575 18924
rect 11517 18915 11575 18921
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 13354 18952 13360 18964
rect 12492 18924 13360 18952
rect 12492 18912 12498 18924
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 22428 18924 22569 18952
rect 22428 18912 22434 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 22557 18915 22615 18921
rect 26142 18912 26148 18964
rect 26200 18952 26206 18964
rect 26200 18924 28948 18952
rect 26200 18912 26206 18924
rect 9766 18884 9772 18896
rect 6472 18856 9772 18884
rect 9766 18844 9772 18856
rect 9824 18844 9830 18896
rect 20162 18884 20168 18896
rect 9876 18856 20168 18884
rect 6822 18776 6828 18828
rect 6880 18816 6886 18828
rect 6880 18776 6914 18816
rect 1762 18708 1768 18760
rect 1820 18748 1826 18760
rect 2130 18757 2136 18760
rect 1857 18751 1915 18757
rect 1857 18748 1869 18751
rect 1820 18720 1869 18748
rect 1820 18708 1826 18720
rect 1857 18717 1869 18720
rect 1903 18717 1915 18751
rect 2124 18748 2136 18757
rect 2091 18720 2136 18748
rect 1857 18711 1915 18717
rect 2124 18711 2136 18720
rect 2130 18708 2136 18711
rect 2188 18708 2194 18760
rect 5166 18708 5172 18760
rect 5224 18708 5230 18760
rect 5436 18751 5494 18757
rect 5436 18717 5448 18751
rect 5482 18748 5494 18751
rect 6362 18748 6368 18760
rect 5482 18720 6368 18748
rect 5482 18717 5494 18720
rect 5436 18711 5494 18717
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 5902 18640 5908 18692
rect 5960 18680 5966 18692
rect 6886 18680 6914 18776
rect 7926 18708 7932 18760
rect 7984 18748 7990 18760
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 7984 18720 9505 18748
rect 7984 18708 7990 18720
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 9641 18751 9699 18757
rect 9641 18717 9653 18751
rect 9687 18748 9699 18751
rect 9876 18748 9904 18856
rect 20162 18844 20168 18856
rect 20220 18844 20226 18896
rect 20625 18887 20683 18893
rect 20625 18853 20637 18887
rect 20671 18884 20683 18887
rect 22278 18884 22284 18896
rect 20671 18856 22284 18884
rect 20671 18853 20683 18856
rect 20625 18847 20683 18853
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 12897 18819 12955 18825
rect 12897 18816 12909 18819
rect 11480 18788 12909 18816
rect 11480 18776 11486 18788
rect 12897 18785 12909 18788
rect 12943 18785 12955 18819
rect 20640 18816 20668 18847
rect 22278 18844 22284 18856
rect 22336 18884 22342 18896
rect 22646 18884 22652 18896
rect 22336 18856 22652 18884
rect 22336 18844 22342 18856
rect 22646 18844 22652 18856
rect 22704 18844 22710 18896
rect 26418 18844 26424 18896
rect 26476 18844 26482 18896
rect 26970 18884 26976 18896
rect 26528 18856 26976 18884
rect 12897 18779 12955 18785
rect 13096 18788 19472 18816
rect 9687 18720 9904 18748
rect 9687 18717 9699 18720
rect 9641 18711 9699 18717
rect 9950 18708 9956 18760
rect 10008 18757 10014 18760
rect 10008 18748 10016 18757
rect 10008 18720 10053 18748
rect 10008 18711 10016 18720
rect 10008 18708 10014 18711
rect 11790 18708 11796 18760
rect 11848 18708 11854 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 13096 18748 13124 18788
rect 11940 18720 13124 18748
rect 13173 18751 13231 18757
rect 11940 18708 11946 18720
rect 13173 18717 13185 18751
rect 13219 18748 13231 18751
rect 16390 18748 16396 18760
rect 13219 18720 16396 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 9769 18683 9827 18689
rect 9769 18680 9781 18683
rect 5960 18652 9781 18680
rect 5960 18640 5966 18652
rect 9769 18649 9781 18652
rect 9815 18649 9827 18683
rect 9769 18643 9827 18649
rect 9784 18612 9812 18643
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 11698 18640 11704 18692
rect 11756 18640 11762 18692
rect 12253 18683 12311 18689
rect 12253 18649 12265 18683
rect 12299 18649 12311 18683
rect 12253 18643 12311 18649
rect 12158 18612 12164 18624
rect 9784 18584 12164 18612
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 12268 18612 12296 18643
rect 12894 18640 12900 18692
rect 12952 18680 12958 18692
rect 13081 18683 13139 18689
rect 13081 18680 13093 18683
rect 12952 18652 13093 18680
rect 12952 18640 12958 18652
rect 13081 18649 13093 18652
rect 13127 18649 13139 18683
rect 13081 18643 13139 18649
rect 19334 18612 19340 18624
rect 12268 18584 19340 18612
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 19444 18612 19472 18788
rect 19536 18788 20668 18816
rect 21177 18819 21235 18825
rect 19536 18757 19564 18788
rect 21177 18785 21189 18819
rect 21223 18816 21235 18819
rect 22741 18819 22799 18825
rect 22741 18816 22753 18819
rect 21223 18788 22753 18816
rect 21223 18785 21235 18788
rect 21177 18779 21235 18785
rect 22741 18785 22753 18788
rect 22787 18785 22799 18819
rect 22741 18779 22799 18785
rect 22925 18819 22983 18825
rect 22925 18785 22937 18819
rect 22971 18816 22983 18819
rect 23658 18816 23664 18828
rect 22971 18788 23664 18816
rect 22971 18785 22983 18788
rect 22925 18779 22983 18785
rect 23658 18776 23664 18788
rect 23716 18776 23722 18828
rect 24762 18776 24768 18828
rect 24820 18816 24826 18828
rect 25590 18816 25596 18828
rect 24820 18788 25596 18816
rect 24820 18776 24826 18788
rect 25590 18776 25596 18788
rect 25648 18816 25654 18828
rect 26528 18816 26556 18856
rect 26970 18844 26976 18856
rect 27028 18884 27034 18896
rect 27338 18884 27344 18896
rect 27028 18856 27344 18884
rect 27028 18844 27034 18856
rect 27338 18844 27344 18856
rect 27396 18844 27402 18896
rect 28920 18884 28948 18924
rect 31386 18912 31392 18964
rect 31444 18912 31450 18964
rect 32582 18912 32588 18964
rect 32640 18952 32646 18964
rect 32640 18924 42932 18952
rect 32640 18912 32646 18924
rect 28920 18856 36492 18884
rect 25648 18788 26556 18816
rect 26605 18819 26663 18825
rect 25648 18776 25654 18788
rect 26605 18785 26617 18819
rect 26651 18816 26663 18819
rect 27154 18816 27160 18828
rect 26651 18788 27160 18816
rect 26651 18785 26663 18788
rect 26605 18779 26663 18785
rect 27154 18776 27160 18788
rect 27212 18776 27218 18828
rect 30098 18776 30104 18828
rect 30156 18816 30162 18828
rect 36464 18816 36492 18856
rect 42426 18844 42432 18896
rect 42484 18844 42490 18896
rect 42705 18887 42763 18893
rect 42705 18853 42717 18887
rect 42751 18884 42763 18887
rect 42794 18884 42800 18896
rect 42751 18856 42800 18884
rect 42751 18853 42763 18856
rect 42705 18847 42763 18853
rect 42794 18844 42800 18856
rect 42852 18844 42858 18896
rect 30156 18788 34836 18816
rect 36464 18788 40356 18816
rect 30156 18776 30162 18788
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18748 19855 18751
rect 20070 18748 20076 18760
rect 19843 18720 20076 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 20070 18708 20076 18720
rect 20128 18708 20134 18760
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18748 20499 18751
rect 20898 18748 20904 18760
rect 20487 18720 20904 18748
rect 20487 18717 20499 18720
rect 20441 18711 20499 18717
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 21048 18720 21373 18748
rect 21048 18708 21054 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 21450 18708 21456 18760
rect 21508 18708 21514 18760
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 21637 18751 21695 18757
rect 21637 18717 21649 18751
rect 21683 18748 21695 18751
rect 21726 18748 21732 18760
rect 21683 18720 21732 18748
rect 21683 18717 21695 18720
rect 21637 18711 21695 18717
rect 19978 18640 19984 18692
rect 20036 18680 20042 18692
rect 21560 18680 21588 18711
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 22830 18708 22836 18760
rect 22888 18708 22894 18760
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18748 23075 18751
rect 23290 18748 23296 18760
rect 23063 18720 23296 18748
rect 23063 18717 23075 18720
rect 23017 18711 23075 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 24854 18748 24860 18760
rect 24688 18720 24860 18748
rect 24688 18680 24716 18720
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 26694 18708 26700 18760
rect 26752 18708 26758 18760
rect 26789 18751 26847 18757
rect 26789 18717 26801 18751
rect 26835 18717 26847 18751
rect 26789 18711 26847 18717
rect 20036 18652 21588 18680
rect 21652 18652 24716 18680
rect 20036 18640 20042 18652
rect 20714 18612 20720 18624
rect 19444 18584 20720 18612
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 21450 18572 21456 18624
rect 21508 18612 21514 18624
rect 21652 18612 21680 18652
rect 24762 18640 24768 18692
rect 24820 18680 24826 18692
rect 26326 18680 26332 18692
rect 24820 18652 26332 18680
rect 24820 18640 24826 18652
rect 26326 18640 26332 18652
rect 26384 18680 26390 18692
rect 26804 18680 26832 18711
rect 26878 18708 26884 18760
rect 26936 18708 26942 18760
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 31018 18748 31024 18760
rect 28776 18720 31024 18748
rect 28776 18708 28782 18720
rect 31018 18708 31024 18720
rect 31076 18708 31082 18760
rect 31110 18708 31116 18760
rect 31168 18748 31174 18760
rect 31570 18748 31576 18760
rect 31168 18720 31576 18748
rect 31168 18708 31174 18720
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 31665 18751 31723 18757
rect 31665 18717 31677 18751
rect 31711 18748 31723 18751
rect 32582 18748 32588 18760
rect 31711 18720 32588 18748
rect 31711 18717 31723 18720
rect 31665 18711 31723 18717
rect 32582 18708 32588 18720
rect 32640 18708 32646 18760
rect 34808 18748 34836 18788
rect 36354 18748 36360 18760
rect 34808 18720 36360 18748
rect 36354 18708 36360 18720
rect 36412 18708 36418 18760
rect 37458 18708 37464 18760
rect 37516 18748 37522 18760
rect 37642 18748 37648 18760
rect 37516 18720 37648 18748
rect 37516 18708 37522 18720
rect 37642 18708 37648 18720
rect 37700 18708 37706 18760
rect 40221 18751 40279 18757
rect 40221 18717 40233 18751
rect 40267 18717 40279 18751
rect 40328 18748 40356 18788
rect 41322 18776 41328 18828
rect 41380 18816 41386 18828
rect 41380 18788 42288 18816
rect 41380 18776 41386 18788
rect 40488 18751 40546 18757
rect 40328 18720 40448 18748
rect 40221 18711 40279 18717
rect 26384 18652 26832 18680
rect 30009 18683 30067 18689
rect 26384 18640 26390 18652
rect 30009 18649 30021 18683
rect 30055 18680 30067 18683
rect 30098 18680 30104 18692
rect 30055 18652 30104 18680
rect 30055 18649 30067 18652
rect 30009 18643 30067 18649
rect 30098 18640 30104 18652
rect 30156 18640 30162 18692
rect 30374 18640 30380 18692
rect 30432 18680 30438 18692
rect 30745 18683 30803 18689
rect 30745 18680 30757 18683
rect 30432 18652 30757 18680
rect 30432 18640 30438 18652
rect 30745 18649 30757 18652
rect 30791 18649 30803 18683
rect 30745 18643 30803 18649
rect 31202 18640 31208 18692
rect 31260 18680 31266 18692
rect 31941 18683 31999 18689
rect 31941 18680 31953 18683
rect 31260 18652 31953 18680
rect 31260 18640 31266 18652
rect 31941 18649 31953 18652
rect 31987 18649 31999 18683
rect 31941 18643 31999 18649
rect 32030 18640 32036 18692
rect 32088 18680 32094 18692
rect 34790 18680 34796 18692
rect 32088 18652 34796 18680
rect 32088 18640 32094 18652
rect 34790 18640 34796 18652
rect 34848 18640 34854 18692
rect 36538 18640 36544 18692
rect 36596 18680 36602 18692
rect 37093 18683 37151 18689
rect 37093 18680 37105 18683
rect 36596 18652 37105 18680
rect 36596 18640 36602 18652
rect 37093 18649 37105 18652
rect 37139 18680 37151 18683
rect 40236 18680 40264 18711
rect 40310 18680 40316 18692
rect 37139 18652 40316 18680
rect 37139 18649 37151 18652
rect 37093 18643 37151 18649
rect 40310 18640 40316 18652
rect 40368 18640 40374 18692
rect 40420 18680 40448 18720
rect 40488 18717 40500 18751
rect 40534 18748 40546 18751
rect 40954 18748 40960 18760
rect 40534 18720 40960 18748
rect 40534 18717 40546 18720
rect 40488 18711 40546 18717
rect 40954 18708 40960 18720
rect 41012 18708 41018 18760
rect 42150 18680 42156 18692
rect 40420 18652 42156 18680
rect 42150 18640 42156 18652
rect 42208 18640 42214 18692
rect 21508 18584 21680 18612
rect 21508 18572 21514 18584
rect 25866 18572 25872 18624
rect 25924 18612 25930 18624
rect 40586 18612 40592 18624
rect 25924 18584 40592 18612
rect 25924 18572 25930 18584
rect 40586 18572 40592 18584
rect 40644 18572 40650 18624
rect 41598 18572 41604 18624
rect 41656 18572 41662 18624
rect 42260 18612 42288 18788
rect 42334 18708 42340 18760
rect 42392 18748 42398 18760
rect 42904 18757 42932 18924
rect 44450 18912 44456 18964
rect 44508 18952 44514 18964
rect 44508 18924 45416 18952
rect 44508 18912 44514 18924
rect 43898 18844 43904 18896
rect 43956 18884 43962 18896
rect 44637 18887 44695 18893
rect 44637 18884 44649 18887
rect 43956 18856 44649 18884
rect 43956 18844 43962 18856
rect 44637 18853 44649 18856
rect 44683 18853 44695 18887
rect 44637 18847 44695 18853
rect 44174 18776 44180 18828
rect 44232 18816 44238 18828
rect 45189 18819 45247 18825
rect 45189 18816 45201 18819
rect 44232 18788 45201 18816
rect 44232 18776 44238 18788
rect 45189 18785 45201 18788
rect 45235 18785 45247 18819
rect 45388 18816 45416 18924
rect 45388 18788 45508 18816
rect 45189 18779 45247 18785
rect 45480 18757 45508 18788
rect 45922 18776 45928 18828
rect 45980 18776 45986 18828
rect 42613 18751 42671 18757
rect 42613 18748 42625 18751
rect 42392 18720 42625 18748
rect 42392 18708 42398 18720
rect 42613 18717 42625 18720
rect 42659 18717 42671 18751
rect 42613 18711 42671 18717
rect 42797 18751 42855 18757
rect 42797 18717 42809 18751
rect 42843 18717 42855 18751
rect 42797 18711 42855 18717
rect 42889 18751 42947 18757
rect 42889 18717 42901 18751
rect 42935 18717 42947 18751
rect 45373 18751 45431 18757
rect 45373 18748 45385 18751
rect 42889 18711 42947 18717
rect 44284 18720 45385 18748
rect 42812 18680 42840 18711
rect 44284 18692 44312 18720
rect 45373 18717 45385 18720
rect 45419 18717 45431 18751
rect 45373 18711 45431 18717
rect 45465 18751 45523 18757
rect 45465 18717 45477 18751
rect 45511 18717 45523 18751
rect 45465 18711 45523 18717
rect 44174 18680 44180 18692
rect 42812 18652 44180 18680
rect 44174 18640 44180 18652
rect 44232 18640 44238 18692
rect 44266 18640 44272 18692
rect 44324 18640 44330 18692
rect 44485 18683 44543 18689
rect 44485 18649 44497 18683
rect 44531 18680 44543 18683
rect 45554 18680 45560 18692
rect 44531 18652 45560 18680
rect 44531 18649 44543 18652
rect 44485 18643 44543 18649
rect 45554 18640 45560 18652
rect 45612 18640 45618 18692
rect 43714 18612 43720 18624
rect 42260 18584 43720 18612
rect 43714 18572 43720 18584
rect 43772 18572 43778 18624
rect 43806 18572 43812 18624
rect 43864 18612 43870 18624
rect 45738 18612 45744 18624
rect 43864 18584 45744 18612
rect 43864 18572 43870 18584
rect 45738 18572 45744 18584
rect 45796 18572 45802 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1026 18368 1032 18420
rect 1084 18408 1090 18420
rect 1084 18380 2636 18408
rect 1084 18368 1090 18380
rect 934 18300 940 18352
rect 992 18340 998 18352
rect 2608 18349 2636 18380
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 11698 18408 11704 18420
rect 2832 18380 11704 18408
rect 2832 18368 2838 18380
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 19705 18411 19763 18417
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 19978 18408 19984 18420
rect 19751 18380 19984 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 22186 18408 22192 18420
rect 21560 18380 22192 18408
rect 1857 18343 1915 18349
rect 1857 18340 1869 18343
rect 992 18312 1869 18340
rect 992 18300 998 18312
rect 1857 18309 1869 18312
rect 1903 18309 1915 18343
rect 1857 18303 1915 18309
rect 2593 18343 2651 18349
rect 2593 18309 2605 18343
rect 2639 18309 2651 18343
rect 2593 18303 2651 18309
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 21450 18340 21456 18352
rect 3476 18312 21456 18340
rect 3476 18300 3482 18312
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 1627 18244 2544 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2516 18204 2544 18244
rect 14734 18232 14740 18284
rect 14792 18272 14798 18284
rect 14792 18244 16988 18272
rect 14792 18232 14798 18244
rect 15010 18204 15016 18216
rect 2516 18176 15016 18204
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 16666 18164 16672 18216
rect 16724 18204 16730 18216
rect 16850 18204 16856 18216
rect 16724 18176 16856 18204
rect 16724 18164 16730 18176
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 16960 18204 16988 18244
rect 17034 18232 17040 18284
rect 17092 18232 17098 18284
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 17184 18244 17233 18272
rect 17184 18232 17190 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 18592 18275 18650 18281
rect 18592 18241 18604 18275
rect 18638 18272 18650 18275
rect 19426 18272 19432 18284
rect 18638 18244 19432 18272
rect 18638 18241 18650 18244
rect 18592 18235 18650 18241
rect 17328 18204 17356 18235
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 16960 18176 17448 18204
rect 2774 18096 2780 18148
rect 2832 18096 2838 18148
rect 9766 18096 9772 18148
rect 9824 18136 9830 18148
rect 17218 18136 17224 18148
rect 9824 18108 17224 18136
rect 9824 18096 9830 18108
rect 17218 18096 17224 18108
rect 17276 18096 17282 18148
rect 16850 18028 16856 18080
rect 16908 18028 16914 18080
rect 17420 18068 17448 18176
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 18012 18176 18337 18204
rect 18012 18164 18018 18176
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 18325 18167 18383 18173
rect 21560 18136 21588 18380
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 22922 18368 22928 18420
rect 22980 18408 22986 18420
rect 24397 18411 24455 18417
rect 24397 18408 24409 18411
rect 22980 18380 24409 18408
rect 22980 18368 22986 18380
rect 24397 18377 24409 18380
rect 24443 18377 24455 18411
rect 24397 18371 24455 18377
rect 25038 18368 25044 18420
rect 25096 18408 25102 18420
rect 25866 18408 25872 18420
rect 25096 18380 25872 18408
rect 25096 18368 25102 18380
rect 25866 18368 25872 18380
rect 25924 18408 25930 18420
rect 26510 18408 26516 18420
rect 25924 18380 26516 18408
rect 25924 18368 25930 18380
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 26694 18368 26700 18420
rect 26752 18408 26758 18420
rect 40494 18408 40500 18420
rect 26752 18380 40500 18408
rect 26752 18368 26758 18380
rect 40494 18368 40500 18380
rect 40552 18368 40558 18420
rect 40586 18368 40592 18420
rect 40644 18368 40650 18420
rect 42150 18368 42156 18420
rect 42208 18408 42214 18420
rect 43901 18411 43959 18417
rect 43901 18408 43913 18411
rect 42208 18380 43913 18408
rect 42208 18368 42214 18380
rect 43901 18377 43913 18380
rect 43947 18377 43959 18411
rect 43901 18371 43959 18377
rect 44450 18368 44456 18420
rect 44508 18408 44514 18420
rect 44637 18411 44695 18417
rect 44637 18408 44649 18411
rect 44508 18380 44649 18408
rect 44508 18368 44514 18380
rect 44637 18377 44649 18380
rect 44683 18377 44695 18411
rect 44637 18371 44695 18377
rect 23934 18340 23940 18352
rect 22020 18312 23940 18340
rect 22020 18281 22048 18312
rect 23934 18300 23940 18312
rect 23992 18300 23998 18352
rect 32674 18340 32680 18352
rect 24780 18312 31754 18340
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22261 18275 22319 18281
rect 22261 18272 22273 18275
rect 22152 18244 22273 18272
rect 22152 18232 22158 18244
rect 22261 18241 22273 18244
rect 22307 18241 22319 18275
rect 22261 18235 22319 18241
rect 24673 18275 24731 18281
rect 24673 18241 24685 18275
rect 24719 18272 24731 18275
rect 24780 18272 24808 18312
rect 24719 18244 24808 18272
rect 24719 18241 24731 18244
rect 24673 18235 24731 18241
rect 24854 18232 24860 18284
rect 24912 18232 24918 18284
rect 24946 18232 24952 18284
rect 25004 18272 25010 18284
rect 25682 18272 25688 18284
rect 25004 18244 25688 18272
rect 25004 18232 25010 18244
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 25777 18275 25835 18281
rect 25777 18241 25789 18275
rect 25823 18272 25835 18275
rect 30466 18272 30472 18284
rect 25823 18244 30472 18272
rect 25823 18241 25835 18244
rect 25777 18235 25835 18241
rect 30466 18232 30472 18244
rect 30524 18232 30530 18284
rect 30650 18281 30656 18284
rect 30644 18235 30656 18281
rect 30650 18232 30656 18235
rect 30708 18232 30714 18284
rect 31018 18232 31024 18284
rect 31076 18272 31082 18284
rect 31570 18272 31576 18284
rect 31076 18244 31576 18272
rect 31076 18232 31082 18244
rect 31570 18232 31576 18244
rect 31628 18232 31634 18284
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 19306 18108 21588 18136
rect 24596 18136 24624 18167
rect 24762 18164 24768 18216
rect 24820 18164 24826 18216
rect 24872 18204 24900 18232
rect 24872 18176 25544 18204
rect 25409 18139 25467 18145
rect 25409 18136 25421 18139
rect 24596 18108 25421 18136
rect 19306 18068 19334 18108
rect 25409 18105 25421 18108
rect 25455 18105 25467 18139
rect 25516 18136 25544 18176
rect 25590 18164 25596 18216
rect 25648 18164 25654 18216
rect 25866 18164 25872 18216
rect 25924 18164 25930 18216
rect 30374 18164 30380 18216
rect 30432 18164 30438 18216
rect 31726 18204 31754 18312
rect 32416 18312 32680 18340
rect 32416 18281 32444 18312
rect 32674 18300 32680 18312
rect 32732 18300 32738 18352
rect 37274 18300 37280 18352
rect 37332 18340 37338 18352
rect 40313 18343 40371 18349
rect 37332 18312 39988 18340
rect 37332 18300 37338 18312
rect 32401 18275 32459 18281
rect 32401 18241 32413 18275
rect 32447 18241 32459 18275
rect 32401 18235 32459 18241
rect 32585 18275 32643 18281
rect 32585 18241 32597 18275
rect 32631 18272 32643 18275
rect 32766 18272 32772 18284
rect 32631 18244 32772 18272
rect 32631 18241 32643 18244
rect 32585 18235 32643 18241
rect 32766 18232 32772 18244
rect 32824 18232 32830 18284
rect 37458 18232 37464 18284
rect 37516 18232 37522 18284
rect 37642 18232 37648 18284
rect 37700 18232 37706 18284
rect 39960 18281 39988 18312
rect 40313 18309 40325 18343
rect 40359 18340 40371 18343
rect 41230 18340 41236 18352
rect 40359 18312 41236 18340
rect 40359 18309 40371 18312
rect 40313 18303 40371 18309
rect 41230 18300 41236 18312
rect 41288 18300 41294 18352
rect 43070 18300 43076 18352
rect 43128 18340 43134 18352
rect 43625 18343 43683 18349
rect 43625 18340 43637 18343
rect 43128 18312 43637 18340
rect 43128 18300 43134 18312
rect 43625 18309 43637 18312
rect 43671 18309 43683 18343
rect 45554 18340 45560 18352
rect 43625 18303 43683 18309
rect 44008 18312 45560 18340
rect 39945 18275 40003 18281
rect 39945 18241 39957 18275
rect 39991 18241 40003 18275
rect 39945 18235 40003 18241
rect 40093 18275 40151 18281
rect 40093 18241 40105 18275
rect 40139 18272 40151 18275
rect 40139 18241 40172 18272
rect 40093 18235 40172 18241
rect 34146 18204 34152 18216
rect 31726 18176 34152 18204
rect 34146 18164 34152 18176
rect 34204 18164 34210 18216
rect 36446 18164 36452 18216
rect 36504 18204 36510 18216
rect 37660 18204 37688 18232
rect 36504 18176 37688 18204
rect 36504 18164 36510 18176
rect 26878 18136 26884 18148
rect 25516 18108 26884 18136
rect 25409 18099 25467 18105
rect 26878 18096 26884 18108
rect 26936 18096 26942 18148
rect 31386 18096 31392 18148
rect 31444 18136 31450 18148
rect 32401 18139 32459 18145
rect 32401 18136 32413 18139
rect 31444 18108 32413 18136
rect 31444 18096 31450 18108
rect 32401 18105 32413 18108
rect 32447 18105 32459 18139
rect 38102 18136 38108 18148
rect 32401 18099 32459 18105
rect 37200 18108 38108 18136
rect 17420 18040 19334 18068
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 22002 18068 22008 18080
rect 20772 18040 22008 18068
rect 20772 18028 20778 18040
rect 22002 18028 22008 18040
rect 22060 18068 22066 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 22060 18040 23397 18068
rect 22060 18028 22066 18040
rect 23385 18037 23397 18040
rect 23431 18037 23443 18071
rect 23385 18031 23443 18037
rect 23658 18028 23664 18080
rect 23716 18068 23722 18080
rect 24762 18068 24768 18080
rect 23716 18040 24768 18068
rect 23716 18028 23722 18040
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 31294 18028 31300 18080
rect 31352 18068 31358 18080
rect 31757 18071 31815 18077
rect 31757 18068 31769 18071
rect 31352 18040 31769 18068
rect 31352 18028 31358 18040
rect 31757 18037 31769 18040
rect 31803 18037 31815 18071
rect 31757 18031 31815 18037
rect 31846 18028 31852 18080
rect 31904 18068 31910 18080
rect 37200 18068 37228 18108
rect 38102 18096 38108 18108
rect 38160 18096 38166 18148
rect 39960 18136 39988 18235
rect 40144 18204 40172 18235
rect 40218 18232 40224 18284
rect 40276 18232 40282 18284
rect 40451 18275 40509 18281
rect 40451 18241 40463 18275
rect 40497 18272 40509 18275
rect 40586 18272 40592 18284
rect 40497 18244 40592 18272
rect 40497 18241 40509 18244
rect 40451 18235 40509 18241
rect 40586 18232 40592 18244
rect 40644 18272 40650 18284
rect 41322 18272 41328 18284
rect 40644 18244 41328 18272
rect 40644 18232 40650 18244
rect 41322 18232 41328 18244
rect 41380 18232 41386 18284
rect 41506 18232 41512 18284
rect 41564 18272 41570 18284
rect 41564 18244 43208 18272
rect 41564 18232 41570 18244
rect 42058 18204 42064 18216
rect 40144 18176 42064 18204
rect 42058 18164 42064 18176
rect 42116 18164 42122 18216
rect 43180 18204 43208 18244
rect 43254 18232 43260 18284
rect 43312 18232 43318 18284
rect 43438 18281 43444 18284
rect 43405 18275 43444 18281
rect 43405 18241 43417 18275
rect 43405 18235 43444 18241
rect 43438 18232 43444 18235
rect 43496 18232 43502 18284
rect 43530 18232 43536 18284
rect 43588 18232 43594 18284
rect 43714 18232 43720 18284
rect 43772 18281 43778 18284
rect 43772 18272 43780 18281
rect 43772 18244 43817 18272
rect 43772 18235 43780 18244
rect 43772 18232 43778 18235
rect 44008 18204 44036 18312
rect 44744 18281 44772 18312
rect 45554 18300 45560 18312
rect 45612 18300 45618 18352
rect 44453 18275 44511 18281
rect 44453 18241 44465 18275
rect 44499 18241 44511 18275
rect 44453 18235 44511 18241
rect 44729 18275 44787 18281
rect 44729 18241 44741 18275
rect 44775 18241 44787 18275
rect 44729 18235 44787 18241
rect 44266 18204 44272 18216
rect 43180 18176 44036 18204
rect 44100 18176 44272 18204
rect 40034 18136 40040 18148
rect 39960 18108 40040 18136
rect 40034 18096 40040 18108
rect 40092 18136 40098 18148
rect 43254 18136 43260 18148
rect 40092 18108 43260 18136
rect 40092 18096 40098 18108
rect 43254 18096 43260 18108
rect 43312 18096 43318 18148
rect 31904 18040 37228 18068
rect 31904 18028 31910 18040
rect 37274 18028 37280 18080
rect 37332 18068 37338 18080
rect 37461 18071 37519 18077
rect 37461 18068 37473 18071
rect 37332 18040 37473 18068
rect 37332 18028 37338 18040
rect 37461 18037 37473 18040
rect 37507 18037 37519 18071
rect 37461 18031 37519 18037
rect 38654 18028 38660 18080
rect 38712 18068 38718 18080
rect 41506 18068 41512 18080
rect 38712 18040 41512 18068
rect 38712 18028 38718 18040
rect 41506 18028 41512 18040
rect 41564 18028 41570 18080
rect 41598 18028 41604 18080
rect 41656 18068 41662 18080
rect 44100 18068 44128 18176
rect 44266 18164 44272 18176
rect 44324 18204 44330 18216
rect 44468 18204 44496 18235
rect 44324 18176 44496 18204
rect 44324 18164 44330 18176
rect 44174 18096 44180 18148
rect 44232 18136 44238 18148
rect 44453 18139 44511 18145
rect 44453 18136 44465 18139
rect 44232 18108 44465 18136
rect 44232 18096 44238 18108
rect 44453 18105 44465 18108
rect 44499 18105 44511 18139
rect 44453 18099 44511 18105
rect 41656 18040 44128 18068
rect 41656 18028 41662 18040
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 5166 17864 5172 17876
rect 3988 17836 5172 17864
rect 1762 17688 1768 17740
rect 1820 17728 1826 17740
rect 3988 17737 4016 17836
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 5350 17824 5356 17876
rect 5408 17824 5414 17876
rect 17126 17864 17132 17876
rect 6886 17836 17132 17864
rect 6886 17796 6914 17836
rect 17126 17824 17132 17836
rect 17184 17864 17190 17876
rect 17773 17867 17831 17873
rect 17773 17864 17785 17867
rect 17184 17836 17785 17864
rect 17184 17824 17190 17836
rect 17773 17833 17785 17836
rect 17819 17833 17831 17867
rect 17773 17827 17831 17833
rect 19426 17824 19432 17876
rect 19484 17824 19490 17876
rect 21637 17867 21695 17873
rect 21637 17833 21649 17867
rect 21683 17864 21695 17867
rect 22094 17864 22100 17876
rect 21683 17836 22100 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 22830 17824 22836 17876
rect 22888 17864 22894 17876
rect 27614 17864 27620 17876
rect 22888 17836 27620 17864
rect 22888 17824 22894 17836
rect 27614 17824 27620 17836
rect 27672 17824 27678 17876
rect 30650 17824 30656 17876
rect 30708 17824 30714 17876
rect 35713 17867 35771 17873
rect 35713 17864 35725 17867
rect 31726 17836 35725 17864
rect 5092 17768 6914 17796
rect 3973 17731 4031 17737
rect 3973 17728 3985 17731
rect 1820 17700 3985 17728
rect 1820 17688 1826 17700
rect 3973 17697 3985 17700
rect 4019 17697 4031 17731
rect 3973 17691 4031 17697
rect 934 17620 940 17672
rect 992 17660 998 17672
rect 2501 17663 2559 17669
rect 992 17632 1808 17660
rect 992 17620 998 17632
rect 1118 17552 1124 17604
rect 1176 17592 1182 17604
rect 1673 17595 1731 17601
rect 1673 17592 1685 17595
rect 1176 17564 1685 17592
rect 1176 17552 1182 17564
rect 1673 17561 1685 17564
rect 1719 17561 1731 17595
rect 1780 17592 1808 17632
rect 2501 17629 2513 17663
rect 2547 17660 2559 17663
rect 5092 17660 5120 17768
rect 8478 17756 8484 17808
rect 8536 17796 8542 17808
rect 8573 17799 8631 17805
rect 8573 17796 8585 17799
rect 8536 17768 8585 17796
rect 8536 17756 8542 17768
rect 8573 17765 8585 17768
rect 8619 17765 8631 17799
rect 8573 17759 8631 17765
rect 19518 17756 19524 17808
rect 19576 17796 19582 17808
rect 28074 17796 28080 17808
rect 19576 17768 28080 17796
rect 19576 17756 19582 17768
rect 28074 17756 28080 17768
rect 28132 17756 28138 17808
rect 15286 17728 15292 17740
rect 13004 17700 15292 17728
rect 13004 17672 13032 17700
rect 15286 17688 15292 17700
rect 15344 17728 15350 17740
rect 16393 17731 16451 17737
rect 16393 17728 16405 17731
rect 15344 17700 16405 17728
rect 15344 17688 15350 17700
rect 16393 17697 16405 17700
rect 16439 17697 16451 17731
rect 23382 17728 23388 17740
rect 16393 17691 16451 17697
rect 19628 17700 23388 17728
rect 2547 17632 5120 17660
rect 2547 17629 2559 17632
rect 2501 17623 2559 17629
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 7190 17660 7196 17672
rect 5224 17632 7196 17660
rect 5224 17620 5230 17632
rect 7190 17620 7196 17632
rect 7248 17660 7254 17672
rect 8202 17660 8208 17672
rect 7248 17632 8208 17660
rect 7248 17620 7254 17632
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 12986 17660 12992 17672
rect 10827 17632 12992 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 14642 17620 14648 17672
rect 14700 17620 14706 17672
rect 14734 17620 14740 17672
rect 14792 17620 14798 17672
rect 16408 17660 16436 17691
rect 17954 17660 17960 17672
rect 16408 17632 17960 17660
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 2777 17595 2835 17601
rect 2777 17592 2789 17595
rect 1780 17564 2789 17592
rect 1673 17555 1731 17561
rect 2777 17561 2789 17564
rect 2823 17561 2835 17595
rect 2777 17555 2835 17561
rect 4240 17595 4298 17601
rect 4240 17561 4252 17595
rect 4286 17592 4298 17595
rect 4982 17592 4988 17604
rect 4286 17564 4988 17592
rect 4286 17561 4298 17564
rect 4240 17555 4298 17561
rect 4982 17552 4988 17564
rect 5040 17552 5046 17604
rect 7460 17595 7518 17601
rect 7460 17561 7472 17595
rect 7506 17592 7518 17595
rect 8938 17592 8944 17604
rect 7506 17564 8944 17592
rect 7506 17561 7518 17564
rect 7460 17555 7518 17561
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 11048 17595 11106 17601
rect 11048 17561 11060 17595
rect 11094 17592 11106 17595
rect 11698 17592 11704 17604
rect 11094 17564 11704 17592
rect 11094 17561 11106 17564
rect 11048 17555 11106 17561
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 16660 17595 16718 17601
rect 16660 17561 16672 17595
rect 16706 17592 16718 17595
rect 16850 17592 16856 17604
rect 16706 17564 16856 17592
rect 16706 17561 16718 17564
rect 16660 17555 16718 17561
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 17218 17552 17224 17604
rect 17276 17592 17282 17604
rect 18248 17592 18276 17623
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19628 17669 19656 17700
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 30466 17688 30472 17740
rect 30524 17728 30530 17740
rect 31205 17731 31263 17737
rect 31205 17728 31217 17731
rect 30524 17700 31217 17728
rect 30524 17688 30530 17700
rect 31205 17697 31217 17700
rect 31251 17728 31263 17731
rect 31294 17728 31300 17740
rect 31251 17700 31300 17728
rect 31251 17697 31263 17700
rect 31205 17691 31263 17697
rect 31294 17688 31300 17700
rect 31352 17688 31358 17740
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 19392 17632 19625 17660
rect 19392 17620 19398 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 20070 17660 20076 17672
rect 19935 17632 20076 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 21818 17620 21824 17672
rect 21876 17620 21882 17672
rect 22002 17620 22008 17672
rect 22060 17620 22066 17672
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17660 22155 17663
rect 22186 17660 22192 17672
rect 22143 17632 22192 17660
rect 22143 17629 22155 17632
rect 22097 17623 22155 17629
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 27522 17620 27528 17672
rect 27580 17660 27586 17672
rect 30837 17663 30895 17669
rect 30837 17660 30849 17663
rect 27580 17632 30849 17660
rect 27580 17620 27586 17632
rect 30837 17629 30849 17632
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 30929 17663 30987 17669
rect 30929 17629 30941 17663
rect 30975 17660 30987 17663
rect 31726 17660 31754 17836
rect 35713 17833 35725 17836
rect 35759 17864 35771 17867
rect 37918 17864 37924 17876
rect 35759 17836 37924 17864
rect 35759 17833 35771 17836
rect 35713 17827 35771 17833
rect 37918 17824 37924 17836
rect 37976 17824 37982 17876
rect 40494 17824 40500 17876
rect 40552 17864 40558 17876
rect 40681 17867 40739 17873
rect 40681 17864 40693 17867
rect 40552 17836 40693 17864
rect 40552 17824 40558 17836
rect 40681 17833 40693 17836
rect 40727 17833 40739 17867
rect 40681 17827 40739 17833
rect 38010 17756 38016 17808
rect 38068 17796 38074 17808
rect 40586 17796 40592 17808
rect 38068 17768 40592 17796
rect 38068 17756 38074 17768
rect 40586 17756 40592 17768
rect 40644 17756 40650 17808
rect 36538 17728 36544 17740
rect 34808 17700 36544 17728
rect 30975 17632 31754 17660
rect 32861 17663 32919 17669
rect 30975 17629 30987 17632
rect 30929 17623 30987 17629
rect 32861 17629 32873 17663
rect 32907 17660 32919 17663
rect 34808 17660 34836 17700
rect 36538 17688 36544 17700
rect 36596 17688 36602 17740
rect 41598 17728 41604 17740
rect 40420 17700 41604 17728
rect 32907 17632 34836 17660
rect 34885 17663 34943 17669
rect 32907 17629 32919 17632
rect 32861 17623 32919 17629
rect 34885 17629 34897 17663
rect 34931 17660 34943 17663
rect 35526 17660 35532 17672
rect 34931 17632 35532 17660
rect 34931 17629 34943 17632
rect 34885 17623 34943 17629
rect 17276 17564 18276 17592
rect 19797 17595 19855 17601
rect 17276 17552 17282 17564
rect 19797 17561 19809 17595
rect 19843 17592 19855 17595
rect 19978 17592 19984 17604
rect 19843 17564 19984 17592
rect 19843 17561 19855 17564
rect 19797 17555 19855 17561
rect 19978 17552 19984 17564
rect 20036 17552 20042 17604
rect 26234 17552 26240 17604
rect 26292 17592 26298 17604
rect 30650 17592 30656 17604
rect 26292 17564 30656 17592
rect 26292 17552 26298 17564
rect 30650 17552 30656 17564
rect 30708 17552 30714 17604
rect 30852 17592 30880 17623
rect 35526 17620 35532 17632
rect 35584 17620 35590 17672
rect 35618 17620 35624 17672
rect 35676 17620 35682 17672
rect 35802 17620 35808 17672
rect 35860 17620 35866 17672
rect 36808 17663 36866 17669
rect 36808 17629 36820 17663
rect 36854 17660 36866 17663
rect 37274 17660 37280 17672
rect 36854 17632 37280 17660
rect 36854 17629 36866 17632
rect 36808 17623 36866 17629
rect 37274 17620 37280 17632
rect 37332 17620 37338 17672
rect 40034 17620 40040 17672
rect 40092 17620 40098 17672
rect 40185 17663 40243 17669
rect 40185 17629 40197 17663
rect 40231 17660 40243 17663
rect 40420 17660 40448 17700
rect 41598 17688 41604 17700
rect 41656 17688 41662 17740
rect 40586 17669 40592 17672
rect 40231 17632 40448 17660
rect 40543 17663 40592 17669
rect 40231 17629 40243 17632
rect 40185 17623 40243 17629
rect 40543 17629 40555 17663
rect 40589 17629 40592 17663
rect 40543 17623 40592 17629
rect 40586 17620 40592 17623
rect 40644 17620 40650 17672
rect 31110 17592 31116 17604
rect 30852 17564 31116 17592
rect 31110 17552 31116 17564
rect 31168 17552 31174 17604
rect 31297 17595 31355 17601
rect 31297 17561 31309 17595
rect 31343 17592 31355 17595
rect 32030 17592 32036 17604
rect 31343 17564 32036 17592
rect 31343 17561 31355 17564
rect 31297 17555 31355 17561
rect 32030 17552 32036 17564
rect 32088 17552 32094 17604
rect 33128 17595 33186 17601
rect 33128 17561 33140 17595
rect 33174 17592 33186 17595
rect 33870 17592 33876 17604
rect 33174 17564 33876 17592
rect 33174 17561 33186 17564
rect 33128 17555 33186 17561
rect 33870 17552 33876 17564
rect 33928 17552 33934 17604
rect 36354 17552 36360 17604
rect 36412 17592 36418 17604
rect 37366 17592 37372 17604
rect 36412 17564 37372 17592
rect 36412 17552 36418 17564
rect 37366 17552 37372 17564
rect 37424 17592 37430 17604
rect 40313 17595 40371 17601
rect 40313 17592 40325 17595
rect 37424 17564 40325 17592
rect 37424 17552 37430 17564
rect 40236 17536 40264 17564
rect 40313 17561 40325 17564
rect 40359 17561 40371 17595
rect 40313 17555 40371 17561
rect 40405 17595 40463 17601
rect 40405 17561 40417 17595
rect 40451 17592 40463 17595
rect 40451 17564 40540 17592
rect 40451 17561 40463 17564
rect 40405 17555 40463 17561
rect 40512 17536 40540 17564
rect 1949 17527 2007 17533
rect 1949 17493 1961 17527
rect 1995 17524 2007 17527
rect 2406 17524 2412 17536
rect 1995 17496 2412 17524
rect 1995 17493 2007 17496
rect 1949 17487 2007 17493
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 11974 17524 11980 17536
rect 11388 17496 11980 17524
rect 11388 17484 11394 17496
rect 11974 17484 11980 17496
rect 12032 17524 12038 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 12032 17496 12173 17524
rect 12032 17484 12038 17496
rect 12161 17493 12173 17496
rect 12207 17493 12219 17527
rect 12161 17487 12219 17493
rect 14274 17484 14280 17536
rect 14332 17484 14338 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 17460 17496 18429 17524
rect 17460 17484 17466 17496
rect 18417 17493 18429 17496
rect 18463 17524 18475 17527
rect 20254 17524 20260 17536
rect 18463 17496 20260 17524
rect 18463 17493 18475 17496
rect 18417 17487 18475 17493
rect 20254 17484 20260 17496
rect 20312 17524 20318 17536
rect 21910 17524 21916 17536
rect 20312 17496 21916 17524
rect 20312 17484 20318 17496
rect 21910 17484 21916 17496
rect 21968 17524 21974 17536
rect 23566 17524 23572 17536
rect 21968 17496 23572 17524
rect 21968 17484 21974 17496
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 34241 17527 34299 17533
rect 34241 17524 34253 17527
rect 25280 17496 34253 17524
rect 25280 17484 25286 17496
rect 34241 17493 34253 17496
rect 34287 17524 34299 17527
rect 34422 17524 34428 17536
rect 34287 17496 34428 17524
rect 34287 17493 34299 17496
rect 34241 17487 34299 17493
rect 34422 17484 34428 17496
rect 34480 17484 34486 17536
rect 34606 17484 34612 17536
rect 34664 17524 34670 17536
rect 35069 17527 35127 17533
rect 35069 17524 35081 17527
rect 34664 17496 35081 17524
rect 34664 17484 34670 17496
rect 35069 17493 35081 17496
rect 35115 17493 35127 17527
rect 35069 17487 35127 17493
rect 36078 17484 36084 17536
rect 36136 17524 36142 17536
rect 37182 17524 37188 17536
rect 36136 17496 37188 17524
rect 36136 17484 36142 17496
rect 37182 17484 37188 17496
rect 37240 17484 37246 17536
rect 37274 17484 37280 17536
rect 37332 17524 37338 17536
rect 37921 17527 37979 17533
rect 37921 17524 37933 17527
rect 37332 17496 37933 17524
rect 37332 17484 37338 17496
rect 37921 17493 37933 17496
rect 37967 17493 37979 17527
rect 37921 17487 37979 17493
rect 40218 17484 40224 17536
rect 40276 17484 40282 17536
rect 40494 17484 40500 17536
rect 40552 17484 40558 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 2317 17323 2375 17329
rect 2317 17289 2329 17323
rect 2363 17320 2375 17323
rect 3418 17320 3424 17332
rect 2363 17292 3424 17320
rect 2363 17289 2375 17292
rect 2317 17283 2375 17289
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 4522 17280 4528 17332
rect 4580 17320 4586 17332
rect 4706 17320 4712 17332
rect 4580 17292 4712 17320
rect 4580 17280 4586 17292
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 4982 17280 4988 17332
rect 5040 17280 5046 17332
rect 7282 17280 7288 17332
rect 7340 17280 7346 17332
rect 8938 17280 8944 17332
rect 8996 17280 9002 17332
rect 11698 17280 11704 17332
rect 11756 17280 11762 17332
rect 16945 17323 17003 17329
rect 11900 17292 14872 17320
rect 934 17212 940 17264
rect 992 17252 998 17264
rect 3237 17255 3295 17261
rect 3237 17252 3249 17255
rect 992 17224 3249 17252
rect 992 17212 998 17224
rect 3237 17221 3249 17224
rect 3283 17221 3295 17255
rect 5626 17252 5632 17264
rect 3237 17215 3295 17221
rect 4356 17224 5632 17252
rect 4356 17193 4384 17224
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 7300 17252 7328 17280
rect 8018 17252 8024 17264
rect 7300 17224 8024 17252
rect 8018 17212 8024 17224
rect 8076 17252 8082 17264
rect 8205 17255 8263 17261
rect 8205 17252 8217 17255
rect 8076 17224 8217 17252
rect 8076 17212 8082 17224
rect 8205 17221 8217 17224
rect 8251 17221 8263 17255
rect 8205 17215 8263 17221
rect 8478 17212 8484 17264
rect 8536 17252 8542 17264
rect 9309 17255 9367 17261
rect 9309 17252 9321 17255
rect 8536 17224 9321 17252
rect 8536 17212 8542 17224
rect 9309 17221 9321 17224
rect 9355 17221 9367 17255
rect 9309 17215 9367 17221
rect 4522 17193 4528 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 4489 17187 4528 17193
rect 4489 17153 4501 17187
rect 4489 17147 4528 17153
rect 4522 17144 4528 17147
rect 4580 17144 4586 17196
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4709 17187 4767 17193
rect 4709 17153 4721 17187
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 4847 17187 4905 17193
rect 4847 17153 4859 17187
rect 4893 17184 4905 17187
rect 4893 17156 6914 17184
rect 4893 17153 4905 17156
rect 4847 17147 4905 17153
rect 2409 17119 2467 17125
rect 2409 17085 2421 17119
rect 2455 17085 2467 17119
rect 2409 17079 2467 17085
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 2682 17116 2688 17128
rect 2639 17088 2688 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 2424 17048 2452 17079
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 3234 17048 3240 17060
rect 2424 17020 3240 17048
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 4632 17048 4660 17147
rect 4724 17116 4752 17147
rect 5350 17116 5356 17128
rect 4724 17088 5356 17116
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 5902 17048 5908 17060
rect 4632 17020 5908 17048
rect 5902 17008 5908 17020
rect 5960 17008 5966 17060
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16980 2007 16983
rect 2038 16980 2044 16992
rect 1995 16952 2044 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 2038 16940 2044 16952
rect 2096 16940 2102 16992
rect 2406 16940 2412 16992
rect 2464 16980 2470 16992
rect 2682 16980 2688 16992
rect 2464 16952 2688 16980
rect 2464 16940 2470 16952
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 3329 16983 3387 16989
rect 3329 16949 3341 16983
rect 3375 16980 3387 16983
rect 6638 16980 6644 16992
rect 3375 16952 6644 16980
rect 3375 16949 3387 16952
rect 3329 16943 3387 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 6730 16940 6736 16992
rect 6788 16980 6794 16992
rect 6886 16980 6914 17156
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7340 17156 7849 17184
rect 7340 17144 7346 17156
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17184 9459 17187
rect 9582 17184 9588 17196
rect 9447 17156 9588 17184
rect 9447 17153 9459 17156
rect 9401 17147 9459 17153
rect 9140 17116 9168 17147
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 11900 17193 11928 17292
rect 11974 17212 11980 17264
rect 12032 17252 12038 17264
rect 12069 17255 12127 17261
rect 12069 17252 12081 17255
rect 12032 17224 12081 17252
rect 12032 17212 12038 17224
rect 12069 17221 12081 17224
rect 12115 17221 12127 17255
rect 12069 17215 12127 17221
rect 13256 17255 13314 17261
rect 13256 17221 13268 17255
rect 13302 17252 13314 17255
rect 14274 17252 14280 17264
rect 13302 17224 14280 17252
rect 13302 17221 13314 17224
rect 13256 17215 13314 17221
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 14844 17252 14872 17292
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 17034 17320 17040 17332
rect 16991 17292 17040 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 17310 17280 17316 17332
rect 17368 17320 17374 17332
rect 18506 17320 18512 17332
rect 17368 17292 18512 17320
rect 17368 17280 17374 17292
rect 18506 17280 18512 17292
rect 18564 17320 18570 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 18564 17292 19349 17320
rect 18564 17280 18570 17292
rect 19337 17289 19349 17292
rect 19383 17289 19395 17323
rect 19337 17283 19395 17289
rect 23569 17323 23627 17329
rect 23569 17289 23581 17323
rect 23615 17289 23627 17323
rect 33686 17320 33692 17332
rect 23569 17283 23627 17289
rect 23860 17292 33692 17320
rect 23584 17252 23612 17283
rect 14844 17224 23612 17252
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 12161 17187 12219 17193
rect 12161 17184 12173 17187
rect 11885 17147 11943 17153
rect 12084 17156 12173 17184
rect 11606 17116 11612 17128
rect 9140 17088 11612 17116
rect 11606 17076 11612 17088
rect 11664 17076 11670 17128
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 10318 17048 10324 17060
rect 9732 17020 10324 17048
rect 9732 17008 9738 17020
rect 10318 17008 10324 17020
rect 10376 17048 10382 17060
rect 12084 17048 12112 17156
rect 12161 17153 12173 17156
rect 12207 17184 12219 17187
rect 14734 17184 14740 17196
rect 12207 17156 14740 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15896 17156 15945 17184
rect 15896 17144 15902 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16390 17144 16396 17196
rect 16448 17184 16454 17196
rect 17313 17187 17371 17193
rect 17313 17184 17325 17187
rect 16448 17156 17325 17184
rect 16448 17144 16454 17156
rect 17313 17153 17325 17156
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17402 17144 17408 17196
rect 17460 17144 17466 17196
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 17954 17184 17960 17196
rect 17552 17156 17960 17184
rect 17552 17144 17558 17156
rect 17954 17144 17960 17156
rect 18012 17144 18018 17196
rect 18230 17193 18236 17196
rect 18224 17147 18236 17193
rect 18230 17144 18236 17147
rect 18288 17144 18294 17196
rect 23566 17144 23572 17196
rect 23624 17184 23630 17196
rect 23860 17193 23888 17292
rect 33686 17280 33692 17292
rect 33744 17280 33750 17332
rect 33870 17280 33876 17332
rect 33928 17280 33934 17332
rect 34146 17280 34152 17332
rect 34204 17320 34210 17332
rect 36725 17323 36783 17329
rect 36725 17320 36737 17323
rect 34204 17292 36737 17320
rect 34204 17280 34210 17292
rect 36725 17289 36737 17292
rect 36771 17289 36783 17323
rect 36725 17283 36783 17289
rect 37458 17280 37464 17332
rect 37516 17280 37522 17332
rect 43530 17280 43536 17332
rect 43588 17280 43594 17332
rect 45738 17280 45744 17332
rect 45796 17280 45802 17332
rect 45833 17323 45891 17329
rect 45833 17289 45845 17323
rect 45879 17320 45891 17323
rect 45922 17320 45928 17332
rect 45879 17292 45928 17320
rect 45879 17289 45891 17292
rect 45833 17283 45891 17289
rect 45922 17280 45928 17292
rect 45980 17320 45986 17332
rect 46382 17320 46388 17332
rect 45980 17292 46388 17320
rect 45980 17280 45986 17292
rect 46382 17280 46388 17292
rect 46440 17320 46446 17332
rect 46440 17292 46980 17320
rect 46440 17280 46446 17292
rect 23934 17212 23940 17264
rect 23992 17252 23998 17264
rect 30374 17252 30380 17264
rect 23992 17224 30380 17252
rect 23992 17212 23998 17224
rect 23753 17187 23811 17193
rect 23753 17184 23765 17187
rect 23624 17156 23765 17184
rect 23624 17144 23630 17156
rect 23753 17153 23765 17156
rect 23799 17153 23811 17187
rect 23753 17147 23811 17153
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17153 23903 17187
rect 23845 17147 23903 17153
rect 24118 17144 24124 17196
rect 24176 17184 24182 17196
rect 27172 17193 27200 17224
rect 30374 17212 30380 17224
rect 30432 17212 30438 17264
rect 34422 17212 34428 17264
rect 34480 17212 34486 17264
rect 34517 17255 34575 17261
rect 34517 17221 34529 17255
rect 34563 17252 34575 17255
rect 34790 17252 34796 17264
rect 34563 17224 34796 17252
rect 34563 17221 34575 17224
rect 34517 17215 34575 17221
rect 34790 17212 34796 17224
rect 34848 17212 34854 17264
rect 35986 17252 35992 17264
rect 34900 17224 35992 17252
rect 27430 17193 27436 17196
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 24176 17156 25053 17184
rect 24176 17144 24182 17156
rect 25041 17153 25053 17156
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27424 17147 27436 17193
rect 27430 17144 27436 17147
rect 27488 17144 27494 17196
rect 29178 17144 29184 17196
rect 29236 17184 29242 17196
rect 29273 17187 29331 17193
rect 29273 17184 29285 17187
rect 29236 17156 29285 17184
rect 29236 17144 29242 17156
rect 29273 17153 29285 17156
rect 29319 17153 29331 17187
rect 29273 17147 29331 17153
rect 29454 17144 29460 17196
rect 29512 17184 29518 17196
rect 30282 17184 30288 17196
rect 29512 17156 30288 17184
rect 29512 17144 29518 17156
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 32306 17144 32312 17196
rect 32364 17144 32370 17196
rect 32674 17144 32680 17196
rect 32732 17184 32738 17196
rect 32861 17187 32919 17193
rect 32861 17184 32873 17187
rect 32732 17156 32873 17184
rect 32732 17144 32738 17156
rect 32861 17153 32873 17156
rect 32907 17153 32919 17187
rect 32861 17147 32919 17153
rect 33244 17156 33456 17184
rect 12986 17076 12992 17128
rect 13044 17076 13050 17128
rect 17126 17076 17132 17128
rect 17184 17076 17190 17128
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 23937 17119 23995 17125
rect 23937 17085 23949 17119
rect 23983 17085 23995 17119
rect 23937 17079 23995 17085
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24210 17116 24216 17128
rect 24075 17088 24216 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 10376 17020 12112 17048
rect 14369 17051 14427 17057
rect 10376 17008 10382 17020
rect 14369 17017 14381 17051
rect 14415 17048 14427 17051
rect 14642 17048 14648 17060
rect 14415 17020 14648 17048
rect 14415 17017 14427 17020
rect 14369 17011 14427 17017
rect 14642 17008 14648 17020
rect 14700 17008 14706 17060
rect 17236 17048 17264 17079
rect 17862 17048 17868 17060
rect 17236 17020 17868 17048
rect 17862 17008 17868 17020
rect 17920 17008 17926 17060
rect 23658 17008 23664 17060
rect 23716 17048 23722 17060
rect 23952 17048 23980 17079
rect 24210 17076 24216 17088
rect 24268 17116 24274 17128
rect 24578 17116 24584 17128
rect 24268 17088 24584 17116
rect 24268 17076 24274 17088
rect 24578 17076 24584 17088
rect 24636 17076 24642 17128
rect 24670 17076 24676 17128
rect 24728 17116 24734 17128
rect 24765 17119 24823 17125
rect 24765 17116 24777 17119
rect 24728 17088 24777 17116
rect 24728 17076 24734 17088
rect 24765 17085 24777 17088
rect 24811 17085 24823 17119
rect 24765 17079 24823 17085
rect 24854 17076 24860 17128
rect 24912 17076 24918 17128
rect 24949 17119 25007 17125
rect 24949 17085 24961 17119
rect 24995 17085 25007 17119
rect 24949 17079 25007 17085
rect 23716 17020 23980 17048
rect 23716 17008 23722 17020
rect 9582 16980 9588 16992
rect 6788 16952 9588 16980
rect 6788 16940 6794 16952
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 16574 16980 16580 16992
rect 16255 16952 16580 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 16574 16940 16580 16952
rect 16632 16980 16638 16992
rect 18966 16980 18972 16992
rect 16632 16952 18972 16980
rect 16632 16940 16638 16952
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 23474 16940 23480 16992
rect 23532 16980 23538 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 23532 16952 24593 16980
rect 23532 16940 23538 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24964 16980 24992 17079
rect 28166 17076 28172 17128
rect 28224 17116 28230 17128
rect 30466 17116 30472 17128
rect 28224 17088 30472 17116
rect 28224 17076 28230 17088
rect 30466 17076 30472 17088
rect 30524 17076 30530 17128
rect 30650 17076 30656 17128
rect 30708 17116 30714 17128
rect 33244 17116 33272 17156
rect 30708 17088 33272 17116
rect 33321 17119 33379 17125
rect 30708 17076 30714 17088
rect 33321 17085 33333 17119
rect 33367 17085 33379 17119
rect 33321 17079 33379 17085
rect 32582 17008 32588 17060
rect 32640 17008 32646 17060
rect 33336 16992 33364 17079
rect 33428 17048 33456 17156
rect 33502 17144 33508 17196
rect 33560 17184 33566 17196
rect 34057 17187 34115 17193
rect 34057 17184 34069 17187
rect 33560 17156 34069 17184
rect 33560 17144 33566 17156
rect 34057 17153 34069 17156
rect 34103 17153 34115 17187
rect 34057 17147 34115 17153
rect 34149 17187 34207 17193
rect 34149 17153 34161 17187
rect 34195 17184 34207 17187
rect 34900 17184 34928 17224
rect 35986 17212 35992 17224
rect 36044 17212 36050 17264
rect 37274 17252 37280 17264
rect 36280 17224 37280 17252
rect 34195 17156 34928 17184
rect 34977 17187 35035 17193
rect 34195 17153 34207 17156
rect 34149 17147 34207 17153
rect 34977 17153 34989 17187
rect 35023 17184 35035 17187
rect 35894 17184 35900 17196
rect 35023 17156 35900 17184
rect 35023 17153 35035 17156
rect 34977 17147 35035 17153
rect 35894 17144 35900 17156
rect 35952 17144 35958 17196
rect 36078 17144 36084 17196
rect 36136 17144 36142 17196
rect 36280 17193 36308 17224
rect 37274 17212 37280 17224
rect 37332 17212 37338 17264
rect 38010 17252 38016 17264
rect 37476 17224 38016 17252
rect 36229 17187 36308 17193
rect 36229 17153 36241 17187
rect 36275 17156 36308 17187
rect 36275 17153 36287 17156
rect 36229 17147 36287 17153
rect 36354 17144 36360 17196
rect 36412 17144 36418 17196
rect 36630 17193 36636 17196
rect 36449 17187 36507 17193
rect 36449 17153 36461 17187
rect 36495 17153 36507 17187
rect 36449 17147 36507 17153
rect 36587 17187 36636 17193
rect 36587 17153 36599 17187
rect 36633 17153 36636 17187
rect 36587 17147 36636 17153
rect 35253 17119 35311 17125
rect 35253 17085 35265 17119
rect 35299 17116 35311 17119
rect 35526 17116 35532 17128
rect 35299 17088 35532 17116
rect 35299 17085 35311 17088
rect 35253 17079 35311 17085
rect 35526 17076 35532 17088
rect 35584 17076 35590 17128
rect 36464 17116 36492 17147
rect 36630 17144 36636 17147
rect 36688 17184 36694 17196
rect 37476 17184 37504 17224
rect 38010 17212 38016 17224
rect 38068 17212 38074 17264
rect 40218 17212 40224 17264
rect 40276 17252 40282 17264
rect 43548 17252 43576 17280
rect 43898 17252 43904 17264
rect 40276 17224 43904 17252
rect 40276 17212 40282 17224
rect 43898 17212 43904 17224
rect 43956 17252 43962 17264
rect 43993 17255 44051 17261
rect 43993 17252 44005 17255
rect 43956 17224 44005 17252
rect 43956 17212 43962 17224
rect 43993 17221 44005 17224
rect 44039 17221 44051 17255
rect 43993 17215 44051 17221
rect 44085 17255 44143 17261
rect 44085 17221 44097 17255
rect 44131 17252 44143 17255
rect 44450 17252 44456 17264
rect 44131 17224 44456 17252
rect 44131 17221 44143 17224
rect 44085 17215 44143 17221
rect 44450 17212 44456 17224
rect 44508 17212 44514 17264
rect 45664 17224 46704 17252
rect 45664 17196 45692 17224
rect 36688 17156 37504 17184
rect 36688 17144 36694 17156
rect 37550 17144 37556 17196
rect 37608 17184 37614 17196
rect 37645 17187 37703 17193
rect 37645 17184 37657 17187
rect 37608 17156 37657 17184
rect 37608 17144 37614 17156
rect 37645 17153 37657 17156
rect 37691 17153 37703 17187
rect 37645 17147 37703 17153
rect 37918 17144 37924 17196
rect 37976 17144 37982 17196
rect 43530 17144 43536 17196
rect 43588 17184 43594 17196
rect 43717 17187 43775 17193
rect 43717 17184 43729 17187
rect 43588 17156 43729 17184
rect 43588 17144 43594 17156
rect 43717 17153 43729 17156
rect 43763 17153 43775 17187
rect 43717 17147 43775 17153
rect 43806 17144 43812 17196
rect 43864 17184 43870 17196
rect 44174 17184 44180 17196
rect 44232 17193 44238 17196
rect 43864 17156 43909 17184
rect 44140 17156 44180 17184
rect 43864 17144 43870 17156
rect 44174 17144 44180 17156
rect 44232 17147 44240 17193
rect 44232 17144 44238 17147
rect 45646 17144 45652 17196
rect 45704 17144 45710 17196
rect 46676 17193 46704 17224
rect 46952 17193 46980 17292
rect 46661 17187 46719 17193
rect 46661 17153 46673 17187
rect 46707 17153 46719 17187
rect 46661 17147 46719 17153
rect 46845 17187 46903 17193
rect 46845 17153 46857 17187
rect 46891 17153 46903 17187
rect 46845 17147 46903 17153
rect 46937 17187 46995 17193
rect 46937 17153 46949 17187
rect 46983 17153 46995 17187
rect 46937 17147 46995 17153
rect 36906 17116 36912 17128
rect 36464 17088 36912 17116
rect 36906 17076 36912 17088
rect 36964 17076 36970 17128
rect 37737 17119 37795 17125
rect 37737 17085 37749 17119
rect 37783 17116 37795 17119
rect 38654 17116 38660 17128
rect 37783 17088 38660 17116
rect 37783 17085 37795 17088
rect 37737 17079 37795 17085
rect 38654 17076 38660 17088
rect 38712 17076 38718 17128
rect 45738 17076 45744 17128
rect 45796 17116 45802 17128
rect 46106 17116 46112 17128
rect 45796 17088 46112 17116
rect 45796 17076 45802 17088
rect 46106 17076 46112 17088
rect 46164 17116 46170 17128
rect 46860 17116 46888 17147
rect 46164 17088 46888 17116
rect 46164 17076 46170 17088
rect 33428 17020 36492 17048
rect 27890 16980 27896 16992
rect 24964 16952 27896 16980
rect 24581 16943 24639 16949
rect 27890 16940 27896 16952
rect 27948 16980 27954 16992
rect 28537 16983 28595 16989
rect 28537 16980 28549 16983
rect 27948 16952 28549 16980
rect 27948 16940 27954 16952
rect 28537 16949 28549 16952
rect 28583 16949 28595 16983
rect 28537 16943 28595 16949
rect 28902 16940 28908 16992
rect 28960 16980 28966 16992
rect 29365 16983 29423 16989
rect 29365 16980 29377 16983
rect 28960 16952 29377 16980
rect 28960 16940 28966 16952
rect 29365 16949 29377 16952
rect 29411 16949 29423 16983
rect 29365 16943 29423 16949
rect 33318 16940 33324 16992
rect 33376 16980 33382 16992
rect 35618 16980 35624 16992
rect 33376 16952 35624 16980
rect 33376 16940 33382 16952
rect 35618 16940 35624 16952
rect 35676 16940 35682 16992
rect 35894 16940 35900 16992
rect 35952 16980 35958 16992
rect 36354 16980 36360 16992
rect 35952 16952 36360 16980
rect 35952 16940 35958 16952
rect 36354 16940 36360 16952
rect 36412 16940 36418 16992
rect 36464 16980 36492 17020
rect 36538 17008 36544 17060
rect 36596 17048 36602 17060
rect 37182 17048 37188 17060
rect 36596 17020 37188 17048
rect 36596 17008 36602 17020
rect 37182 17008 37188 17020
rect 37240 17008 37246 17060
rect 37826 17008 37832 17060
rect 37884 17008 37890 17060
rect 45462 17008 45468 17060
rect 45520 17008 45526 17060
rect 45830 17008 45836 17060
rect 45888 17048 45894 17060
rect 46477 17051 46535 17057
rect 46477 17048 46489 17051
rect 45888 17020 46489 17048
rect 45888 17008 45894 17020
rect 46477 17017 46489 17020
rect 46523 17017 46535 17051
rect 46477 17011 46535 17017
rect 44361 16983 44419 16989
rect 44361 16980 44373 16983
rect 36464 16952 44373 16980
rect 44361 16949 44373 16952
rect 44407 16949 44419 16983
rect 44361 16943 44419 16949
rect 45278 16940 45284 16992
rect 45336 16980 45342 16992
rect 46017 16983 46075 16989
rect 46017 16980 46029 16983
rect 45336 16952 46029 16980
rect 45336 16940 45342 16952
rect 46017 16949 46029 16952
rect 46063 16949 46075 16983
rect 46017 16943 46075 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 6273 16779 6331 16785
rect 6273 16745 6285 16779
rect 6319 16776 6331 16779
rect 7006 16776 7012 16788
rect 6319 16748 7012 16776
rect 6319 16745 6331 16748
rect 6273 16739 6331 16745
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 9401 16779 9459 16785
rect 9401 16745 9413 16779
rect 9447 16776 9459 16779
rect 10502 16776 10508 16788
rect 9447 16748 10508 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 23293 16779 23351 16785
rect 23293 16776 23305 16779
rect 14516 16748 23305 16776
rect 14516 16736 14522 16748
rect 23293 16745 23305 16748
rect 23339 16745 23351 16779
rect 23293 16739 23351 16745
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 24762 16776 24768 16788
rect 24084 16748 24768 16776
rect 24084 16736 24090 16748
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 24946 16736 24952 16788
rect 25004 16776 25010 16788
rect 27341 16779 27399 16785
rect 25004 16748 27200 16776
rect 25004 16736 25010 16748
rect 4249 16711 4307 16717
rect 4249 16677 4261 16711
rect 4295 16708 4307 16711
rect 6178 16708 6184 16720
rect 4295 16680 6184 16708
rect 4295 16677 4307 16680
rect 4249 16671 4307 16677
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 20714 16708 20720 16720
rect 16684 16680 20720 16708
rect 1762 16600 1768 16652
rect 1820 16600 1826 16652
rect 2038 16600 2044 16652
rect 2096 16600 2102 16652
rect 5166 16600 5172 16652
rect 5224 16640 5230 16652
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 5224 16612 6745 16640
rect 5224 16600 5230 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 6733 16603 6791 16609
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16640 10195 16643
rect 14829 16643 14887 16649
rect 10183 16612 14596 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 14568 16584 14596 16612
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 15194 16640 15200 16652
rect 14875 16612 15200 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 16684 16649 16712 16680
rect 20714 16668 20720 16680
rect 20772 16668 20778 16720
rect 21358 16668 21364 16720
rect 21416 16708 21422 16720
rect 27172 16708 27200 16748
rect 27341 16745 27353 16779
rect 27387 16776 27399 16779
rect 27430 16776 27436 16788
rect 27387 16748 27436 16776
rect 27387 16745 27399 16748
rect 27341 16739 27399 16745
rect 27430 16736 27436 16748
rect 27488 16736 27494 16788
rect 28902 16736 28908 16788
rect 28960 16736 28966 16788
rect 30374 16776 30380 16788
rect 29748 16748 30380 16776
rect 28166 16708 28172 16720
rect 21416 16680 25452 16708
rect 27172 16680 28172 16708
rect 21416 16668 21422 16680
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 15436 16612 16681 16640
rect 15436 16600 15442 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16609 16911 16643
rect 17034 16640 17040 16652
rect 16853 16606 16911 16609
rect 16960 16612 17040 16640
rect 16960 16606 16988 16612
rect 16853 16603 16988 16606
rect 934 16532 940 16584
rect 992 16572 998 16584
rect 992 16544 2728 16572
rect 992 16532 998 16544
rect 2700 16504 2728 16544
rect 3418 16532 3424 16584
rect 3476 16532 3482 16584
rect 5626 16532 5632 16584
rect 5684 16532 5690 16584
rect 5810 16581 5816 16584
rect 5777 16575 5816 16581
rect 5777 16541 5789 16575
rect 5777 16535 5816 16541
rect 5810 16532 5816 16535
rect 5868 16532 5874 16584
rect 5902 16532 5908 16584
rect 5960 16532 5966 16584
rect 5994 16532 6000 16584
rect 6052 16532 6058 16584
rect 6135 16575 6193 16581
rect 6135 16541 6147 16575
rect 6181 16572 6193 16575
rect 6638 16572 6644 16584
rect 6181 16544 6644 16572
rect 6181 16541 6193 16544
rect 6135 16535 6193 16541
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 7006 16581 7012 16584
rect 7000 16535 7012 16581
rect 7006 16532 7012 16535
rect 7064 16532 7070 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 9766 16572 9772 16584
rect 9723 16544 9772 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 9766 16532 9772 16544
rect 9824 16572 9830 16584
rect 11790 16572 11796 16584
rect 9824 16544 11796 16572
rect 9824 16532 9830 16544
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 15013 16575 15071 16581
rect 15013 16572 15025 16575
rect 14608 16544 15025 16572
rect 14608 16532 14614 16544
rect 15013 16541 15025 16544
rect 15059 16541 15071 16575
rect 15013 16535 15071 16541
rect 15286 16532 15292 16584
rect 15344 16532 15350 16584
rect 16574 16572 16580 16584
rect 16536 16544 16580 16572
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 16761 16575 16819 16581
rect 16868 16578 16988 16603
rect 17034 16600 17040 16612
rect 17092 16640 17098 16652
rect 17310 16640 17316 16652
rect 17092 16612 17316 16640
rect 17092 16600 17098 16612
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16640 18475 16643
rect 19426 16640 19432 16652
rect 18463 16612 19432 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 23474 16600 23480 16652
rect 23532 16600 23538 16652
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16640 23627 16643
rect 24946 16640 24952 16652
rect 23615 16612 24952 16640
rect 23615 16609 23627 16612
rect 23569 16603 23627 16609
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 25314 16600 25320 16652
rect 25372 16600 25378 16652
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 4065 16507 4123 16513
rect 4065 16504 4077 16507
rect 2700 16476 4077 16504
rect 4065 16473 4077 16476
rect 4111 16473 4123 16507
rect 4065 16467 4123 16473
rect 6012 16436 6040 16532
rect 6822 16464 6828 16516
rect 6880 16504 6886 16516
rect 9585 16507 9643 16513
rect 9585 16504 9597 16507
rect 6880 16476 9597 16504
rect 6880 16464 6886 16476
rect 9585 16473 9597 16476
rect 9631 16473 9643 16507
rect 16776 16504 16804 16535
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17736 16544 18061 16572
rect 17736 16532 17742 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 9585 16467 9643 16473
rect 16316 16476 16804 16504
rect 16316 16448 16344 16476
rect 17034 16464 17040 16516
rect 17092 16504 17098 16516
rect 17865 16507 17923 16513
rect 17865 16504 17877 16507
rect 17092 16476 17877 16504
rect 17092 16464 17098 16476
rect 17865 16473 17877 16476
rect 17911 16473 17923 16507
rect 18064 16504 18092 16535
rect 21174 16532 21180 16584
rect 21232 16572 21238 16584
rect 23658 16572 23664 16584
rect 21232 16544 23664 16572
rect 21232 16532 21238 16544
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 23753 16575 23811 16581
rect 23753 16541 23765 16575
rect 23799 16572 23811 16575
rect 24210 16572 24216 16584
rect 23799 16544 24216 16572
rect 23799 16541 23811 16544
rect 23753 16535 23811 16541
rect 20806 16504 20812 16516
rect 18064 16476 20812 16504
rect 17865 16467 17923 16473
rect 20806 16464 20812 16476
rect 20864 16504 20870 16516
rect 22186 16504 22192 16516
rect 20864 16476 22192 16504
rect 20864 16464 20870 16476
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 23290 16464 23296 16516
rect 23348 16504 23354 16516
rect 23768 16504 23796 16535
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 25038 16572 25044 16584
rect 24728 16544 25044 16572
rect 24728 16532 24734 16544
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16541 25191 16575
rect 25133 16535 25191 16541
rect 23348 16476 23796 16504
rect 23348 16464 23354 16476
rect 23842 16464 23848 16516
rect 23900 16504 23906 16516
rect 24688 16504 24716 16532
rect 23900 16476 24716 16504
rect 23900 16464 23906 16476
rect 24762 16464 24768 16516
rect 24820 16504 24826 16516
rect 25148 16504 25176 16535
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 24820 16476 25176 16504
rect 25424 16504 25452 16680
rect 28166 16668 28172 16680
rect 28224 16668 28230 16720
rect 27522 16600 27528 16652
rect 27580 16600 27586 16652
rect 28920 16640 28948 16736
rect 27632 16612 28948 16640
rect 27632 16581 27660 16612
rect 29086 16600 29092 16652
rect 29144 16600 29150 16652
rect 29748 16649 29776 16748
rect 30374 16736 30380 16748
rect 30432 16776 30438 16788
rect 31294 16776 31300 16788
rect 30432 16748 31300 16776
rect 30432 16736 30438 16748
rect 31294 16736 31300 16748
rect 31352 16736 31358 16788
rect 32582 16736 32588 16788
rect 32640 16776 32646 16788
rect 35894 16776 35900 16788
rect 32640 16748 35900 16776
rect 32640 16736 32646 16748
rect 35894 16736 35900 16748
rect 35952 16736 35958 16788
rect 36633 16779 36691 16785
rect 36633 16745 36645 16779
rect 36679 16776 36691 16779
rect 37826 16776 37832 16788
rect 36679 16748 37832 16776
rect 36679 16745 36691 16748
rect 36633 16739 36691 16745
rect 37826 16736 37832 16748
rect 37884 16736 37890 16788
rect 43533 16779 43591 16785
rect 43533 16745 43545 16779
rect 43579 16776 43591 16779
rect 43806 16776 43812 16788
rect 43579 16748 43812 16776
rect 43579 16745 43591 16748
rect 43533 16739 43591 16745
rect 43806 16736 43812 16748
rect 43864 16736 43870 16788
rect 34146 16668 34152 16720
rect 34204 16708 34210 16720
rect 36722 16708 36728 16720
rect 34204 16680 36728 16708
rect 34204 16668 34210 16680
rect 36722 16668 36728 16680
rect 36780 16668 36786 16720
rect 43714 16668 43720 16720
rect 43772 16708 43778 16720
rect 47949 16711 48007 16717
rect 47949 16708 47961 16711
rect 43772 16680 47961 16708
rect 43772 16668 43778 16680
rect 47949 16677 47961 16680
rect 47995 16677 48007 16711
rect 47949 16671 48007 16677
rect 29733 16643 29791 16649
rect 29733 16609 29745 16643
rect 29779 16609 29791 16643
rect 33318 16640 33324 16652
rect 29733 16603 29791 16609
rect 30760 16612 33324 16640
rect 27617 16575 27675 16581
rect 27617 16541 27629 16575
rect 27663 16541 27675 16575
rect 27617 16535 27675 16541
rect 27890 16532 27896 16584
rect 27948 16532 27954 16584
rect 28813 16575 28871 16581
rect 28813 16572 28825 16575
rect 28552 16544 28825 16572
rect 27985 16507 28043 16513
rect 27985 16504 27997 16507
rect 25424 16476 27997 16504
rect 24820 16464 24826 16476
rect 27985 16473 27997 16476
rect 28031 16473 28043 16507
rect 27985 16467 28043 16473
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 6012 16408 8125 16436
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 11514 16396 11520 16448
rect 11572 16436 11578 16448
rect 11698 16436 11704 16448
rect 11572 16408 11704 16436
rect 11572 16396 11578 16408
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 16298 16436 16304 16448
rect 15243 16408 16304 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16393 16439 16451 16445
rect 16393 16405 16405 16439
rect 16439 16436 16451 16439
rect 17126 16436 17132 16448
rect 16439 16408 17132 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 20070 16436 20076 16448
rect 17460 16408 20076 16436
rect 17460 16396 17466 16408
rect 20070 16396 20076 16408
rect 20128 16436 20134 16448
rect 21358 16436 21364 16448
rect 20128 16408 21364 16436
rect 20128 16396 20134 16408
rect 21358 16396 21364 16408
rect 21416 16396 21422 16448
rect 23566 16396 23572 16448
rect 23624 16436 23630 16448
rect 24857 16439 24915 16445
rect 24857 16436 24869 16439
rect 23624 16408 24869 16436
rect 23624 16396 23630 16408
rect 24857 16405 24869 16408
rect 24903 16405 24915 16439
rect 24857 16399 24915 16405
rect 27522 16396 27528 16448
rect 27580 16436 27586 16448
rect 28552 16436 28580 16544
rect 28813 16541 28825 16544
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 29178 16532 29184 16584
rect 29236 16572 29242 16584
rect 30760 16572 30788 16612
rect 33318 16600 33324 16612
rect 33376 16600 33382 16652
rect 37274 16640 37280 16652
rect 36832 16612 37280 16640
rect 29236 16544 30788 16572
rect 29236 16532 29242 16544
rect 34606 16532 34612 16584
rect 34664 16572 34670 16584
rect 36832 16581 36860 16612
rect 37274 16600 37280 16612
rect 37332 16600 37338 16652
rect 38013 16643 38071 16649
rect 38013 16609 38025 16643
rect 38059 16640 38071 16643
rect 38654 16640 38660 16652
rect 38059 16612 38660 16640
rect 38059 16609 38071 16612
rect 38013 16603 38071 16609
rect 38654 16600 38660 16612
rect 38712 16600 38718 16652
rect 40310 16600 40316 16652
rect 40368 16600 40374 16652
rect 42153 16643 42211 16649
rect 42153 16640 42165 16643
rect 41386 16612 42165 16640
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34664 16544 34897 16572
rect 34664 16532 34670 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 35069 16575 35127 16581
rect 35069 16541 35081 16575
rect 35115 16541 35127 16575
rect 35069 16535 35127 16541
rect 36633 16575 36691 16581
rect 36633 16541 36645 16575
rect 36679 16541 36691 16575
rect 36633 16535 36691 16541
rect 36817 16575 36875 16581
rect 36817 16541 36829 16575
rect 36863 16541 36875 16575
rect 40328 16572 40356 16600
rect 41386 16572 41414 16612
rect 42153 16609 42165 16612
rect 42199 16609 42211 16643
rect 42153 16603 42211 16609
rect 45738 16600 45744 16652
rect 45796 16640 45802 16652
rect 46293 16643 46351 16649
rect 46293 16640 46305 16643
rect 45796 16612 46305 16640
rect 45796 16600 45802 16612
rect 46293 16609 46305 16612
rect 46339 16640 46351 16643
rect 47489 16643 47547 16649
rect 47489 16640 47501 16643
rect 46339 16612 47501 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47489 16609 47501 16612
rect 47535 16609 47547 16643
rect 47489 16603 47547 16609
rect 40328 16544 41414 16572
rect 36817 16535 36875 16541
rect 29089 16507 29147 16513
rect 29089 16473 29101 16507
rect 29135 16504 29147 16507
rect 29978 16507 30036 16513
rect 29978 16504 29990 16507
rect 29135 16476 29990 16504
rect 29135 16473 29147 16476
rect 29089 16467 29147 16473
rect 29978 16473 29990 16476
rect 30024 16473 30036 16507
rect 29978 16467 30036 16473
rect 34514 16464 34520 16516
rect 34572 16504 34578 16516
rect 35084 16504 35112 16535
rect 34572 16476 35112 16504
rect 34572 16464 34578 16476
rect 27580 16408 28580 16436
rect 27580 16396 27586 16408
rect 30742 16396 30748 16448
rect 30800 16436 30806 16448
rect 31113 16439 31171 16445
rect 31113 16436 31125 16439
rect 30800 16408 31125 16436
rect 30800 16396 30806 16408
rect 31113 16405 31125 16408
rect 31159 16405 31171 16439
rect 31113 16399 31171 16405
rect 34790 16396 34796 16448
rect 34848 16436 34854 16448
rect 34977 16439 35035 16445
rect 34977 16436 34989 16439
rect 34848 16408 34989 16436
rect 34848 16396 34854 16408
rect 34977 16405 34989 16408
rect 35023 16405 35035 16439
rect 36648 16436 36676 16535
rect 43806 16532 43812 16584
rect 43864 16572 43870 16584
rect 45646 16572 45652 16584
rect 43864 16544 45652 16572
rect 43864 16532 43870 16544
rect 45646 16532 45652 16544
rect 45704 16572 45710 16584
rect 45925 16575 45983 16581
rect 45925 16572 45937 16575
rect 45704 16544 45937 16572
rect 45704 16532 45710 16544
rect 45925 16541 45937 16544
rect 45971 16541 45983 16575
rect 45925 16535 45983 16541
rect 46106 16532 46112 16584
rect 46164 16532 46170 16584
rect 46382 16532 46388 16584
rect 46440 16532 46446 16584
rect 47581 16575 47639 16581
rect 47581 16572 47593 16575
rect 47504 16544 47593 16572
rect 36722 16464 36728 16516
rect 36780 16504 36786 16516
rect 37553 16507 37611 16513
rect 37553 16504 37565 16507
rect 36780 16476 37565 16504
rect 36780 16464 36786 16476
rect 37553 16473 37565 16476
rect 37599 16473 37611 16507
rect 37553 16467 37611 16473
rect 37642 16464 37648 16516
rect 37700 16464 37706 16516
rect 40034 16464 40040 16516
rect 40092 16504 40098 16516
rect 40558 16507 40616 16513
rect 40558 16504 40570 16507
rect 40092 16476 40570 16504
rect 40092 16464 40098 16476
rect 40558 16473 40570 16476
rect 40604 16473 40616 16507
rect 40558 16467 40616 16473
rect 42420 16507 42478 16513
rect 42420 16473 42432 16507
rect 42466 16504 42478 16507
rect 45554 16504 45560 16516
rect 42466 16476 45560 16504
rect 42466 16473 42478 16476
rect 42420 16467 42478 16473
rect 45554 16464 45560 16476
rect 45612 16464 45618 16516
rect 37274 16436 37280 16448
rect 36648 16408 37280 16436
rect 34977 16399 35035 16405
rect 37274 16396 37280 16408
rect 37332 16396 37338 16448
rect 37458 16396 37464 16448
rect 37516 16436 37522 16448
rect 38838 16436 38844 16448
rect 37516 16408 38844 16436
rect 37516 16396 37522 16408
rect 38838 16396 38844 16408
rect 38896 16396 38902 16448
rect 41693 16439 41751 16445
rect 41693 16405 41705 16439
rect 41739 16436 41751 16439
rect 43622 16436 43628 16448
rect 41739 16408 43628 16436
rect 41739 16405 41751 16408
rect 41693 16399 41751 16405
rect 43622 16396 43628 16408
rect 43680 16436 43686 16448
rect 45462 16436 45468 16448
rect 43680 16408 45468 16436
rect 43680 16396 43686 16408
rect 45462 16396 45468 16408
rect 45520 16436 45526 16448
rect 47504 16436 47532 16544
rect 47581 16541 47593 16544
rect 47627 16541 47639 16575
rect 47581 16535 47639 16541
rect 45520 16408 47532 16436
rect 45520 16396 45526 16408
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 2832 16204 3433 16232
rect 2832 16192 2838 16204
rect 3421 16201 3433 16204
rect 3467 16201 3479 16235
rect 3421 16195 3479 16201
rect 5810 16192 5816 16244
rect 5868 16232 5874 16244
rect 5868 16204 11744 16232
rect 5868 16192 5874 16204
rect 934 16124 940 16176
rect 992 16164 998 16176
rect 1857 16167 1915 16173
rect 1857 16164 1869 16167
rect 992 16136 1869 16164
rect 992 16124 998 16136
rect 1857 16133 1869 16136
rect 1903 16133 1915 16167
rect 11514 16164 11520 16176
rect 1857 16127 1915 16133
rect 3252 16136 11520 16164
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 3252 16096 3280 16136
rect 11514 16124 11520 16136
rect 11572 16124 11578 16176
rect 1627 16068 3280 16096
rect 3329 16099 3387 16105
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 4062 16096 4068 16108
rect 3375 16068 4068 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7248 16068 7665 16096
rect 7248 16056 7254 16068
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 7909 16099 7967 16105
rect 7909 16096 7921 16099
rect 7800 16068 7921 16096
rect 7800 16056 7806 16068
rect 7909 16065 7921 16068
rect 7955 16065 7967 16099
rect 7909 16059 7967 16065
rect 2590 15988 2596 16040
rect 2648 16028 2654 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 2648 16000 3617 16028
rect 2648 15988 2654 16000
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 3620 15960 3648 15991
rect 6730 15988 6736 16040
rect 6788 15988 6794 16040
rect 3620 15932 6914 15960
rect 2958 15852 2964 15904
rect 3016 15852 3022 15904
rect 6886 15892 6914 15932
rect 8018 15892 8024 15904
rect 6886 15864 8024 15892
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 9033 15895 9091 15901
rect 9033 15861 9045 15895
rect 9079 15892 9091 15895
rect 9306 15892 9312 15904
rect 9079 15864 9312 15892
rect 9079 15861 9091 15864
rect 9033 15855 9091 15861
rect 9306 15852 9312 15864
rect 9364 15852 9370 15904
rect 11716 15892 11744 16204
rect 14182 16192 14188 16244
rect 14240 16232 14246 16244
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 14240 16204 14381 16232
rect 14240 16192 14246 16204
rect 14369 16201 14381 16204
rect 14415 16232 14427 16235
rect 14642 16232 14648 16244
rect 14415 16204 14648 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 16298 16192 16304 16244
rect 16356 16192 16362 16244
rect 18141 16235 18199 16241
rect 18141 16201 18153 16235
rect 18187 16232 18199 16235
rect 18230 16232 18236 16244
rect 18187 16204 18236 16232
rect 18187 16201 18199 16204
rect 18141 16195 18199 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18506 16192 18512 16244
rect 18564 16192 18570 16244
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 31018 16232 31024 16244
rect 25188 16204 31024 16232
rect 25188 16192 25194 16204
rect 31018 16192 31024 16204
rect 31076 16192 31082 16244
rect 33686 16192 33692 16244
rect 33744 16232 33750 16244
rect 34517 16235 34575 16241
rect 34517 16232 34529 16235
rect 33744 16204 34529 16232
rect 33744 16192 33750 16204
rect 34517 16201 34529 16204
rect 34563 16201 34575 16235
rect 34517 16195 34575 16201
rect 37274 16192 37280 16244
rect 37332 16232 37338 16244
rect 37829 16235 37887 16241
rect 37829 16232 37841 16235
rect 37332 16204 37841 16232
rect 37332 16192 37338 16204
rect 37829 16201 37841 16204
rect 37875 16201 37887 16235
rect 37829 16195 37887 16201
rect 40034 16192 40040 16244
rect 40092 16192 40098 16244
rect 40402 16192 40408 16244
rect 40460 16192 40466 16244
rect 44910 16232 44916 16244
rect 43916 16204 44916 16232
rect 12986 16124 12992 16176
rect 13044 16164 13050 16176
rect 15194 16173 15200 16176
rect 15188 16164 15200 16173
rect 13044 16136 14964 16164
rect 15155 16136 15200 16164
rect 13044 16124 13050 16136
rect 13256 16099 13314 16105
rect 13256 16065 13268 16099
rect 13302 16096 13314 16099
rect 14826 16096 14832 16108
rect 13302 16068 14832 16096
rect 13302 16065 13314 16068
rect 13256 16059 13314 16065
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 14936 16105 14964 16136
rect 15188 16127 15200 16136
rect 15194 16124 15200 16127
rect 15252 16124 15258 16176
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 17586 16164 17592 16176
rect 17083 16136 17592 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 17586 16124 17592 16136
rect 17644 16164 17650 16176
rect 18874 16164 18880 16176
rect 17644 16136 18880 16164
rect 17644 16124 17650 16136
rect 18874 16124 18880 16136
rect 18932 16124 18938 16176
rect 18966 16124 18972 16176
rect 19024 16164 19030 16176
rect 20990 16164 20996 16176
rect 19024 16136 20996 16164
rect 19024 16124 19030 16136
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15028 16068 15976 16096
rect 12986 15988 12992 16040
rect 13044 15988 13050 16040
rect 15028 16028 15056 16068
rect 14844 16000 15056 16028
rect 15948 16028 15976 16068
rect 16942 16056 16948 16108
rect 17000 16056 17006 16108
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16065 18383 16099
rect 18325 16059 18383 16065
rect 18046 16028 18052 16040
rect 15948 16000 18052 16028
rect 14844 15892 14872 16000
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18340 16028 18368 16059
rect 18598 16056 18604 16108
rect 18656 16056 18662 16108
rect 20640 16105 20668 16136
rect 20990 16124 20996 16136
rect 21048 16124 21054 16176
rect 25038 16124 25044 16176
rect 25096 16164 25102 16176
rect 25590 16164 25596 16176
rect 25096 16136 25596 16164
rect 25096 16124 25102 16136
rect 25590 16124 25596 16136
rect 25648 16164 25654 16176
rect 26053 16167 26111 16173
rect 26053 16164 26065 16167
rect 25648 16136 26065 16164
rect 25648 16124 25654 16136
rect 26053 16133 26065 16136
rect 26099 16133 26111 16167
rect 26053 16127 26111 16133
rect 29178 16124 29184 16176
rect 29236 16164 29242 16176
rect 29825 16167 29883 16173
rect 29825 16164 29837 16167
rect 29236 16136 29837 16164
rect 29236 16124 29242 16136
rect 29825 16133 29837 16136
rect 29871 16133 29883 16167
rect 29825 16127 29883 16133
rect 30466 16124 30472 16176
rect 30524 16164 30530 16176
rect 33778 16164 33784 16176
rect 30524 16136 33784 16164
rect 30524 16124 30530 16136
rect 33778 16124 33784 16136
rect 33836 16124 33842 16176
rect 36633 16167 36691 16173
rect 36633 16164 36645 16167
rect 33981 16136 36645 16164
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 20625 16099 20683 16105
rect 19659 16068 20484 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 18340 16000 19441 16028
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 19705 16031 19763 16037
rect 19705 15997 19717 16031
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 11716 15864 14872 15892
rect 18046 15852 18052 15904
rect 18104 15892 18110 15904
rect 18782 15892 18788 15904
rect 18104 15864 18788 15892
rect 18104 15852 18110 15864
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19720 15892 19748 15991
rect 19794 15988 19800 16040
rect 19852 15988 19858 16040
rect 19889 16031 19947 16037
rect 19889 15997 19901 16031
rect 19935 16028 19947 16031
rect 20254 16028 20260 16040
rect 19935 16000 20260 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 20456 16037 20484 16068
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 20714 16056 20720 16108
rect 20772 16056 20778 16108
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 21266 16096 21272 16108
rect 20947 16068 21272 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21266 16056 21272 16068
rect 21324 16096 21330 16108
rect 21726 16096 21732 16108
rect 21324 16068 21732 16096
rect 21324 16056 21330 16068
rect 21726 16056 21732 16068
rect 21784 16056 21790 16108
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22261 16099 22319 16105
rect 22261 16096 22273 16099
rect 22152 16068 22273 16096
rect 22152 16056 22158 16068
rect 22261 16065 22273 16068
rect 22307 16065 22319 16099
rect 22261 16059 22319 16065
rect 24486 16056 24492 16108
rect 24544 16056 24550 16108
rect 24670 16056 24676 16108
rect 24728 16056 24734 16108
rect 25682 16056 25688 16108
rect 25740 16096 25746 16108
rect 25869 16099 25927 16105
rect 25869 16096 25881 16099
rect 25740 16068 25881 16096
rect 25740 16056 25746 16068
rect 25869 16065 25881 16068
rect 25915 16065 25927 16099
rect 25869 16059 25927 16065
rect 26142 16056 26148 16108
rect 26200 16056 26206 16108
rect 29454 16056 29460 16108
rect 29512 16056 29518 16108
rect 29914 16056 29920 16108
rect 29972 16096 29978 16108
rect 30561 16099 30619 16105
rect 30561 16096 30573 16099
rect 29972 16068 30573 16096
rect 29972 16056 29978 16068
rect 30561 16065 30573 16068
rect 30607 16065 30619 16099
rect 30561 16059 30619 16065
rect 20441 16031 20499 16037
rect 20441 15997 20453 16031
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 20714 15892 20720 15904
rect 19720 15864 20720 15892
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 20824 15892 20852 15991
rect 21082 15988 21088 16040
rect 21140 16028 21146 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21140 16000 22017 16028
rect 21140 15988 21146 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 26605 16031 26663 16037
rect 26605 15997 26617 16031
rect 26651 15997 26663 16031
rect 30576 16028 30604 16059
rect 30742 16056 30748 16108
rect 30800 16056 30806 16108
rect 33134 16056 33140 16108
rect 33192 16096 33198 16108
rect 33870 16096 33876 16108
rect 33192 16068 33876 16096
rect 33192 16056 33198 16068
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 33981 16105 34009 16136
rect 36633 16133 36645 16136
rect 36679 16164 36691 16167
rect 37458 16164 37464 16176
rect 36679 16136 37464 16164
rect 36679 16133 36691 16136
rect 36633 16127 36691 16133
rect 37458 16124 37464 16136
rect 37516 16124 37522 16176
rect 37642 16164 37648 16176
rect 37700 16173 37706 16176
rect 37700 16167 37719 16173
rect 37568 16136 37648 16164
rect 33966 16099 34024 16105
rect 33966 16065 33978 16099
rect 34012 16065 34024 16099
rect 33966 16059 34024 16065
rect 34054 16056 34060 16108
rect 34112 16096 34118 16108
rect 34149 16099 34207 16105
rect 34149 16096 34161 16099
rect 34112 16068 34161 16096
rect 34112 16056 34118 16068
rect 34149 16065 34161 16068
rect 34195 16065 34207 16099
rect 34149 16059 34207 16065
rect 34238 16056 34244 16108
rect 34296 16056 34302 16108
rect 34379 16099 34437 16105
rect 34379 16065 34391 16099
rect 34425 16096 34437 16099
rect 34514 16096 34520 16108
rect 34425 16068 34520 16096
rect 34425 16065 34437 16068
rect 34379 16059 34437 16065
rect 34514 16056 34520 16068
rect 34572 16056 34578 16108
rect 36722 16056 36728 16108
rect 36780 16096 36786 16108
rect 36817 16099 36875 16105
rect 36817 16096 36829 16099
rect 36780 16068 36829 16096
rect 36780 16056 36786 16068
rect 36817 16065 36829 16068
rect 36863 16065 36875 16099
rect 36817 16059 36875 16065
rect 36909 16099 36967 16105
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37568 16096 37596 16136
rect 37642 16124 37648 16136
rect 37707 16133 37719 16167
rect 43714 16164 43720 16176
rect 37700 16127 37719 16133
rect 41386 16136 43720 16164
rect 37700 16124 37706 16127
rect 36955 16068 37596 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 36924 16028 36952 16059
rect 40218 16056 40224 16108
rect 40276 16056 40282 16108
rect 40497 16099 40555 16105
rect 40497 16065 40509 16099
rect 40543 16096 40555 16099
rect 41386 16096 41414 16136
rect 43714 16124 43720 16136
rect 43772 16124 43778 16176
rect 40543 16068 41414 16096
rect 40543 16065 40555 16068
rect 40497 16059 40555 16065
rect 43530 16056 43536 16108
rect 43588 16056 43594 16108
rect 43622 16056 43628 16108
rect 43680 16096 43686 16108
rect 43680 16068 43725 16096
rect 43680 16056 43686 16068
rect 43806 16056 43812 16108
rect 43864 16056 43870 16108
rect 43916 16105 43944 16204
rect 44910 16192 44916 16204
rect 44968 16192 44974 16244
rect 45554 16192 45560 16244
rect 45612 16192 45618 16244
rect 43901 16099 43959 16105
rect 43901 16065 43913 16099
rect 43947 16065 43959 16099
rect 43901 16059 43959 16065
rect 43990 16056 43996 16108
rect 44048 16105 44054 16108
rect 44048 16096 44056 16105
rect 46017 16099 46075 16105
rect 46017 16096 46029 16099
rect 44048 16068 44093 16096
rect 44192 16068 46029 16096
rect 44048 16059 44056 16068
rect 44048 16056 44054 16059
rect 30576 16000 36952 16028
rect 26605 15991 26663 15997
rect 26620 15960 26648 15991
rect 38102 15988 38108 16040
rect 38160 16028 38166 16040
rect 44192 16028 44220 16068
rect 46017 16065 46029 16068
rect 46063 16065 46075 16099
rect 46017 16059 46075 16065
rect 38160 16000 44220 16028
rect 38160 15988 38166 16000
rect 45738 15988 45744 16040
rect 45796 15988 45802 16040
rect 45830 15988 45836 16040
rect 45888 15988 45894 16040
rect 45925 16031 45983 16037
rect 45925 15997 45937 16031
rect 45971 15997 45983 16031
rect 45925 15991 45983 15997
rect 36262 15960 36268 15972
rect 26620 15932 36268 15960
rect 36262 15920 36268 15932
rect 36320 15920 36326 15972
rect 36722 15920 36728 15972
rect 36780 15960 36786 15972
rect 36780 15932 37688 15960
rect 36780 15920 36786 15932
rect 22002 15892 22008 15904
rect 20824 15864 22008 15892
rect 22002 15852 22008 15864
rect 22060 15892 22066 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 22060 15864 23397 15892
rect 22060 15852 22066 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 24581 15895 24639 15901
rect 24581 15861 24593 15895
rect 24627 15892 24639 15895
rect 24670 15892 24676 15904
rect 24627 15864 24676 15892
rect 24627 15861 24639 15864
rect 24581 15855 24639 15861
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 30190 15852 30196 15904
rect 30248 15892 30254 15904
rect 30561 15895 30619 15901
rect 30561 15892 30573 15895
rect 30248 15864 30573 15892
rect 30248 15852 30254 15864
rect 30561 15861 30573 15864
rect 30607 15861 30619 15895
rect 30561 15855 30619 15861
rect 33870 15852 33876 15904
rect 33928 15892 33934 15904
rect 36078 15892 36084 15904
rect 33928 15864 36084 15892
rect 33928 15852 33934 15864
rect 36078 15852 36084 15864
rect 36136 15852 36142 15904
rect 36633 15895 36691 15901
rect 36633 15861 36645 15895
rect 36679 15892 36691 15895
rect 36814 15892 36820 15904
rect 36679 15864 36820 15892
rect 36679 15861 36691 15864
rect 36633 15855 36691 15861
rect 36814 15852 36820 15864
rect 36872 15852 36878 15904
rect 37660 15901 37688 15932
rect 44174 15920 44180 15972
rect 44232 15920 44238 15972
rect 37645 15895 37703 15901
rect 37645 15861 37657 15895
rect 37691 15861 37703 15895
rect 37645 15855 37703 15861
rect 42978 15852 42984 15904
rect 43036 15892 43042 15904
rect 45940 15892 45968 15991
rect 43036 15864 45968 15892
rect 43036 15852 43042 15864
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7742 15688 7748 15700
rect 7423 15660 7748 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 11882 15688 11888 15700
rect 11756 15660 11888 15688
rect 11756 15648 11762 15660
rect 11882 15648 11888 15660
rect 11940 15688 11946 15700
rect 11940 15660 14780 15688
rect 11940 15648 11946 15660
rect 5626 15580 5632 15632
rect 5684 15620 5690 15632
rect 7926 15620 7932 15632
rect 5684 15592 7932 15620
rect 5684 15580 5690 15592
rect 7926 15580 7932 15592
rect 7984 15620 7990 15632
rect 14752 15620 14780 15660
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 14921 15691 14979 15697
rect 14921 15688 14933 15691
rect 14884 15660 14933 15688
rect 14884 15648 14890 15660
rect 14921 15657 14933 15660
rect 14967 15657 14979 15691
rect 14921 15651 14979 15657
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 21082 15688 21088 15700
rect 17552 15660 21088 15688
rect 17552 15648 17558 15660
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 22094 15648 22100 15700
rect 22152 15648 22158 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23440 15660 27936 15688
rect 23440 15648 23446 15660
rect 17034 15620 17040 15632
rect 7984 15592 14320 15620
rect 14752 15592 17040 15620
rect 7984 15580 7990 15592
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 7837 15555 7895 15561
rect 7837 15552 7849 15555
rect 6236 15524 7849 15552
rect 6236 15512 6242 15524
rect 7837 15521 7849 15524
rect 7883 15521 7895 15555
rect 7837 15515 7895 15521
rect 8018 15512 8024 15564
rect 8076 15512 8082 15564
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 14090 15484 14096 15496
rect 1627 15456 14096 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 14292 15493 14320 15592
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 27433 15623 27491 15629
rect 27433 15589 27445 15623
rect 27479 15620 27491 15623
rect 27798 15620 27804 15632
rect 27479 15592 27804 15620
rect 27479 15589 27491 15592
rect 27433 15583 27491 15589
rect 27798 15580 27804 15592
rect 27856 15580 27862 15632
rect 27908 15620 27936 15660
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 29733 15691 29791 15697
rect 29733 15688 29745 15691
rect 29144 15660 29745 15688
rect 29144 15648 29150 15660
rect 29733 15657 29745 15660
rect 29779 15657 29791 15691
rect 32398 15688 32404 15700
rect 29733 15651 29791 15657
rect 29840 15660 32404 15688
rect 29840 15620 29868 15660
rect 32398 15648 32404 15660
rect 32456 15688 32462 15700
rect 33042 15688 33048 15700
rect 32456 15660 33048 15688
rect 32456 15648 32462 15660
rect 33042 15648 33048 15660
rect 33100 15648 33106 15700
rect 33778 15648 33784 15700
rect 33836 15688 33842 15700
rect 33873 15691 33931 15697
rect 33873 15688 33885 15691
rect 33836 15660 33885 15688
rect 33836 15648 33842 15660
rect 33873 15657 33885 15660
rect 33919 15657 33931 15691
rect 33873 15651 33931 15657
rect 34146 15648 34152 15700
rect 34204 15688 34210 15700
rect 34514 15688 34520 15700
rect 34204 15660 34520 15688
rect 34204 15648 34210 15660
rect 34514 15648 34520 15660
rect 34572 15648 34578 15700
rect 40218 15688 40224 15700
rect 36004 15660 40224 15688
rect 27908 15592 29868 15620
rect 31018 15580 31024 15632
rect 31076 15620 31082 15632
rect 36004 15620 36032 15660
rect 40218 15648 40224 15660
rect 40276 15648 40282 15700
rect 36722 15620 36728 15632
rect 31076 15592 36032 15620
rect 36556 15592 36728 15620
rect 31076 15580 31082 15592
rect 14568 15524 17356 15552
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14425 15487 14483 15493
rect 14425 15453 14437 15487
rect 14471 15484 14483 15487
rect 14568 15484 14596 15524
rect 14471 15456 14596 15484
rect 14471 15453 14483 15456
rect 14425 15447 14483 15453
rect 14642 15444 14648 15496
rect 14700 15444 14706 15496
rect 14734 15444 14740 15496
rect 14792 15493 14798 15496
rect 14792 15484 14800 15493
rect 17328 15484 17356 15524
rect 17494 15512 17500 15564
rect 17552 15512 17558 15564
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 20165 15555 20223 15561
rect 20165 15552 20177 15555
rect 19852 15524 20177 15552
rect 19852 15512 19858 15524
rect 20165 15521 20177 15524
rect 20211 15552 20223 15555
rect 21174 15552 21180 15564
rect 20211 15524 21180 15552
rect 20211 15521 20223 15524
rect 20165 15515 20223 15521
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 22002 15512 22008 15564
rect 22060 15552 22066 15564
rect 22649 15555 22707 15561
rect 22649 15552 22661 15555
rect 22060 15524 22661 15552
rect 22060 15512 22066 15524
rect 22649 15521 22661 15524
rect 22695 15521 22707 15555
rect 27522 15552 27528 15564
rect 22649 15515 22707 15521
rect 26620 15524 27528 15552
rect 19058 15484 19064 15496
rect 14792 15456 14837 15484
rect 17328 15456 19064 15484
rect 14792 15447 14800 15456
rect 14792 15444 14798 15447
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 22094 15484 22100 15496
rect 21039 15456 22100 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1857 15419 1915 15425
rect 1857 15416 1869 15419
rect 992 15388 1869 15416
rect 992 15376 998 15388
rect 1857 15385 1869 15388
rect 1903 15385 1915 15419
rect 1857 15379 1915 15385
rect 2593 15419 2651 15425
rect 2593 15385 2605 15419
rect 2639 15385 2651 15419
rect 2593 15379 2651 15385
rect 2777 15419 2835 15425
rect 2777 15385 2789 15419
rect 2823 15416 2835 15419
rect 5534 15416 5540 15428
rect 2823 15388 5540 15416
rect 2823 15385 2835 15388
rect 2777 15379 2835 15385
rect 1026 15308 1032 15360
rect 1084 15348 1090 15360
rect 2608 15348 2636 15379
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 12434 15376 12440 15428
rect 12492 15416 12498 15428
rect 12802 15416 12808 15428
rect 12492 15388 12808 15416
rect 12492 15376 12498 15388
rect 12802 15376 12808 15388
rect 12860 15416 12866 15428
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 12860 15388 14565 15416
rect 12860 15376 12866 15388
rect 14553 15385 14565 15388
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 17764 15419 17822 15425
rect 17764 15385 17776 15419
rect 17810 15416 17822 15419
rect 19426 15416 19432 15428
rect 17810 15388 19432 15416
rect 17810 15385 17822 15388
rect 17764 15379 17822 15385
rect 19426 15376 19432 15388
rect 19484 15376 19490 15428
rect 19996 15416 20024 15447
rect 22094 15444 22100 15456
rect 22152 15444 22158 15496
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 22244 15456 22293 15484
rect 22244 15444 22250 15456
rect 22281 15453 22293 15456
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 22373 15487 22431 15493
rect 22373 15453 22385 15487
rect 22419 15484 22431 15487
rect 24581 15487 24639 15493
rect 22419 15456 23888 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 21266 15416 21272 15428
rect 19996 15388 21272 15416
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 22738 15376 22744 15428
rect 22796 15376 22802 15428
rect 23860 15416 23888 15456
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 26326 15484 26332 15496
rect 24627 15456 26332 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 24670 15416 24676 15428
rect 23860 15388 24676 15416
rect 24670 15376 24676 15388
rect 24728 15376 24734 15428
rect 24857 15419 24915 15425
rect 24857 15385 24869 15419
rect 24903 15416 24915 15419
rect 24946 15416 24952 15428
rect 24903 15388 24952 15416
rect 24903 15385 24915 15388
rect 24857 15379 24915 15385
rect 24946 15376 24952 15388
rect 25004 15416 25010 15428
rect 26620 15416 26648 15524
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 30742 15552 30748 15564
rect 30024 15524 30748 15552
rect 26694 15444 26700 15496
rect 26752 15484 26758 15496
rect 27709 15487 27767 15493
rect 27709 15484 27721 15487
rect 26752 15456 27721 15484
rect 26752 15444 26758 15456
rect 27709 15453 27721 15456
rect 27755 15453 27767 15487
rect 27709 15447 27767 15453
rect 29914 15444 29920 15496
rect 29972 15444 29978 15496
rect 30024 15493 30052 15524
rect 30742 15512 30748 15524
rect 30800 15552 30806 15564
rect 36556 15552 36584 15592
rect 36722 15580 36728 15592
rect 36780 15580 36786 15632
rect 36814 15580 36820 15632
rect 36872 15580 36878 15632
rect 36909 15623 36967 15629
rect 36909 15589 36921 15623
rect 36955 15620 36967 15623
rect 37274 15620 37280 15632
rect 36955 15592 37280 15620
rect 36955 15589 36967 15592
rect 36909 15583 36967 15589
rect 37274 15580 37280 15592
rect 37332 15580 37338 15632
rect 30800 15524 36584 15552
rect 30800 15512 30806 15524
rect 30009 15487 30067 15493
rect 30009 15453 30021 15487
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 30190 15444 30196 15496
rect 30248 15444 30254 15496
rect 30285 15487 30343 15493
rect 30285 15453 30297 15487
rect 30331 15453 30343 15487
rect 30285 15447 30343 15453
rect 25004 15388 26648 15416
rect 27433 15419 27491 15425
rect 25004 15376 25010 15388
rect 27433 15385 27445 15419
rect 27479 15416 27491 15419
rect 27522 15416 27528 15428
rect 27479 15388 27528 15416
rect 27479 15385 27491 15388
rect 27433 15379 27491 15385
rect 27522 15376 27528 15388
rect 27580 15376 27586 15428
rect 28074 15376 28080 15428
rect 28132 15416 28138 15428
rect 30300 15416 30328 15447
rect 33134 15444 33140 15496
rect 33192 15484 33198 15496
rect 33336 15493 33364 15524
rect 40310 15512 40316 15564
rect 40368 15552 40374 15564
rect 41141 15555 41199 15561
rect 41141 15552 41153 15555
rect 40368 15524 41153 15552
rect 40368 15512 40374 15524
rect 41141 15521 41153 15524
rect 41187 15521 41199 15555
rect 41141 15515 41199 15521
rect 33229 15487 33287 15493
rect 33229 15484 33241 15487
rect 33192 15456 33241 15484
rect 33192 15444 33198 15456
rect 33229 15453 33241 15456
rect 33275 15453 33287 15487
rect 33229 15447 33287 15453
rect 33322 15487 33380 15493
rect 33322 15453 33334 15487
rect 33368 15453 33380 15487
rect 33322 15447 33380 15453
rect 33686 15444 33692 15496
rect 33744 15493 33750 15496
rect 33744 15484 33752 15493
rect 34146 15484 34152 15496
rect 33744 15456 34152 15484
rect 33744 15447 33752 15456
rect 33744 15444 33750 15447
rect 34146 15444 34152 15456
rect 34204 15444 34210 15496
rect 36722 15444 36728 15496
rect 36780 15444 36786 15496
rect 37001 15487 37059 15493
rect 37001 15453 37013 15487
rect 37047 15484 37059 15487
rect 37047 15456 37136 15484
rect 37047 15453 37059 15456
rect 37001 15447 37059 15453
rect 28132 15388 30328 15416
rect 28132 15376 28138 15388
rect 33410 15376 33416 15428
rect 33468 15416 33474 15428
rect 33505 15419 33563 15425
rect 33505 15416 33517 15419
rect 33468 15388 33517 15416
rect 33468 15376 33474 15388
rect 33505 15385 33517 15388
rect 33551 15385 33563 15419
rect 33505 15379 33563 15385
rect 33597 15419 33655 15425
rect 33597 15385 33609 15419
rect 33643 15416 33655 15419
rect 34698 15416 34704 15428
rect 33643 15388 34704 15416
rect 33643 15385 33655 15388
rect 33597 15379 33655 15385
rect 1084 15320 2636 15348
rect 7745 15351 7803 15357
rect 1084 15308 1090 15320
rect 7745 15317 7757 15351
rect 7791 15348 7803 15351
rect 9306 15348 9312 15360
rect 7791 15320 9312 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 18877 15351 18935 15357
rect 18877 15348 18889 15351
rect 11572 15320 18889 15348
rect 11572 15308 11578 15320
rect 18877 15317 18889 15320
rect 18923 15348 18935 15351
rect 19978 15348 19984 15360
rect 18923 15320 19984 15348
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 27617 15351 27675 15357
rect 27617 15317 27629 15351
rect 27663 15348 27675 15351
rect 27706 15348 27712 15360
rect 27663 15320 27712 15348
rect 27663 15317 27675 15320
rect 27617 15311 27675 15317
rect 27706 15308 27712 15320
rect 27764 15308 27770 15360
rect 33520 15348 33548 15379
rect 34698 15376 34704 15388
rect 34756 15376 34762 15428
rect 35986 15376 35992 15428
rect 36044 15416 36050 15428
rect 36630 15416 36636 15428
rect 36044 15388 36636 15416
rect 36044 15376 36050 15388
rect 36630 15376 36636 15388
rect 36688 15416 36694 15428
rect 37108 15416 37136 15456
rect 36688 15388 37136 15416
rect 41408 15419 41466 15425
rect 36688 15376 36694 15388
rect 41408 15385 41420 15419
rect 41454 15416 41466 15419
rect 42610 15416 42616 15428
rect 41454 15388 42616 15416
rect 41454 15385 41466 15388
rect 41408 15379 41466 15385
rect 42610 15376 42616 15388
rect 42668 15376 42674 15428
rect 34054 15348 34060 15360
rect 33520 15320 34060 15348
rect 34054 15308 34060 15320
rect 34112 15308 34118 15360
rect 35894 15308 35900 15360
rect 35952 15348 35958 15360
rect 36541 15351 36599 15357
rect 36541 15348 36553 15351
rect 35952 15320 36553 15348
rect 35952 15308 35958 15320
rect 36541 15317 36553 15320
rect 36587 15317 36599 15351
rect 36541 15311 36599 15317
rect 36722 15308 36728 15360
rect 36780 15348 36786 15360
rect 37550 15348 37556 15360
rect 36780 15320 37556 15348
rect 36780 15308 36786 15320
rect 37550 15308 37556 15320
rect 37608 15308 37614 15360
rect 42521 15351 42579 15357
rect 42521 15317 42533 15351
rect 42567 15348 42579 15351
rect 43806 15348 43812 15360
rect 42567 15320 43812 15348
rect 42567 15317 42579 15320
rect 42521 15311 42579 15317
rect 43806 15308 43812 15320
rect 43864 15308 43870 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 11057 15147 11115 15153
rect 11057 15113 11069 15147
rect 11103 15144 11115 15147
rect 11238 15144 11244 15156
rect 11103 15116 11244 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 19484 15116 19533 15144
rect 19484 15104 19490 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 19521 15107 19579 15113
rect 19628 15116 20024 15144
rect 1118 15036 1124 15088
rect 1176 15076 1182 15088
rect 2958 15085 2964 15088
rect 1673 15079 1731 15085
rect 1673 15076 1685 15079
rect 1176 15048 1685 15076
rect 1176 15036 1182 15048
rect 1673 15045 1685 15048
rect 1719 15045 1731 15079
rect 2952 15076 2964 15085
rect 2919 15048 2964 15076
rect 1673 15039 1731 15045
rect 2952 15039 2964 15048
rect 2958 15036 2964 15039
rect 3016 15036 3022 15088
rect 11698 15076 11704 15088
rect 6886 15048 9628 15076
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 6886 15008 6914 15048
rect 7098 15017 7104 15020
rect 1903 14980 6914 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 7092 14971 7104 15017
rect 7098 14968 7104 14971
rect 7156 14968 7162 15020
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 2700 14804 2728 14903
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 3970 14804 3976 14816
rect 2700 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4890 14804 4896 14816
rect 4120 14776 4896 14804
rect 4120 14764 4126 14776
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14804 8263 14807
rect 8294 14804 8300 14816
rect 8251 14776 8300 14804
rect 8251 14773 8263 14776
rect 8205 14767 8263 14773
rect 8294 14764 8300 14776
rect 8352 14804 8358 14816
rect 9214 14804 9220 14816
rect 8352 14776 9220 14804
rect 8352 14764 8358 14776
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 9600 14804 9628 15048
rect 9692 15048 11704 15076
rect 9692 15017 9720 15048
rect 11698 15036 11704 15048
rect 11756 15076 11762 15088
rect 12342 15076 12348 15088
rect 11756 15048 12348 15076
rect 11756 15036 11762 15048
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9944 15011 10002 15017
rect 9944 14977 9956 15011
rect 9990 15008 10002 15011
rect 11790 15008 11796 15020
rect 9990 14980 11796 15008
rect 9990 14977 10002 14980
rect 9944 14971 10002 14977
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 19628 15008 19656 15116
rect 19886 15036 19892 15088
rect 19944 15036 19950 15088
rect 19996 15017 20024 15116
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 26605 15147 26663 15153
rect 26605 15144 26617 15147
rect 20772 15116 26617 15144
rect 20772 15104 20778 15116
rect 26605 15113 26617 15116
rect 26651 15113 26663 15147
rect 26605 15107 26663 15113
rect 27801 15147 27859 15153
rect 27801 15113 27813 15147
rect 27847 15144 27859 15147
rect 27847 15116 31064 15144
rect 27847 15113 27859 15116
rect 27801 15107 27859 15113
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 24118 15076 24124 15088
rect 22152 15048 24124 15076
rect 22152 15036 22158 15048
rect 24118 15036 24124 15048
rect 24176 15036 24182 15088
rect 28074 15036 28080 15088
rect 28132 15036 28138 15088
rect 31036 15085 31064 15116
rect 31128 15116 32996 15144
rect 31021 15079 31079 15085
rect 31021 15045 31033 15079
rect 31067 15045 31079 15079
rect 31021 15039 31079 15045
rect 18656 14980 19656 15008
rect 19705 15014 19763 15017
rect 19705 15011 19840 15014
rect 18656 14968 18662 14980
rect 19705 14977 19717 15011
rect 19751 15008 19840 15011
rect 19981 15011 20039 15017
rect 19751 14986 19932 15008
rect 19751 14977 19763 14986
rect 19812 14980 19932 14986
rect 19705 14971 19763 14977
rect 15010 14900 15016 14952
rect 15068 14940 15074 14952
rect 17494 14940 17500 14952
rect 15068 14912 17500 14940
rect 15068 14900 15074 14912
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 19904 14940 19932 14980
rect 19981 14977 19993 15011
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 21266 14968 21272 15020
rect 21324 15008 21330 15020
rect 23198 15008 23204 15020
rect 21324 14980 23204 15008
rect 21324 14968 21330 14980
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 23934 14968 23940 15020
rect 23992 14968 23998 15020
rect 24204 15011 24262 15017
rect 24204 14977 24216 15011
rect 24250 15008 24262 15011
rect 24762 15008 24768 15020
rect 24250 14980 24768 15008
rect 24250 14977 24262 14980
rect 24204 14971 24262 14977
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 25498 14968 25504 15020
rect 25556 15008 25562 15020
rect 25961 15011 26019 15017
rect 25961 15008 25973 15011
rect 25556 14980 25973 15008
rect 25556 14968 25562 14980
rect 25961 14977 25973 14980
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 26109 15011 26167 15017
rect 26109 14977 26121 15011
rect 26155 14977 26167 15011
rect 26109 14971 26167 14977
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26329 15011 26387 15017
rect 26329 14977 26341 15011
rect 26375 14977 26387 15011
rect 26329 14971 26387 14977
rect 22833 14943 22891 14949
rect 22833 14940 22845 14943
rect 19904 14912 22845 14940
rect 22833 14909 22845 14912
rect 22879 14909 22891 14943
rect 22833 14903 22891 14909
rect 23014 14900 23020 14952
rect 23072 14900 23078 14952
rect 23109 14943 23167 14949
rect 23109 14909 23121 14943
rect 23155 14909 23167 14943
rect 23109 14903 23167 14909
rect 11330 14832 11336 14884
rect 11388 14872 11394 14884
rect 22922 14872 22928 14884
rect 11388 14844 22928 14872
rect 11388 14832 11394 14844
rect 22922 14832 22928 14844
rect 22980 14832 22986 14884
rect 23124 14872 23152 14903
rect 23290 14900 23296 14952
rect 23348 14900 23354 14952
rect 26124 14940 26152 14971
rect 25332 14912 26152 14940
rect 25332 14884 25360 14912
rect 23124 14844 23980 14872
rect 12250 14804 12256 14816
rect 9600 14776 12256 14804
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 23842 14804 23848 14816
rect 13504 14776 23848 14804
rect 13504 14764 13510 14776
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 23952 14804 23980 14844
rect 25314 14832 25320 14884
rect 25372 14832 25378 14884
rect 26252 14872 26280 14971
rect 26344 14940 26372 14971
rect 26418 14968 26424 15020
rect 26476 15017 26482 15020
rect 26476 15008 26484 15017
rect 26476 14980 26521 15008
rect 26476 14971 26484 14980
rect 26476 14968 26482 14971
rect 27798 14968 27804 15020
rect 27856 14968 27862 15020
rect 27893 15011 27951 15017
rect 27893 14977 27905 15011
rect 27939 15008 27951 15011
rect 28994 15008 29000 15020
rect 27939 14980 29000 15008
rect 27939 14977 27951 14980
rect 27893 14971 27951 14977
rect 28994 14968 29000 14980
rect 29052 15008 29058 15020
rect 29914 15008 29920 15020
rect 29052 14980 29920 15008
rect 29052 14968 29058 14980
rect 29914 14968 29920 14980
rect 29972 14968 29978 15020
rect 27338 14940 27344 14952
rect 26344 14912 27344 14940
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 27614 14900 27620 14952
rect 27672 14940 27678 14952
rect 31128 14940 31156 15116
rect 31389 15079 31447 15085
rect 31389 15045 31401 15079
rect 31435 15076 31447 15079
rect 32554 15079 32612 15085
rect 32554 15076 32566 15079
rect 31435 15048 32566 15076
rect 31435 15045 31447 15048
rect 31389 15039 31447 15045
rect 32554 15045 32566 15048
rect 32600 15045 32612 15079
rect 32554 15039 32612 15045
rect 31202 14968 31208 15020
rect 31260 14968 31266 15020
rect 31294 14968 31300 15020
rect 31352 15008 31358 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 31352 14980 32321 15008
rect 31352 14968 31358 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32968 15008 32996 15116
rect 35820 15116 37872 15144
rect 33042 15036 33048 15088
rect 33100 15076 33106 15088
rect 35820 15076 35848 15116
rect 36523 15079 36581 15085
rect 36523 15076 36535 15079
rect 33100 15048 35848 15076
rect 35912 15048 36535 15076
rect 33100 15036 33106 15048
rect 32968 14980 33824 15008
rect 32309 14971 32367 14977
rect 27672 14912 31156 14940
rect 27672 14900 27678 14912
rect 28626 14872 28632 14884
rect 26252 14844 28632 14872
rect 28626 14832 28632 14844
rect 28684 14832 28690 14884
rect 27614 14804 27620 14816
rect 23952 14776 27620 14804
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 30190 14764 30196 14816
rect 30248 14804 30254 14816
rect 33318 14804 33324 14816
rect 30248 14776 33324 14804
rect 30248 14764 30254 14776
rect 33318 14764 33324 14776
rect 33376 14804 33382 14816
rect 33689 14807 33747 14813
rect 33689 14804 33701 14807
rect 33376 14776 33701 14804
rect 33376 14764 33382 14776
rect 33689 14773 33701 14776
rect 33735 14773 33747 14807
rect 33796 14804 33824 14980
rect 35802 14968 35808 15020
rect 35860 14968 35866 15020
rect 34514 14900 34520 14952
rect 34572 14940 34578 14952
rect 35912 14940 35940 15048
rect 36523 15045 36535 15048
rect 36569 15045 36581 15079
rect 37844 15076 37872 15116
rect 38838 15104 38844 15156
rect 38896 15104 38902 15156
rect 42610 15104 42616 15156
rect 42668 15104 42674 15156
rect 42978 15104 42984 15156
rect 43036 15104 43042 15156
rect 43806 15104 43812 15156
rect 43864 15144 43870 15156
rect 43864 15116 45140 15144
rect 43864 15104 43870 15116
rect 37844 15048 41414 15076
rect 36523 15039 36581 15045
rect 35989 15011 36047 15017
rect 35989 14977 36001 15011
rect 36035 14977 36047 15011
rect 35989 14971 36047 14977
rect 34572 14912 35940 14940
rect 36004 14940 36032 14971
rect 37182 14968 37188 15020
rect 37240 15008 37246 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 37240 14980 37473 15008
rect 37240 14968 37246 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37717 15011 37775 15017
rect 37717 15008 37729 15011
rect 37461 14971 37519 14977
rect 37568 14980 37729 15008
rect 36446 14940 36452 14952
rect 36004 14912 36452 14940
rect 34572 14900 34578 14912
rect 36446 14900 36452 14912
rect 36504 14940 36510 14952
rect 36817 14943 36875 14949
rect 36817 14940 36829 14943
rect 36504 14912 36829 14940
rect 36504 14900 36510 14912
rect 36817 14909 36829 14912
rect 36863 14909 36875 14943
rect 37568 14940 37596 14980
rect 37717 14977 37729 14980
rect 37763 14977 37775 15011
rect 41386 15008 41414 15048
rect 43898 15036 43904 15088
rect 43956 15076 43962 15088
rect 43993 15079 44051 15085
rect 43993 15076 44005 15079
rect 43956 15048 44005 15076
rect 43956 15036 43962 15048
rect 43993 15045 44005 15048
rect 44039 15045 44051 15079
rect 43993 15039 44051 15045
rect 42797 15011 42855 15017
rect 42797 15008 42809 15011
rect 41386 14980 42809 15008
rect 37717 14971 37775 14977
rect 42797 14977 42809 14980
rect 42843 14977 42855 15011
rect 42797 14971 42855 14977
rect 43073 15011 43131 15017
rect 43073 14977 43085 15011
rect 43119 14977 43131 15011
rect 43073 14971 43131 14977
rect 36817 14903 36875 14909
rect 37467 14912 37596 14940
rect 43088 14940 43116 14971
rect 43714 14968 43720 15020
rect 43772 14968 43778 15020
rect 43806 14968 43812 15020
rect 43864 15008 43870 15020
rect 43864 14980 43909 15008
rect 43864 14968 43870 14980
rect 44082 14968 44088 15020
rect 44140 14968 44146 15020
rect 44174 14968 44180 15020
rect 44232 15017 44238 15020
rect 45112 15017 45140 15116
rect 44232 15008 44240 15017
rect 45097 15011 45155 15017
rect 44232 14980 44277 15008
rect 44232 14971 44240 14980
rect 45097 14977 45109 15011
rect 45143 14977 45155 15011
rect 45097 14971 45155 14977
rect 44232 14968 44238 14971
rect 45189 14943 45247 14949
rect 43088 14912 44680 14940
rect 35805 14875 35863 14881
rect 35805 14841 35817 14875
rect 35851 14872 35863 14875
rect 37467 14872 37495 14912
rect 44361 14875 44419 14881
rect 44361 14872 44373 14875
rect 35851 14844 37495 14872
rect 41386 14844 44373 14872
rect 35851 14841 35863 14844
rect 35805 14835 35863 14841
rect 41386 14804 41414 14844
rect 44361 14841 44373 14844
rect 44407 14841 44419 14875
rect 44652 14872 44680 14912
rect 45189 14909 45201 14943
rect 45235 14940 45247 14943
rect 45278 14940 45284 14952
rect 45235 14912 45284 14940
rect 45235 14909 45247 14912
rect 45189 14903 45247 14909
rect 45278 14900 45284 14912
rect 45336 14900 45342 14952
rect 45465 14875 45523 14881
rect 45465 14872 45477 14875
rect 44652 14844 45477 14872
rect 44361 14835 44419 14841
rect 45465 14841 45477 14844
rect 45511 14841 45523 14875
rect 45465 14835 45523 14841
rect 33796 14776 41414 14804
rect 33689 14767 33747 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7098 14600 7104 14612
rect 7055 14572 7104 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 11790 14560 11796 14612
rect 11848 14560 11854 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 33778 14600 33784 14612
rect 12032 14572 33784 14600
rect 12032 14560 12038 14572
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 36630 14560 36636 14612
rect 36688 14560 36694 14612
rect 36998 14560 37004 14612
rect 37056 14600 37062 14612
rect 40310 14600 40316 14612
rect 37056 14572 40316 14600
rect 37056 14560 37062 14572
rect 40310 14560 40316 14572
rect 40368 14560 40374 14612
rect 11238 14492 11244 14544
rect 11296 14492 11302 14544
rect 12713 14535 12771 14541
rect 12713 14501 12725 14535
rect 12759 14532 12771 14535
rect 16206 14532 16212 14544
rect 12759 14504 16212 14532
rect 12759 14501 12771 14504
rect 12713 14495 12771 14501
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 17494 14492 17500 14544
rect 17552 14532 17558 14544
rect 17589 14535 17647 14541
rect 17589 14532 17601 14535
rect 17552 14504 17601 14532
rect 17552 14492 17558 14504
rect 17589 14501 17601 14504
rect 17635 14501 17647 14535
rect 17589 14495 17647 14501
rect 18233 14535 18291 14541
rect 18233 14501 18245 14535
rect 18279 14532 18291 14535
rect 18598 14532 18604 14544
rect 18279 14504 18604 14532
rect 18279 14501 18291 14504
rect 18233 14495 18291 14501
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 24670 14492 24676 14544
rect 24728 14492 24734 14544
rect 24762 14492 24768 14544
rect 24820 14492 24826 14544
rect 26234 14492 26240 14544
rect 26292 14532 26298 14544
rect 26694 14532 26700 14544
rect 26292 14504 26700 14532
rect 26292 14492 26298 14504
rect 26694 14492 26700 14504
rect 26752 14492 26758 14544
rect 26789 14535 26847 14541
rect 26789 14501 26801 14535
rect 26835 14501 26847 14535
rect 26789 14495 26847 14501
rect 934 14424 940 14476
rect 992 14464 998 14476
rect 992 14436 2636 14464
rect 992 14424 998 14436
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 2498 14396 2504 14408
rect 1627 14368 2504 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2608 14405 2636 14436
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 6822 14464 6828 14476
rect 4028 14436 6828 14464
rect 4028 14424 4034 14436
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 7650 14464 7656 14476
rect 7432 14436 7656 14464
rect 7432 14424 7438 14436
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 11256 14464 11284 14492
rect 11256 14436 11560 14464
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4120 14368 4261 14396
rect 4120 14356 4126 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 5592 14368 7481 14396
rect 5592 14356 5598 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 11146 14356 11152 14408
rect 11204 14356 11210 14408
rect 11330 14405 11336 14408
rect 11297 14399 11336 14405
rect 11297 14365 11309 14399
rect 11297 14359 11336 14365
rect 11330 14356 11336 14359
rect 11388 14356 11394 14408
rect 11532 14405 11560 14436
rect 11808 14436 13400 14464
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 11655 14399 11713 14405
rect 11655 14365 11667 14399
rect 11701 14396 11713 14399
rect 11808 14396 11836 14436
rect 12802 14396 12808 14408
rect 11701 14368 11836 14396
rect 11900 14368 12808 14396
rect 11701 14365 11713 14368
rect 11655 14359 11713 14365
rect 934 14288 940 14340
rect 992 14328 998 14340
rect 1857 14331 1915 14337
rect 1857 14328 1869 14331
rect 992 14300 1869 14328
rect 992 14288 998 14300
rect 1857 14297 1869 14300
rect 1903 14297 1915 14331
rect 1857 14291 1915 14297
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 3786 14328 3792 14340
rect 2823 14300 3792 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 3786 14288 3792 14300
rect 3844 14288 3850 14340
rect 5626 14288 5632 14340
rect 5684 14328 5690 14340
rect 8202 14328 8208 14340
rect 5684 14300 8208 14328
rect 5684 14288 5690 14300
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 10778 14288 10784 14340
rect 10836 14328 10842 14340
rect 11425 14331 11483 14337
rect 11425 14328 11437 14331
rect 10836 14300 11437 14328
rect 10836 14288 10842 14300
rect 11425 14297 11437 14300
rect 11471 14328 11483 14331
rect 11900 14328 11928 14368
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 13372 14396 13400 14436
rect 13446 14424 13452 14476
rect 13504 14424 13510 14476
rect 24857 14467 24915 14473
rect 24857 14433 24869 14467
rect 24903 14464 24915 14467
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 24903 14436 25697 14464
rect 24903 14433 24915 14436
rect 24857 14427 24915 14433
rect 25685 14433 25697 14436
rect 25731 14433 25743 14467
rect 26804 14464 26832 14495
rect 28626 14492 28632 14544
rect 28684 14532 28690 14544
rect 33410 14532 33416 14544
rect 28684 14504 33416 14532
rect 28684 14492 28690 14504
rect 33410 14492 33416 14504
rect 33468 14492 33474 14544
rect 40129 14535 40187 14541
rect 40129 14501 40141 14535
rect 40175 14501 40187 14535
rect 40129 14495 40187 14501
rect 25685 14427 25743 14433
rect 25884 14436 26832 14464
rect 14918 14396 14924 14408
rect 13372 14368 14924 14396
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 17494 14396 17500 14408
rect 16255 14368 17500 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16592 14340 16620 14368
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 18046 14356 18052 14408
rect 18104 14356 18110 14408
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14396 24639 14399
rect 24946 14396 24952 14408
rect 24627 14368 24952 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 24946 14356 24952 14368
rect 25004 14356 25010 14408
rect 25884 14405 25912 14436
rect 26878 14424 26884 14476
rect 26936 14424 26942 14476
rect 27706 14464 27712 14476
rect 26988 14436 27712 14464
rect 25869 14399 25927 14405
rect 25869 14365 25881 14399
rect 25915 14365 25927 14399
rect 25869 14359 25927 14365
rect 26145 14399 26203 14405
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26234 14396 26240 14408
rect 26191 14368 26240 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 26602 14356 26608 14408
rect 26660 14396 26666 14408
rect 26988 14396 27016 14436
rect 27706 14424 27712 14436
rect 27764 14424 27770 14476
rect 28261 14467 28319 14473
rect 28261 14433 28273 14467
rect 28307 14464 28319 14467
rect 28994 14464 29000 14476
rect 28307 14436 29000 14464
rect 28307 14433 28319 14436
rect 28261 14427 28319 14433
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 31205 14467 31263 14473
rect 31205 14433 31217 14467
rect 31251 14464 31263 14467
rect 31386 14464 31392 14476
rect 31251 14436 31392 14464
rect 31251 14433 31263 14436
rect 31205 14427 31263 14433
rect 31386 14424 31392 14436
rect 31444 14424 31450 14476
rect 40144 14464 40172 14495
rect 40218 14492 40224 14544
rect 40276 14532 40282 14544
rect 40276 14504 41368 14532
rect 40276 14492 40282 14504
rect 40144 14436 41184 14464
rect 30098 14396 30104 14408
rect 26660 14368 27016 14396
rect 27448 14368 30104 14396
rect 26660 14356 26666 14368
rect 12897 14331 12955 14337
rect 12897 14328 12909 14331
rect 11471 14300 11928 14328
rect 12406 14300 12909 14328
rect 11471 14297 11483 14300
rect 11425 14291 11483 14297
rect 7377 14263 7435 14269
rect 7377 14229 7389 14263
rect 7423 14260 7435 14263
rect 8294 14260 8300 14272
rect 7423 14232 8300 14260
rect 7423 14229 7435 14232
rect 7377 14223 7435 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 12158 14260 12164 14272
rect 11204 14232 12164 14260
rect 11204 14220 11210 14232
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 12250 14220 12256 14272
rect 12308 14260 12314 14272
rect 12406 14260 12434 14300
rect 12897 14297 12909 14300
rect 12943 14297 12955 14331
rect 12897 14291 12955 14297
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 16298 14328 16304 14340
rect 13688 14300 16304 14328
rect 13688 14288 13694 14300
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 16482 14337 16488 14340
rect 16476 14291 16488 14337
rect 16482 14288 16488 14291
rect 16540 14288 16546 14340
rect 16574 14288 16580 14340
rect 16632 14288 16638 14340
rect 16684 14300 18368 14328
rect 12308 14232 12434 14260
rect 12308 14220 12314 14232
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 16684 14260 16712 14300
rect 15160 14232 16712 14260
rect 18340 14260 18368 14300
rect 21910 14288 21916 14340
rect 21968 14328 21974 14340
rect 22005 14331 22063 14337
rect 22005 14328 22017 14331
rect 21968 14300 22017 14328
rect 21968 14288 21974 14300
rect 22005 14297 22017 14300
rect 22051 14297 22063 14331
rect 27448 14328 27476 14368
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 30558 14356 30564 14408
rect 30616 14396 30622 14408
rect 30742 14396 30748 14408
rect 30616 14368 30748 14396
rect 30616 14356 30622 14368
rect 30742 14356 30748 14368
rect 30800 14396 30806 14408
rect 30929 14399 30987 14405
rect 30929 14396 30941 14399
rect 30800 14368 30941 14396
rect 30800 14356 30806 14368
rect 30929 14365 30941 14368
rect 30975 14365 30987 14399
rect 30929 14359 30987 14365
rect 35618 14356 35624 14408
rect 35676 14396 35682 14408
rect 36541 14399 36599 14405
rect 36541 14396 36553 14399
rect 35676 14368 36553 14396
rect 35676 14356 35682 14368
rect 36541 14365 36553 14368
rect 36587 14365 36599 14399
rect 36541 14359 36599 14365
rect 36725 14399 36783 14405
rect 36725 14365 36737 14399
rect 36771 14396 36783 14399
rect 36998 14396 37004 14408
rect 36771 14368 37004 14396
rect 36771 14365 36783 14368
rect 36725 14359 36783 14365
rect 36998 14356 37004 14368
rect 37056 14356 37062 14408
rect 38838 14356 38844 14408
rect 38896 14396 38902 14408
rect 41156 14405 41184 14436
rect 41340 14405 41368 14504
rect 40405 14399 40463 14405
rect 40405 14396 40417 14399
rect 38896 14368 40417 14396
rect 38896 14356 38902 14368
rect 40405 14365 40417 14368
rect 40451 14365 40463 14399
rect 40405 14359 40463 14365
rect 41141 14399 41199 14405
rect 41141 14365 41153 14399
rect 41187 14365 41199 14399
rect 41141 14359 41199 14365
rect 41325 14399 41383 14405
rect 41325 14365 41337 14399
rect 41371 14365 41383 14399
rect 41325 14359 41383 14365
rect 22005 14291 22063 14297
rect 23308 14300 27476 14328
rect 23308 14269 23336 14300
rect 27522 14288 27528 14340
rect 27580 14288 27586 14340
rect 27801 14331 27859 14337
rect 27801 14328 27813 14331
rect 27632 14300 27813 14328
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 18340 14232 23305 14260
rect 15160 14220 15166 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 25314 14220 25320 14272
rect 25372 14260 25378 14272
rect 26053 14263 26111 14269
rect 26053 14260 26065 14263
rect 25372 14232 26065 14260
rect 25372 14220 25378 14232
rect 26053 14229 26065 14232
rect 26099 14260 26111 14263
rect 26602 14260 26608 14272
rect 26099 14232 26608 14260
rect 26099 14229 26111 14232
rect 26053 14223 26111 14229
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 27246 14220 27252 14272
rect 27304 14260 27310 14272
rect 27632 14260 27660 14300
rect 27801 14297 27813 14300
rect 27847 14297 27859 14331
rect 27801 14291 27859 14297
rect 27890 14288 27896 14340
rect 27948 14288 27954 14340
rect 29822 14288 29828 14340
rect 29880 14328 29886 14340
rect 31021 14331 31079 14337
rect 31021 14328 31033 14331
rect 29880 14300 31033 14328
rect 29880 14288 29886 14300
rect 31021 14297 31033 14300
rect 31067 14297 31079 14331
rect 31021 14291 31079 14297
rect 34514 14288 34520 14340
rect 34572 14328 34578 14340
rect 40034 14328 40040 14340
rect 34572 14300 40040 14328
rect 34572 14288 34578 14300
rect 40034 14288 40040 14300
rect 40092 14288 40098 14340
rect 40126 14288 40132 14340
rect 40184 14288 40190 14340
rect 44174 14328 44180 14340
rect 40236 14300 44180 14328
rect 27304 14232 27660 14260
rect 27304 14220 27310 14232
rect 27706 14220 27712 14272
rect 27764 14220 27770 14272
rect 28810 14220 28816 14272
rect 28868 14260 28874 14272
rect 30466 14260 30472 14272
rect 28868 14232 30472 14260
rect 28868 14220 28874 14232
rect 30466 14220 30472 14232
rect 30524 14220 30530 14272
rect 30558 14220 30564 14272
rect 30616 14220 30622 14272
rect 34238 14220 34244 14272
rect 34296 14260 34302 14272
rect 35802 14260 35808 14272
rect 34296 14232 35808 14260
rect 34296 14220 34302 14232
rect 35802 14220 35808 14232
rect 35860 14220 35866 14272
rect 36722 14220 36728 14272
rect 36780 14260 36786 14272
rect 40236 14260 40264 14300
rect 44174 14288 44180 14300
rect 44232 14288 44238 14340
rect 36780 14232 40264 14260
rect 36780 14220 36786 14232
rect 40310 14220 40316 14272
rect 40368 14220 40374 14272
rect 41233 14263 41291 14269
rect 41233 14229 41245 14263
rect 41279 14260 41291 14263
rect 41598 14260 41604 14272
rect 41279 14232 41604 14260
rect 41279 14229 41291 14232
rect 41233 14223 41291 14229
rect 41598 14220 41604 14232
rect 41656 14220 41662 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 4062 14016 4068 14068
rect 4120 14016 4126 14068
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 5626 14056 5632 14068
rect 4479 14028 5632 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 12986 14056 12992 14068
rect 10652 14028 12992 14056
rect 10652 14016 10658 14028
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 14090 14016 14096 14068
rect 14148 14056 14154 14068
rect 14826 14056 14832 14068
rect 14148 14028 14832 14056
rect 14148 14016 14154 14028
rect 14826 14016 14832 14028
rect 14884 14056 14890 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 14884 14028 15117 14056
rect 14884 14016 14890 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 16540 14028 17049 14056
rect 16540 14016 16546 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 17037 14019 17095 14025
rect 17402 14016 17408 14068
rect 17460 14016 17466 14068
rect 20901 14059 20959 14065
rect 20901 14025 20913 14059
rect 20947 14056 20959 14059
rect 21818 14056 21824 14068
rect 20947 14028 21824 14056
rect 20947 14025 20959 14028
rect 20901 14019 20959 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 23014 14016 23020 14068
rect 23072 14056 23078 14068
rect 23661 14059 23719 14065
rect 23661 14056 23673 14059
rect 23072 14028 23673 14056
rect 23072 14016 23078 14028
rect 23661 14025 23673 14028
rect 23707 14025 23719 14059
rect 23661 14019 23719 14025
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 30190 14056 30196 14068
rect 27580 14028 30196 14056
rect 27580 14016 27586 14028
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 30742 14016 30748 14068
rect 30800 14016 30806 14068
rect 33778 14016 33784 14068
rect 33836 14016 33842 14068
rect 38013 14059 38071 14065
rect 38013 14025 38025 14059
rect 38059 14025 38071 14059
rect 38013 14019 38071 14025
rect 3970 13988 3976 14000
rect 1688 13960 3976 13988
rect 1688 13929 1716 13960
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 10284 13960 12296 13988
rect 10284 13948 10290 13960
rect 1946 13929 1952 13932
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 1940 13883 1952 13929
rect 1946 13880 1952 13883
rect 2004 13880 2010 13932
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 4798 13920 4804 13932
rect 4571 13892 4804 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 8288 13923 8346 13929
rect 8288 13889 8300 13923
rect 8334 13920 8346 13923
rect 9122 13920 9128 13932
rect 8334 13892 9128 13920
rect 8334 13889 8346 13892
rect 8288 13883 8346 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 11974 13880 11980 13932
rect 12032 13880 12038 13932
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 12268 13920 12296 13960
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 16574 13988 16580 14000
rect 12400 13960 16580 13988
rect 12400 13948 12406 13960
rect 12713 13923 12771 13929
rect 12713 13920 12725 13923
rect 12268 13892 12725 13920
rect 12713 13889 12725 13892
rect 12759 13889 12771 13923
rect 13630 13920 13636 13932
rect 12713 13883 12771 13889
rect 12820 13892 13636 13920
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4755 13824 4844 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 2700 13756 3188 13784
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2700 13716 2728 13756
rect 2648 13688 2728 13716
rect 2648 13676 2654 13688
rect 3050 13676 3056 13728
rect 3108 13676 3114 13728
rect 3160 13716 3188 13756
rect 4816 13716 4844 13824
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 6880 13824 8033 13852
rect 6880 13812 6886 13824
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11664 13824 11713 13852
rect 11664 13812 11670 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 11882 13812 11888 13864
rect 11940 13812 11946 13864
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13852 12127 13855
rect 12820 13852 12848 13892
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 13740 13929 13768 13960
rect 16574 13948 16580 13960
rect 16632 13948 16638 14000
rect 18138 13988 18144 14000
rect 17144 13960 18144 13988
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 13992 13923 14050 13929
rect 13992 13889 14004 13923
rect 14038 13920 14050 13923
rect 14458 13920 14464 13932
rect 14038 13892 14464 13920
rect 14038 13889 14050 13892
rect 13992 13883 14050 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 17144 13920 17172 13960
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 23750 13988 23756 14000
rect 21192 13960 23756 13988
rect 16264 13892 17172 13920
rect 17221 13923 17279 13929
rect 16264 13880 16270 13892
rect 17221 13889 17233 13923
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17497 13923 17555 13929
rect 17497 13889 17509 13923
rect 17543 13920 17555 13923
rect 18598 13920 18604 13932
rect 17543 13892 18604 13920
rect 17543 13889 17555 13892
rect 17497 13883 17555 13889
rect 12115 13824 12848 13852
rect 12115 13821 12127 13824
rect 12069 13815 12127 13821
rect 12894 13812 12900 13864
rect 12952 13812 12958 13864
rect 17236 13852 17264 13883
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 21192 13929 21220 13960
rect 23750 13948 23756 13960
rect 23808 13948 23814 14000
rect 30282 13988 30288 14000
rect 29380 13960 30288 13988
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 21266 13880 21272 13932
rect 21324 13920 21330 13932
rect 21542 13920 21548 13932
rect 21324 13892 21548 13920
rect 21324 13880 21330 13892
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 22002 13880 22008 13932
rect 22060 13880 22066 13932
rect 23658 13880 23664 13932
rect 23716 13920 23722 13932
rect 23845 13923 23903 13929
rect 23845 13920 23857 13923
rect 23716 13892 23857 13920
rect 23716 13880 23722 13892
rect 23845 13889 23857 13892
rect 23891 13889 23903 13923
rect 23845 13883 23903 13889
rect 23934 13880 23940 13932
rect 23992 13880 23998 13932
rect 24029 13923 24087 13929
rect 24029 13889 24041 13923
rect 24075 13920 24087 13923
rect 24854 13920 24860 13932
rect 24075 13892 24860 13920
rect 24075 13889 24087 13892
rect 24029 13883 24087 13889
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 29380 13929 29408 13960
rect 30282 13948 30288 13960
rect 30340 13948 30346 14000
rect 33410 13948 33416 14000
rect 33468 13948 33474 14000
rect 37734 13948 37740 14000
rect 37792 13948 37798 14000
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13889 29423 13923
rect 29365 13883 29423 13889
rect 29632 13923 29690 13929
rect 29632 13889 29644 13923
rect 29678 13920 29690 13923
rect 29914 13920 29920 13932
rect 29678 13892 29920 13920
rect 29678 13889 29690 13892
rect 29632 13883 29690 13889
rect 29914 13880 29920 13892
rect 29972 13880 29978 13932
rect 33134 13920 33140 13932
rect 30392 13892 33140 13920
rect 20622 13852 20628 13864
rect 17236 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 21082 13812 21088 13864
rect 21140 13812 21146 13864
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 22189 13855 22247 13861
rect 22189 13852 22201 13855
rect 21407 13824 22201 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 22189 13821 22201 13824
rect 22235 13852 22247 13855
rect 23290 13852 23296 13864
rect 22235 13824 23296 13852
rect 22235 13821 22247 13824
rect 22189 13815 22247 13821
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 24118 13812 24124 13864
rect 24176 13812 24182 13864
rect 4982 13744 4988 13796
rect 5040 13784 5046 13796
rect 12158 13784 12164 13796
rect 5040 13756 8064 13784
rect 5040 13744 5046 13756
rect 7650 13716 7656 13728
rect 3160 13688 7656 13716
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 8036 13716 8064 13756
rect 8956 13756 12164 13784
rect 8956 13716 8984 13756
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 28994 13784 29000 13796
rect 14844 13756 29000 13784
rect 8036 13688 8984 13716
rect 9398 13676 9404 13728
rect 9456 13676 9462 13728
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 14844 13716 14872 13756
rect 28994 13744 29000 13756
rect 29052 13744 29058 13796
rect 12124 13688 14872 13716
rect 12124 13676 12130 13688
rect 17862 13676 17868 13728
rect 17920 13716 17926 13728
rect 22462 13716 22468 13728
rect 17920 13688 22468 13716
rect 17920 13676 17926 13688
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 28258 13676 28264 13728
rect 28316 13716 28322 13728
rect 30392 13716 30420 13892
rect 33134 13880 33140 13892
rect 33192 13880 33198 13932
rect 33318 13929 33324 13932
rect 33285 13923 33324 13929
rect 33285 13889 33297 13923
rect 33285 13883 33324 13889
rect 33318 13880 33324 13883
rect 33376 13880 33382 13932
rect 33502 13880 33508 13932
rect 33560 13880 33566 13932
rect 33594 13880 33600 13932
rect 33652 13929 33658 13932
rect 33652 13920 33660 13929
rect 33652 13892 33697 13920
rect 33652 13883 33660 13892
rect 33652 13880 33658 13883
rect 37458 13880 37464 13932
rect 37516 13880 37522 13932
rect 37642 13880 37648 13932
rect 37700 13880 37706 13932
rect 37829 13923 37887 13929
rect 37829 13889 37841 13923
rect 37875 13889 37887 13923
rect 38028 13920 38056 14019
rect 38102 14016 38108 14068
rect 38160 14056 38166 14068
rect 41049 14059 41107 14065
rect 41049 14056 41061 14059
rect 38160 14028 41061 14056
rect 38160 14016 38166 14028
rect 41049 14025 41061 14028
rect 41095 14025 41107 14059
rect 41049 14019 41107 14025
rect 40770 13988 40776 14000
rect 39684 13960 40776 13988
rect 39684 13929 39712 13960
rect 40770 13948 40776 13960
rect 40828 13948 40834 14000
rect 38841 13923 38899 13929
rect 38841 13920 38853 13923
rect 38028 13892 38853 13920
rect 37829 13883 37887 13889
rect 38841 13889 38853 13892
rect 38887 13889 38899 13923
rect 38841 13883 38899 13889
rect 39669 13923 39727 13929
rect 39669 13889 39681 13923
rect 39715 13889 39727 13923
rect 39925 13923 39983 13929
rect 39925 13920 39937 13923
rect 39669 13883 39727 13889
rect 39776 13892 39937 13920
rect 30466 13812 30472 13864
rect 30524 13852 30530 13864
rect 36722 13852 36728 13864
rect 30524 13824 36728 13852
rect 30524 13812 30530 13824
rect 36722 13812 36728 13824
rect 36780 13812 36786 13864
rect 32030 13744 32036 13796
rect 32088 13784 32094 13796
rect 32858 13784 32864 13796
rect 32088 13756 32864 13784
rect 32088 13744 32094 13756
rect 32858 13744 32864 13756
rect 32916 13784 32922 13796
rect 37844 13784 37872 13883
rect 38657 13855 38715 13861
rect 38657 13821 38669 13855
rect 38703 13852 38715 13855
rect 38930 13852 38936 13864
rect 38703 13824 38936 13852
rect 38703 13821 38715 13824
rect 38657 13815 38715 13821
rect 38930 13812 38936 13824
rect 38988 13812 38994 13864
rect 39025 13855 39083 13861
rect 39025 13821 39037 13855
rect 39071 13852 39083 13855
rect 39776 13852 39804 13892
rect 39925 13889 39937 13892
rect 39971 13889 39983 13923
rect 39925 13883 39983 13889
rect 39071 13824 39804 13852
rect 39071 13821 39083 13824
rect 39025 13815 39083 13821
rect 32916 13756 37872 13784
rect 32916 13744 32922 13756
rect 28316 13688 30420 13716
rect 28316 13676 28322 13688
rect 31478 13676 31484 13728
rect 31536 13716 31542 13728
rect 35986 13716 35992 13728
rect 31536 13688 35992 13716
rect 31536 13676 31542 13688
rect 35986 13676 35992 13688
rect 36044 13676 36050 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1946 13472 1952 13524
rect 2004 13472 2010 13524
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 4982 13512 4988 13524
rect 2556 13484 4988 13512
rect 2556 13472 2562 13484
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 9122 13472 9128 13524
rect 9180 13472 9186 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 11977 13515 12035 13521
rect 11977 13512 11989 13515
rect 11940 13484 11989 13512
rect 11940 13472 11946 13484
rect 11977 13481 11989 13484
rect 12023 13481 12035 13515
rect 11977 13475 12035 13481
rect 14458 13472 14464 13524
rect 14516 13472 14522 13524
rect 16224 13484 16712 13512
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 15378 13444 15384 13456
rect 8260 13416 15384 13444
rect 8260 13404 8266 13416
rect 2590 13336 2596 13388
rect 2648 13336 2654 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 12268 13385 12296 13416
rect 15378 13404 15384 13416
rect 15436 13404 15442 13456
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 7708 13348 9689 13376
rect 7708 13336 7714 13348
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13345 12311 13379
rect 12253 13339 12311 13345
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 12894 13376 12900 13388
rect 12483 13348 12900 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 12894 13336 12900 13348
rect 12952 13376 12958 13388
rect 13170 13376 13176 13388
rect 12952 13348 13176 13376
rect 12952 13336 12958 13348
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 16224 13376 16252 13484
rect 16574 13404 16580 13456
rect 16632 13404 16638 13456
rect 16684 13444 16712 13484
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 16942 13512 16948 13524
rect 16816 13484 16948 13512
rect 16816 13472 16822 13484
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 19150 13512 19156 13524
rect 17052 13484 19156 13512
rect 17052 13444 17080 13484
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21637 13515 21695 13521
rect 21637 13512 21649 13515
rect 21140 13484 21649 13512
rect 21140 13472 21146 13484
rect 21637 13481 21649 13484
rect 21683 13481 21695 13515
rect 21637 13475 21695 13481
rect 26694 13472 26700 13524
rect 26752 13512 26758 13524
rect 26970 13512 26976 13524
rect 26752 13484 26976 13512
rect 26752 13472 26758 13484
rect 26970 13472 26976 13484
rect 27028 13512 27034 13524
rect 27525 13515 27583 13521
rect 27525 13512 27537 13515
rect 27028 13484 27537 13512
rect 27028 13472 27034 13484
rect 27525 13481 27537 13484
rect 27571 13481 27583 13515
rect 27525 13475 27583 13481
rect 29914 13472 29920 13524
rect 29972 13472 29978 13524
rect 30285 13515 30343 13521
rect 30285 13481 30297 13515
rect 30331 13512 30343 13515
rect 30558 13512 30564 13524
rect 30331 13484 30564 13512
rect 30331 13481 30343 13484
rect 30285 13475 30343 13481
rect 30558 13472 30564 13484
rect 30616 13472 30622 13524
rect 53098 13512 53104 13524
rect 31726 13484 53104 13512
rect 16684 13416 17080 13444
rect 21928 13416 22784 13444
rect 14660 13348 16252 13376
rect 16393 13379 16451 13385
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 2455 13280 4261 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 4249 13277 4261 13280
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 5350 13268 5356 13320
rect 5408 13268 5414 13320
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 5902 13308 5908 13320
rect 5583 13280 5908 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 6822 13308 6828 13320
rect 6043 13280 6828 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 10134 13308 10140 13320
rect 9088 13280 10140 13308
rect 9088 13268 9094 13280
rect 10134 13268 10140 13280
rect 10192 13308 10198 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 10192 13280 12173 13308
rect 10192 13268 10198 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12342 13268 12348 13320
rect 12400 13268 12406 13320
rect 14660 13317 14688 13348
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 16592 13376 16620 13404
rect 16850 13376 16856 13388
rect 16439 13348 16856 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 21821 13379 21879 13385
rect 21821 13345 21833 13379
rect 21867 13376 21879 13379
rect 21928 13376 21956 13416
rect 21867 13348 21956 13376
rect 22005 13379 22063 13385
rect 21867 13345 21879 13348
rect 21821 13339 21879 13345
rect 22005 13345 22017 13379
rect 22051 13376 22063 13379
rect 22554 13376 22560 13388
rect 22051 13348 22560 13376
rect 22051 13345 22063 13348
rect 22005 13339 22063 13345
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14826 13268 14832 13320
rect 14884 13268 14890 13320
rect 14918 13268 14924 13320
rect 14976 13268 14982 13320
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 16666 13308 16672 13320
rect 16623 13280 16672 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 17494 13268 17500 13320
rect 17552 13268 17558 13320
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 21726 13308 21732 13320
rect 20864 13280 21732 13308
rect 20864 13268 20870 13280
rect 21726 13268 21732 13280
rect 21784 13308 21790 13320
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21784 13280 21925 13308
rect 21784 13268 21790 13280
rect 21913 13277 21925 13280
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 22094 13268 22100 13320
rect 22152 13268 22158 13320
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13277 22707 13311
rect 22756 13308 22784 13416
rect 22922 13404 22928 13456
rect 22980 13444 22986 13456
rect 31726 13444 31754 13484
rect 53098 13472 53104 13484
rect 53156 13472 53162 13524
rect 34606 13444 34612 13456
rect 22980 13416 31754 13444
rect 31956 13416 34612 13444
rect 22980 13404 22986 13416
rect 28994 13336 29000 13388
rect 29052 13376 29058 13388
rect 30190 13376 30196 13388
rect 29052 13348 30196 13376
rect 29052 13336 29058 13348
rect 30190 13336 30196 13348
rect 30248 13336 30254 13388
rect 30377 13379 30435 13385
rect 30377 13345 30389 13379
rect 30423 13376 30435 13379
rect 30929 13379 30987 13385
rect 30929 13376 30941 13379
rect 30423 13348 30941 13376
rect 30423 13345 30435 13348
rect 30377 13339 30435 13345
rect 30929 13345 30941 13348
rect 30975 13345 30987 13379
rect 31956 13376 31984 13416
rect 34606 13404 34612 13416
rect 34664 13444 34670 13456
rect 37458 13444 37464 13456
rect 34664 13416 37464 13444
rect 34664 13404 34670 13416
rect 30929 13339 30987 13345
rect 31680 13348 31984 13376
rect 22925 13311 22983 13317
rect 22925 13308 22937 13311
rect 22756 13280 22937 13308
rect 22649 13271 22707 13277
rect 22925 13277 22937 13280
rect 22971 13308 22983 13311
rect 23658 13308 23664 13320
rect 22971 13280 23664 13308
rect 22971 13277 22983 13280
rect 22925 13271 22983 13277
rect 934 13200 940 13252
rect 992 13240 998 13252
rect 3237 13243 3295 13249
rect 3237 13240 3249 13243
rect 992 13212 3249 13240
rect 992 13200 998 13212
rect 3237 13209 3249 13212
rect 3283 13209 3295 13243
rect 3237 13203 3295 13209
rect 4062 13200 4068 13252
rect 4120 13200 4126 13252
rect 5445 13243 5503 13249
rect 5445 13209 5457 13243
rect 5491 13240 5503 13243
rect 6242 13243 6300 13249
rect 6242 13240 6254 13243
rect 5491 13212 6254 13240
rect 5491 13209 5503 13212
rect 5445 13203 5503 13209
rect 6242 13209 6254 13212
rect 6288 13209 6300 13243
rect 6242 13203 6300 13209
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 12894 13240 12900 13252
rect 6420 13212 12900 13240
rect 6420 13200 6426 13212
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 17764 13243 17822 13249
rect 16592 13212 16712 13240
rect 2317 13175 2375 13181
rect 2317 13141 2329 13175
rect 2363 13172 2375 13175
rect 3050 13172 3056 13184
rect 2363 13144 3056 13172
rect 2363 13141 2375 13144
rect 2317 13135 2375 13141
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 3326 13132 3332 13184
rect 3384 13132 3390 13184
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9456 13144 9505 13172
rect 9456 13132 9462 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 16592 13172 16620 13212
rect 11020 13144 16620 13172
rect 16684 13172 16712 13212
rect 17764 13209 17776 13243
rect 17810 13240 17822 13243
rect 18506 13240 18512 13252
rect 17810 13212 18512 13240
rect 17810 13209 17822 13212
rect 17764 13203 17822 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 18616 13212 19012 13240
rect 18616 13172 18644 13212
rect 16684 13144 18644 13172
rect 11020 13132 11026 13144
rect 18874 13132 18880 13184
rect 18932 13132 18938 13184
rect 18984 13172 19012 13212
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 22664 13240 22692 13271
rect 23658 13268 23664 13280
rect 23716 13268 23722 13320
rect 27246 13268 27252 13320
rect 27304 13268 27310 13320
rect 27341 13311 27399 13317
rect 27341 13277 27353 13311
rect 27387 13308 27399 13311
rect 27890 13308 27896 13320
rect 27387 13280 27896 13308
rect 27387 13277 27399 13280
rect 27341 13271 27399 13277
rect 27890 13268 27896 13280
rect 27948 13268 27954 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30742 13308 30748 13320
rect 30147 13280 30748 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 31680 13317 31708 13348
rect 30837 13311 30895 13317
rect 30837 13277 30849 13311
rect 30883 13308 30895 13311
rect 31665 13311 31723 13317
rect 31665 13308 31677 13311
rect 30883 13280 31677 13308
rect 30883 13277 30895 13280
rect 30837 13271 30895 13277
rect 31665 13277 31677 13280
rect 31711 13277 31723 13311
rect 31665 13271 31723 13277
rect 32030 13268 32036 13320
rect 32088 13268 32094 13320
rect 35728 13317 35756 13416
rect 37458 13404 37464 13416
rect 37516 13404 37522 13456
rect 37274 13336 37280 13388
rect 37332 13376 37338 13388
rect 37369 13379 37427 13385
rect 37369 13376 37381 13379
rect 37332 13348 37381 13376
rect 37332 13336 37338 13348
rect 37369 13345 37381 13348
rect 37415 13345 37427 13379
rect 37369 13339 37427 13345
rect 35713 13311 35771 13317
rect 35713 13277 35725 13311
rect 35759 13277 35771 13311
rect 35713 13271 35771 13277
rect 35986 13268 35992 13320
rect 36044 13268 36050 13320
rect 36081 13311 36139 13317
rect 36081 13277 36093 13311
rect 36127 13277 36139 13311
rect 36081 13271 36139 13277
rect 21048 13212 22692 13240
rect 21048 13200 21054 13212
rect 23750 13200 23756 13252
rect 23808 13240 23814 13252
rect 27982 13240 27988 13252
rect 23808 13212 27988 13240
rect 23808 13200 23814 13212
rect 27982 13200 27988 13212
rect 28040 13200 28046 13252
rect 31846 13200 31852 13252
rect 31904 13200 31910 13252
rect 31941 13243 31999 13249
rect 31941 13209 31953 13243
rect 31987 13240 31999 13243
rect 32490 13240 32496 13252
rect 31987 13212 32496 13240
rect 31987 13209 31999 13212
rect 31941 13203 31999 13209
rect 32490 13200 32496 13212
rect 32548 13200 32554 13252
rect 35894 13200 35900 13252
rect 35952 13200 35958 13252
rect 36096 13240 36124 13271
rect 37090 13268 37096 13320
rect 37148 13268 37154 13320
rect 40770 13268 40776 13320
rect 40828 13308 40834 13320
rect 41322 13308 41328 13320
rect 40828 13280 41328 13308
rect 40828 13268 40834 13280
rect 41322 13268 41328 13280
rect 41380 13308 41386 13320
rect 41509 13311 41567 13317
rect 41509 13308 41521 13311
rect 41380 13280 41521 13308
rect 41380 13268 41386 13280
rect 41509 13277 41521 13280
rect 41555 13277 41567 13311
rect 41509 13271 41567 13277
rect 41598 13268 41604 13320
rect 41656 13308 41662 13320
rect 41765 13311 41823 13317
rect 41765 13308 41777 13311
rect 41656 13280 41777 13308
rect 41656 13268 41662 13280
rect 41765 13277 41777 13280
rect 41811 13277 41823 13311
rect 41765 13271 41823 13277
rect 37550 13240 37556 13252
rect 36096 13212 37556 13240
rect 37550 13200 37556 13212
rect 37608 13200 37614 13252
rect 27430 13172 27436 13184
rect 18984 13144 27436 13172
rect 27430 13132 27436 13144
rect 27488 13132 27494 13184
rect 31570 13132 31576 13184
rect 31628 13172 31634 13184
rect 32217 13175 32275 13181
rect 32217 13172 32229 13175
rect 31628 13144 32229 13172
rect 31628 13132 31634 13144
rect 32217 13141 32229 13144
rect 32263 13141 32275 13175
rect 32217 13135 32275 13141
rect 36262 13132 36268 13184
rect 36320 13132 36326 13184
rect 39850 13132 39856 13184
rect 39908 13172 39914 13184
rect 42889 13175 42947 13181
rect 42889 13172 42901 13175
rect 39908 13144 42901 13172
rect 39908 13132 39914 13144
rect 42889 13141 42901 13144
rect 42935 13172 42947 13175
rect 43806 13172 43812 13184
rect 42935 13144 43812 13172
rect 42935 13141 42947 13144
rect 42889 13135 42947 13141
rect 43806 13132 43812 13144
rect 43864 13132 43870 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 934 12928 940 12980
rect 992 12968 998 12980
rect 4062 12968 4068 12980
rect 992 12940 4068 12968
rect 992 12928 998 12940
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 8996 12940 9720 12968
rect 8996 12928 9002 12940
rect 1026 12860 1032 12912
rect 1084 12900 1090 12912
rect 2593 12903 2651 12909
rect 2593 12900 2605 12903
rect 1084 12872 2605 12900
rect 1084 12860 1090 12872
rect 2593 12869 2605 12872
rect 2639 12869 2651 12903
rect 2593 12863 2651 12869
rect 2777 12903 2835 12909
rect 2777 12869 2789 12903
rect 2823 12900 2835 12903
rect 9582 12900 9588 12912
rect 2823 12872 9588 12900
rect 2823 12869 2835 12872
rect 2777 12863 2835 12869
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 6362 12832 6368 12844
rect 1627 12804 6368 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 9030 12792 9036 12844
rect 9088 12792 9094 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9692 12832 9720 12940
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 10928 12940 12112 12968
rect 10928 12928 10934 12940
rect 10410 12832 10416 12844
rect 9539 12804 10416 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 11974 12841 11980 12844
rect 11968 12795 11980 12841
rect 11974 12792 11980 12795
rect 12032 12792 12038 12844
rect 12084 12832 12112 12940
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12400 12940 13093 12968
rect 12400 12928 12406 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 13081 12931 13139 12937
rect 16666 12928 16672 12980
rect 16724 12968 16730 12980
rect 16850 12968 16856 12980
rect 16724 12940 16856 12968
rect 16724 12928 16730 12940
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 18506 12928 18512 12980
rect 18564 12928 18570 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 18656 12940 19012 12968
rect 18656 12928 18662 12940
rect 12158 12860 12164 12912
rect 12216 12900 12222 12912
rect 18874 12900 18880 12912
rect 12216 12872 18880 12900
rect 12216 12860 12222 12872
rect 18874 12860 18880 12872
rect 18932 12860 18938 12912
rect 12084 12804 16804 12832
rect 934 12724 940 12776
rect 992 12764 998 12776
rect 1765 12767 1823 12773
rect 1765 12764 1777 12767
rect 992 12736 1777 12764
rect 992 12724 998 12736
rect 1765 12733 1777 12736
rect 1811 12733 1823 12767
rect 1765 12727 1823 12733
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 9125 12767 9183 12773
rect 3384 12736 9076 12764
rect 3384 12724 3390 12736
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 8938 12696 8944 12708
rect 3108 12668 8944 12696
rect 3108 12656 3114 12668
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 9048 12696 9076 12736
rect 9125 12733 9137 12767
rect 9171 12764 9183 12767
rect 9306 12764 9312 12776
rect 9171 12736 9312 12764
rect 9171 12733 9183 12736
rect 9125 12727 9183 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 16776 12696 16804 12804
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17218 12832 17224 12844
rect 17083 12804 17224 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17218 12792 17224 12804
rect 17276 12792 17282 12844
rect 18984 12841 19012 12940
rect 21726 12928 21732 12980
rect 21784 12968 21790 12980
rect 23934 12968 23940 12980
rect 21784 12940 23940 12968
rect 21784 12928 21790 12940
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 24854 12928 24860 12980
rect 24912 12928 24918 12980
rect 26418 12968 26424 12980
rect 26252 12940 26424 12968
rect 22094 12860 22100 12912
rect 22152 12900 22158 12912
rect 22646 12900 22652 12912
rect 22152 12872 22652 12900
rect 22152 12860 22158 12872
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 26252 12900 26280 12940
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 27430 12928 27436 12980
rect 27488 12968 27494 12980
rect 27617 12971 27675 12977
rect 27617 12968 27629 12971
rect 27488 12940 27629 12968
rect 27488 12928 27494 12940
rect 27617 12937 27629 12940
rect 27663 12937 27675 12971
rect 27617 12931 27675 12937
rect 23676 12872 26280 12900
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 18708 12764 18736 12795
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 22278 12792 22284 12844
rect 22336 12792 22342 12844
rect 23676 12832 23704 12872
rect 22480 12804 23704 12832
rect 23744 12835 23802 12841
rect 19426 12764 19432 12776
rect 18708 12736 19432 12764
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 22480 12696 22508 12804
rect 23744 12801 23756 12835
rect 23790 12832 23802 12835
rect 24578 12832 24584 12844
rect 23790 12804 24584 12832
rect 23790 12801 23802 12804
rect 23744 12795 23802 12801
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 25774 12792 25780 12844
rect 25832 12832 25838 12844
rect 25961 12835 26019 12841
rect 25961 12832 25973 12835
rect 25832 12804 25973 12832
rect 25832 12792 25838 12804
rect 25961 12801 25973 12804
rect 26007 12801 26019 12835
rect 25961 12795 26019 12801
rect 22554 12724 22560 12776
rect 22612 12724 22618 12776
rect 22649 12767 22707 12773
rect 22649 12733 22661 12767
rect 22695 12764 22707 12767
rect 22738 12764 22744 12776
rect 22695 12736 22744 12764
rect 22695 12733 22707 12736
rect 22649 12727 22707 12733
rect 22664 12696 22692 12727
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 23474 12724 23480 12776
rect 23532 12724 23538 12776
rect 26252 12764 26280 12872
rect 26326 12860 26332 12912
rect 26384 12860 26390 12912
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 27632 12832 27660 12931
rect 31846 12928 31852 12980
rect 31904 12968 31910 12980
rect 32769 12971 32827 12977
rect 32769 12968 32781 12971
rect 31904 12940 32781 12968
rect 31904 12928 31910 12940
rect 32769 12937 32781 12940
rect 32815 12937 32827 12971
rect 32769 12931 32827 12937
rect 34054 12928 34060 12980
rect 34112 12968 34118 12980
rect 37274 12968 37280 12980
rect 34112 12940 37280 12968
rect 34112 12928 34118 12940
rect 37274 12928 37280 12940
rect 37332 12928 37338 12980
rect 37461 12971 37519 12977
rect 37461 12937 37473 12971
rect 37507 12968 37519 12971
rect 37642 12968 37648 12980
rect 37507 12940 37648 12968
rect 37507 12937 37519 12940
rect 37461 12931 37519 12937
rect 37642 12928 37648 12940
rect 37700 12928 37706 12980
rect 37829 12971 37887 12977
rect 37829 12937 37841 12971
rect 37875 12968 37887 12971
rect 38102 12968 38108 12980
rect 37875 12940 38108 12968
rect 37875 12937 37887 12940
rect 37829 12931 37887 12937
rect 38102 12928 38108 12940
rect 38160 12928 38166 12980
rect 40034 12928 40040 12980
rect 40092 12968 40098 12980
rect 40770 12968 40776 12980
rect 40092 12940 40776 12968
rect 40092 12928 40098 12940
rect 40770 12928 40776 12940
rect 40828 12928 40834 12980
rect 43714 12900 43720 12912
rect 28000 12872 43720 12900
rect 28000 12841 28028 12872
rect 43714 12860 43720 12872
rect 43772 12860 43778 12912
rect 27985 12835 28043 12841
rect 27985 12832 27997 12835
rect 27632 12804 27997 12832
rect 27985 12801 27997 12804
rect 28031 12801 28043 12835
rect 27985 12795 28043 12801
rect 28258 12792 28264 12844
rect 28316 12792 28322 12844
rect 28810 12792 28816 12844
rect 28868 12832 28874 12844
rect 28905 12835 28963 12841
rect 28905 12832 28917 12835
rect 28868 12804 28917 12832
rect 28868 12792 28874 12804
rect 28905 12801 28917 12804
rect 28951 12801 28963 12835
rect 28905 12795 28963 12801
rect 28920 12764 28948 12795
rect 31570 12792 31576 12844
rect 31628 12792 31634 12844
rect 33134 12792 33140 12844
rect 33192 12792 33198 12844
rect 33229 12835 33287 12841
rect 33229 12801 33241 12835
rect 33275 12832 33287 12835
rect 34238 12832 34244 12844
rect 33275 12804 34244 12832
rect 33275 12801 33287 12804
rect 33229 12795 33287 12801
rect 34238 12792 34244 12804
rect 34296 12792 34302 12844
rect 35618 12841 35624 12844
rect 35612 12795 35624 12841
rect 35618 12792 35624 12795
rect 35676 12792 35682 12844
rect 37921 12835 37979 12841
rect 37921 12801 37933 12835
rect 37967 12832 37979 12835
rect 39850 12832 39856 12844
rect 37967 12804 39856 12832
rect 37967 12801 37979 12804
rect 37921 12795 37979 12801
rect 39850 12792 39856 12804
rect 39908 12792 39914 12844
rect 40034 12792 40040 12844
rect 40092 12832 40098 12844
rect 40681 12835 40739 12841
rect 40681 12832 40693 12835
rect 40092 12804 40693 12832
rect 40092 12792 40098 12804
rect 40681 12801 40693 12804
rect 40727 12801 40739 12835
rect 40681 12795 40739 12801
rect 40770 12792 40776 12844
rect 40828 12832 40834 12844
rect 40865 12835 40923 12841
rect 40865 12832 40877 12835
rect 40828 12804 40877 12832
rect 40828 12792 40834 12804
rect 40865 12801 40877 12804
rect 40911 12801 40923 12835
rect 40865 12795 40923 12801
rect 26252 12736 28948 12764
rect 29181 12767 29239 12773
rect 29181 12733 29193 12767
rect 29227 12733 29239 12767
rect 29181 12727 29239 12733
rect 9048 12668 9536 12696
rect 16776 12668 22508 12696
rect 22572 12668 22692 12696
rect 8754 12588 8760 12640
rect 8812 12588 8818 12640
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9398 12628 9404 12640
rect 9355 12600 9404 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9508 12628 9536 12668
rect 15286 12628 15292 12640
rect 9508 12600 15292 12628
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 16022 12588 16028 12640
rect 16080 12628 16086 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 16080 12600 16865 12628
rect 16080 12588 16086 12600
rect 16853 12597 16865 12600
rect 16899 12597 16911 12631
rect 16853 12591 16911 12597
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 22005 12631 22063 12637
rect 22005 12628 22017 12631
rect 21416 12600 22017 12628
rect 21416 12588 21422 12600
rect 22005 12597 22017 12600
rect 22051 12597 22063 12631
rect 22005 12591 22063 12597
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22572 12628 22600 12668
rect 25038 12656 25044 12708
rect 25096 12696 25102 12708
rect 26878 12696 26884 12708
rect 25096 12668 26884 12696
rect 25096 12656 25102 12668
rect 26878 12656 26884 12668
rect 26936 12656 26942 12708
rect 28810 12656 28816 12708
rect 28868 12696 28874 12708
rect 29196 12696 29224 12727
rect 31294 12724 31300 12776
rect 31352 12764 31358 12776
rect 31389 12767 31447 12773
rect 31389 12764 31401 12767
rect 31352 12736 31401 12764
rect 31352 12724 31358 12736
rect 31389 12733 31401 12736
rect 31435 12733 31447 12767
rect 31389 12727 31447 12733
rect 33413 12767 33471 12773
rect 33413 12733 33425 12767
rect 33459 12764 33471 12767
rect 34054 12764 34060 12776
rect 33459 12736 34060 12764
rect 33459 12733 33471 12736
rect 33413 12727 33471 12733
rect 34054 12724 34060 12736
rect 34112 12724 34118 12776
rect 35342 12724 35348 12776
rect 35400 12724 35406 12776
rect 37274 12724 37280 12776
rect 37332 12764 37338 12776
rect 38013 12767 38071 12773
rect 38013 12764 38025 12767
rect 37332 12736 38025 12764
rect 37332 12724 37338 12736
rect 38013 12733 38025 12736
rect 38059 12764 38071 12767
rect 38286 12764 38292 12776
rect 38059 12736 38292 12764
rect 38059 12733 38071 12736
rect 38013 12727 38071 12733
rect 38286 12724 38292 12736
rect 38344 12724 38350 12776
rect 33594 12696 33600 12708
rect 28868 12668 33600 12696
rect 28868 12656 28874 12668
rect 33594 12656 33600 12668
rect 33652 12656 33658 12708
rect 22152 12600 22600 12628
rect 22152 12588 22158 12600
rect 26786 12588 26792 12640
rect 26844 12628 26850 12640
rect 27249 12631 27307 12637
rect 27249 12628 27261 12631
rect 26844 12600 27261 12628
rect 26844 12588 26850 12600
rect 27249 12597 27261 12600
rect 27295 12597 27307 12631
rect 27249 12591 27307 12597
rect 31757 12631 31815 12637
rect 31757 12597 31769 12631
rect 31803 12628 31815 12631
rect 31846 12628 31852 12640
rect 31803 12600 31852 12628
rect 31803 12597 31815 12600
rect 31757 12591 31815 12597
rect 31846 12588 31852 12600
rect 31904 12588 31910 12640
rect 34238 12588 34244 12640
rect 34296 12628 34302 12640
rect 36722 12628 36728 12640
rect 34296 12600 36728 12628
rect 34296 12588 34302 12600
rect 36722 12588 36728 12600
rect 36780 12588 36786 12640
rect 40681 12631 40739 12637
rect 40681 12597 40693 12631
rect 40727 12628 40739 12631
rect 41414 12628 41420 12640
rect 40727 12600 41420 12628
rect 40727 12597 40739 12600
rect 40681 12591 40739 12597
rect 41414 12588 41420 12600
rect 41472 12588 41478 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 3786 12384 3792 12436
rect 3844 12424 3850 12436
rect 11885 12427 11943 12433
rect 3844 12396 10732 12424
rect 3844 12384 3850 12396
rect 7374 12316 7380 12368
rect 7432 12356 7438 12368
rect 10597 12359 10655 12365
rect 10597 12356 10609 12359
rect 7432 12328 10609 12356
rect 7432 12316 7438 12328
rect 10597 12325 10609 12328
rect 10643 12325 10655 12359
rect 10597 12319 10655 12325
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 4108 12288
rect 2832 12248 2838 12260
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1673 12223 1731 12229
rect 1673 12220 1685 12223
rect 992 12192 1685 12220
rect 992 12180 998 12192
rect 1673 12189 1685 12192
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4080 12220 4108 12260
rect 7193 12223 7251 12229
rect 4080 12192 7144 12220
rect 1026 12112 1032 12164
rect 1084 12152 1090 12164
rect 2593 12155 2651 12161
rect 2593 12152 2605 12155
rect 1084 12124 2605 12152
rect 1084 12112 1090 12124
rect 2593 12121 2605 12124
rect 2639 12121 2651 12155
rect 2593 12115 2651 12121
rect 2777 12155 2835 12161
rect 2777 12121 2789 12155
rect 2823 12152 2835 12155
rect 3878 12152 3884 12164
rect 2823 12124 3884 12152
rect 2823 12121 2835 12124
rect 2777 12115 2835 12121
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4218 12155 4276 12161
rect 4218 12152 4230 12155
rect 3988 12124 4230 12152
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 2682 12084 2688 12096
rect 1995 12056 2688 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3988 12084 4016 12124
rect 4218 12121 4230 12124
rect 4264 12121 4276 12155
rect 7116 12152 7144 12192
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7282 12220 7288 12232
rect 7239 12192 7288 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8168 12192 8493 12220
rect 8168 12180 8174 12192
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 10042 12152 10048 12164
rect 7116 12124 10048 12152
rect 4218 12115 4276 12121
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10318 12152 10324 12164
rect 10244 12124 10324 12152
rect 3476 12056 4016 12084
rect 3476 12044 3482 12056
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4982 12084 4988 12096
rect 4396 12056 4988 12084
rect 4396 12044 4402 12056
rect 4982 12044 4988 12056
rect 5040 12084 5046 12096
rect 5353 12087 5411 12093
rect 5353 12084 5365 12087
rect 5040 12056 5365 12084
rect 5040 12044 5046 12056
rect 5353 12053 5365 12056
rect 5399 12053 5411 12087
rect 5353 12047 5411 12053
rect 8297 12087 8355 12093
rect 8297 12053 8309 12087
rect 8343 12084 8355 12087
rect 10244 12084 10272 12124
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 10704 12152 10732 12396
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 11974 12424 11980 12436
rect 11931 12396 11980 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 13262 12384 13268 12436
rect 13320 12424 13326 12436
rect 13320 12396 15424 12424
rect 13320 12384 13326 12396
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 15396 12288 15424 12396
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 17405 12427 17463 12433
rect 17405 12424 17417 12427
rect 16908 12396 17417 12424
rect 16908 12384 16914 12396
rect 17405 12393 17417 12396
rect 17451 12393 17463 12427
rect 22465 12427 22523 12433
rect 17405 12387 17463 12393
rect 17512 12396 22094 12424
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 17512 12356 17540 12396
rect 15528 12328 17540 12356
rect 22066 12356 22094 12396
rect 22465 12393 22477 12427
rect 22511 12424 22523 12427
rect 22554 12424 22560 12436
rect 22511 12396 22560 12424
rect 22511 12393 22523 12396
rect 22465 12387 22523 12393
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 24578 12384 24584 12436
rect 24636 12384 24642 12436
rect 25700 12396 27844 12424
rect 25700 12356 25728 12396
rect 22066 12328 25728 12356
rect 25777 12359 25835 12365
rect 15528 12316 15534 12328
rect 25777 12325 25789 12359
rect 25823 12356 25835 12359
rect 27246 12356 27252 12368
rect 25823 12328 27252 12356
rect 25823 12325 25835 12328
rect 25777 12319 25835 12325
rect 27246 12316 27252 12328
rect 27304 12316 27310 12368
rect 27816 12356 27844 12396
rect 27890 12384 27896 12436
rect 27948 12384 27954 12436
rect 27982 12384 27988 12436
rect 28040 12424 28046 12436
rect 28997 12427 29055 12433
rect 28997 12424 29009 12427
rect 28040 12396 29009 12424
rect 28040 12384 28046 12396
rect 28997 12393 29009 12396
rect 29043 12393 29055 12427
rect 28997 12387 29055 12393
rect 31202 12384 31208 12436
rect 31260 12424 31266 12436
rect 31260 12396 35572 12424
rect 31260 12384 31266 12396
rect 35544 12356 35572 12396
rect 35618 12384 35624 12436
rect 35676 12424 35682 12436
rect 35805 12427 35863 12433
rect 35805 12424 35817 12427
rect 35676 12396 35817 12424
rect 35676 12384 35682 12396
rect 35805 12393 35817 12396
rect 35851 12393 35863 12427
rect 35805 12387 35863 12393
rect 35894 12384 35900 12436
rect 35952 12424 35958 12436
rect 36541 12427 36599 12433
rect 36541 12424 36553 12427
rect 35952 12396 36553 12424
rect 35952 12384 35958 12396
rect 36541 12393 36553 12396
rect 36587 12393 36599 12427
rect 36541 12387 36599 12393
rect 35986 12356 35992 12368
rect 27816 12328 28672 12356
rect 35544 12328 35992 12356
rect 16298 12288 16304 12300
rect 11664 12260 14412 12288
rect 15396 12260 16304 12288
rect 11664 12248 11670 12260
rect 14384 12232 14412 12260
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 16482 12248 16488 12300
rect 16540 12288 16546 12300
rect 16540 12260 17632 12288
rect 16540 12248 16546 12260
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 12066 12220 12072 12232
rect 11112 12192 12072 12220
rect 11112 12180 11118 12192
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 14182 12220 14188 12232
rect 12391 12192 14188 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14568 12192 16436 12220
rect 14568 12152 14596 12192
rect 10704 12124 14596 12152
rect 14636 12155 14694 12161
rect 14636 12121 14648 12155
rect 14682 12152 14694 12155
rect 15562 12152 15568 12164
rect 14682 12124 15568 12152
rect 14682 12121 14694 12124
rect 14636 12115 14694 12121
rect 15562 12112 15568 12124
rect 15620 12112 15626 12164
rect 16408 12152 16436 12192
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16632 12192 16681 12220
rect 16632 12180 16638 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 17604 12229 17632 12260
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 21085 12291 21143 12297
rect 21085 12288 21097 12291
rect 17828 12260 21097 12288
rect 17828 12248 17834 12260
rect 21085 12257 21097 12260
rect 21131 12257 21143 12291
rect 26326 12288 26332 12300
rect 21085 12251 21143 12257
rect 25792 12260 26332 12288
rect 21358 12229 21364 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 16816 12192 17417 12220
rect 16816 12180 16822 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12220 20131 12223
rect 20119 12192 21312 12220
rect 20119 12189 20131 12192
rect 20073 12183 20131 12189
rect 20162 12152 20168 12164
rect 16408 12124 20168 12152
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 20346 12112 20352 12164
rect 20404 12112 20410 12164
rect 21284 12152 21312 12192
rect 21352 12183 21364 12229
rect 21358 12180 21364 12183
rect 21416 12180 21422 12232
rect 23842 12180 23848 12232
rect 23900 12220 23906 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 23900 12192 24777 12220
rect 23900 12180 23906 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 21634 12152 21640 12164
rect 21284 12124 21640 12152
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 24780 12152 24808 12183
rect 24854 12180 24860 12232
rect 24912 12220 24918 12232
rect 24949 12223 25007 12229
rect 24949 12220 24961 12223
rect 24912 12192 24961 12220
rect 24912 12180 24918 12192
rect 24949 12189 24961 12192
rect 24995 12189 25007 12223
rect 24949 12183 25007 12189
rect 25038 12180 25044 12232
rect 25096 12180 25102 12232
rect 25222 12152 25228 12164
rect 24780 12124 25228 12152
rect 25222 12112 25228 12124
rect 25280 12112 25286 12164
rect 25792 12161 25820 12260
rect 26326 12248 26332 12260
rect 26384 12248 26390 12300
rect 27154 12248 27160 12300
rect 27212 12288 27218 12300
rect 27525 12291 27583 12297
rect 27525 12288 27537 12291
rect 27212 12260 27537 12288
rect 27212 12248 27218 12260
rect 27525 12257 27537 12260
rect 27571 12288 27583 12291
rect 28644 12288 28672 12328
rect 35986 12316 35992 12328
rect 36044 12316 36050 12368
rect 38102 12356 38108 12368
rect 37016 12328 38108 12356
rect 31202 12288 31208 12300
rect 27571 12260 28488 12288
rect 28644 12260 31208 12288
rect 27571 12257 27583 12260
rect 27525 12251 27583 12257
rect 28460 12232 28488 12260
rect 31202 12248 31208 12260
rect 31260 12248 31266 12300
rect 37016 12297 37044 12328
rect 38102 12316 38108 12328
rect 38160 12316 38166 12368
rect 39209 12359 39267 12365
rect 39209 12325 39221 12359
rect 39255 12325 39267 12359
rect 39209 12319 39267 12325
rect 37001 12291 37059 12297
rect 37001 12288 37013 12291
rect 35365 12260 37013 12288
rect 26053 12223 26111 12229
rect 26053 12189 26065 12223
rect 26099 12220 26111 12223
rect 26513 12223 26571 12229
rect 26513 12220 26525 12223
rect 26099 12192 26525 12220
rect 26099 12189 26111 12192
rect 26053 12183 26111 12189
rect 26513 12189 26525 12192
rect 26559 12189 26571 12223
rect 26513 12183 26571 12189
rect 26694 12180 26700 12232
rect 26752 12180 26758 12232
rect 26786 12180 26792 12232
rect 26844 12180 26850 12232
rect 26970 12180 26976 12232
rect 27028 12180 27034 12232
rect 27065 12223 27123 12229
rect 27065 12189 27077 12223
rect 27111 12189 27123 12223
rect 27065 12183 27123 12189
rect 25777 12155 25835 12161
rect 25777 12121 25789 12155
rect 25823 12121 25835 12155
rect 27080 12152 27108 12183
rect 27338 12180 27344 12232
rect 27396 12220 27402 12232
rect 27709 12223 27767 12229
rect 27709 12220 27721 12223
rect 27396 12192 27721 12220
rect 27396 12180 27402 12192
rect 27709 12189 27721 12192
rect 27755 12189 27767 12223
rect 27709 12183 27767 12189
rect 28350 12180 28356 12232
rect 28408 12180 28414 12232
rect 28442 12180 28448 12232
rect 28500 12180 28506 12232
rect 28810 12180 28816 12232
rect 28868 12229 28874 12232
rect 28868 12220 28876 12229
rect 28868 12192 28913 12220
rect 28868 12183 28876 12192
rect 28868 12180 28874 12183
rect 31754 12180 31760 12232
rect 31812 12180 31818 12232
rect 31846 12180 31852 12232
rect 31904 12220 31910 12232
rect 32013 12223 32071 12229
rect 32013 12220 32025 12223
rect 31904 12192 32025 12220
rect 31904 12180 31910 12192
rect 32013 12189 32025 12192
rect 32059 12189 32071 12223
rect 32013 12183 32071 12189
rect 32490 12180 32496 12232
rect 32548 12220 32554 12232
rect 35365 12220 35393 12260
rect 37001 12257 37013 12260
rect 37047 12257 37059 12291
rect 37001 12251 37059 12257
rect 37182 12248 37188 12300
rect 37240 12248 37246 12300
rect 38746 12248 38752 12300
rect 38804 12288 38810 12300
rect 39224 12288 39252 12319
rect 44082 12316 44088 12368
rect 44140 12356 44146 12368
rect 47946 12356 47952 12368
rect 44140 12328 47952 12356
rect 44140 12316 44146 12328
rect 47946 12316 47952 12328
rect 48004 12316 48010 12368
rect 38804 12260 39160 12288
rect 39224 12260 40264 12288
rect 38804 12248 38810 12260
rect 32548 12192 35393 12220
rect 35437 12223 35495 12229
rect 32548 12180 32554 12192
rect 35437 12189 35449 12223
rect 35483 12189 35495 12223
rect 35437 12183 35495 12189
rect 35621 12223 35679 12229
rect 35621 12189 35633 12223
rect 35667 12220 35679 12223
rect 36262 12220 36268 12232
rect 35667 12192 36268 12220
rect 35667 12189 35679 12192
rect 35621 12183 35679 12189
rect 28534 12152 28540 12164
rect 25777 12115 25835 12121
rect 25884 12124 26096 12152
rect 27080 12124 28540 12152
rect 8343 12056 10272 12084
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 10781 12087 10839 12093
rect 10781 12084 10793 12087
rect 10744 12056 10793 12084
rect 10744 12044 10750 12056
rect 10781 12053 10793 12056
rect 10827 12053 10839 12087
rect 10781 12047 10839 12053
rect 12253 12087 12311 12093
rect 12253 12053 12265 12087
rect 12299 12084 12311 12087
rect 12342 12084 12348 12096
rect 12299 12056 12348 12084
rect 12299 12053 12311 12056
rect 12253 12047 12311 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 15436 12056 15761 12084
rect 15436 12044 15442 12056
rect 15749 12053 15761 12056
rect 15795 12084 15807 12087
rect 16482 12084 16488 12096
rect 15795 12056 16488 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 16577 12087 16635 12093
rect 16577 12053 16589 12087
rect 16623 12084 16635 12087
rect 16666 12084 16672 12096
rect 16623 12056 16672 12084
rect 16623 12053 16635 12056
rect 16577 12047 16635 12053
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 18414 12084 18420 12096
rect 16899 12056 18420 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 25884 12084 25912 12124
rect 19116 12056 25912 12084
rect 19116 12044 19122 12056
rect 25958 12044 25964 12096
rect 26016 12044 26022 12096
rect 26068 12084 26096 12124
rect 28534 12112 28540 12124
rect 28592 12112 28598 12164
rect 28626 12112 28632 12164
rect 28684 12112 28690 12164
rect 28718 12112 28724 12164
rect 28776 12112 28782 12164
rect 28902 12112 28908 12164
rect 28960 12152 28966 12164
rect 28960 12124 30144 12152
rect 28960 12112 28966 12124
rect 30006 12084 30012 12096
rect 26068 12056 30012 12084
rect 30006 12044 30012 12056
rect 30064 12044 30070 12096
rect 30116 12084 30144 12124
rect 30650 12112 30656 12164
rect 30708 12152 30714 12164
rect 35452 12152 35480 12183
rect 36262 12180 36268 12192
rect 36320 12180 36326 12232
rect 36722 12180 36728 12232
rect 36780 12220 36786 12232
rect 36909 12223 36967 12229
rect 36909 12220 36921 12223
rect 36780 12192 36921 12220
rect 36780 12180 36786 12192
rect 36909 12189 36921 12192
rect 36955 12189 36967 12223
rect 38654 12220 38660 12232
rect 36909 12183 36967 12189
rect 37108 12192 38660 12220
rect 30708 12124 35480 12152
rect 30708 12112 30714 12124
rect 35526 12112 35532 12164
rect 35584 12152 35590 12164
rect 37108 12152 37136 12192
rect 38654 12180 38660 12192
rect 38712 12180 38718 12232
rect 39022 12180 39028 12232
rect 39080 12180 39086 12232
rect 39132 12220 39160 12260
rect 39206 12220 39212 12232
rect 39132 12192 39212 12220
rect 39206 12180 39212 12192
rect 39264 12220 39270 12232
rect 40236 12229 40264 12260
rect 40037 12223 40095 12229
rect 40037 12220 40049 12223
rect 39264 12192 40049 12220
rect 39264 12180 39270 12192
rect 40037 12189 40049 12192
rect 40083 12189 40095 12223
rect 40037 12183 40095 12189
rect 40221 12223 40279 12229
rect 40221 12189 40233 12223
rect 40267 12189 40279 12223
rect 40221 12183 40279 12189
rect 35584 12124 37136 12152
rect 38841 12155 38899 12161
rect 35584 12112 35590 12124
rect 38841 12121 38853 12155
rect 38887 12121 38899 12155
rect 38841 12115 38899 12121
rect 33134 12084 33140 12096
rect 30116 12056 33140 12084
rect 33134 12044 33140 12056
rect 33192 12044 33198 12096
rect 38856 12084 38884 12115
rect 38930 12112 38936 12164
rect 38988 12112 38994 12164
rect 40052 12152 40080 12183
rect 41322 12180 41328 12232
rect 41380 12180 41386 12232
rect 41414 12180 41420 12232
rect 41472 12220 41478 12232
rect 41581 12223 41639 12229
rect 41581 12220 41593 12223
rect 41472 12192 41593 12220
rect 41472 12180 41478 12192
rect 41581 12189 41593 12192
rect 41627 12189 41639 12223
rect 41581 12183 41639 12189
rect 42334 12152 42340 12164
rect 40052 12124 42340 12152
rect 42334 12112 42340 12124
rect 42392 12112 42398 12164
rect 40218 12084 40224 12096
rect 38856 12056 40224 12084
rect 40218 12044 40224 12056
rect 40276 12044 40282 12096
rect 40402 12044 40408 12096
rect 40460 12044 40466 12096
rect 42426 12044 42432 12096
rect 42484 12084 42490 12096
rect 42705 12087 42763 12093
rect 42705 12084 42717 12087
rect 42484 12056 42717 12084
rect 42484 12044 42490 12056
rect 42705 12053 42717 12056
rect 42751 12053 42763 12087
rect 42705 12047 42763 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 3418 11840 3424 11892
rect 3476 11840 3482 11892
rect 3878 11840 3884 11892
rect 3936 11840 3942 11892
rect 4816 11852 7236 11880
rect 1118 11772 1124 11824
rect 1176 11812 1182 11824
rect 2593 11815 2651 11821
rect 2593 11812 2605 11815
rect 1176 11784 2605 11812
rect 1176 11772 1182 11784
rect 2593 11781 2605 11784
rect 2639 11781 2651 11815
rect 2593 11775 2651 11781
rect 2774 11772 2780 11824
rect 2832 11772 2838 11824
rect 3050 11772 3056 11824
rect 3108 11812 3114 11824
rect 4816 11812 4844 11852
rect 5350 11812 5356 11824
rect 3108 11784 4844 11812
rect 4908 11784 5356 11812
rect 3108 11772 3114 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 3694 11744 3700 11756
rect 1627 11716 3700 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 4246 11744 4252 11756
rect 3835 11716 4252 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4908 11753 4936 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 7208 11753 7236 11852
rect 7282 11840 7288 11892
rect 7340 11840 7346 11892
rect 10226 11840 10232 11892
rect 10284 11840 10290 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 15470 11880 15476 11892
rect 12124 11852 15476 11880
rect 12124 11840 12130 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15562 11840 15568 11892
rect 15620 11840 15626 11892
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 17053 11883 17111 11889
rect 17053 11880 17065 11883
rect 16632 11852 17065 11880
rect 16632 11840 16638 11852
rect 17053 11849 17065 11852
rect 17099 11849 17111 11883
rect 17053 11843 17111 11849
rect 17218 11840 17224 11892
rect 17276 11840 17282 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17770 11880 17776 11892
rect 17552 11852 17776 11880
rect 17552 11840 17558 11852
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 20346 11880 20352 11892
rect 18196 11852 20352 11880
rect 18196 11840 18202 11852
rect 8754 11812 8760 11824
rect 8128 11784 8760 11812
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4356 11716 4905 11744
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1765 11679 1823 11685
rect 1765 11676 1777 11679
rect 992 11648 1777 11676
rect 992 11636 998 11648
rect 1765 11645 1777 11648
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 3973 11679 4031 11685
rect 2556 11648 3372 11676
rect 2556 11636 2562 11648
rect 3344 11608 3372 11648
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 3988 11608 4016 11639
rect 3344 11580 4016 11608
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 4356 11540 4384 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 8018 11744 8024 11756
rect 7239 11716 8024 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 5092 11676 5120 11707
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8128 11753 8156 11784
rect 8754 11772 8760 11784
rect 8812 11772 8818 11824
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 15933 11815 15991 11821
rect 15933 11812 15945 11815
rect 14240 11784 15945 11812
rect 14240 11772 14246 11784
rect 15933 11781 15945 11784
rect 15979 11812 15991 11815
rect 15979 11784 16436 11812
rect 15979 11781 15991 11784
rect 15933 11775 15991 11781
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11744 9919 11747
rect 10502 11744 10508 11756
rect 9907 11716 10508 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 7374 11676 7380 11688
rect 5092 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 9876 11676 9904 11707
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 16022 11704 16028 11756
rect 16080 11704 16086 11756
rect 16408 11744 16436 11784
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 16853 11815 16911 11821
rect 16853 11812 16865 11815
rect 16540 11784 16865 11812
rect 16540 11772 16546 11784
rect 16853 11781 16865 11784
rect 16899 11781 16911 11815
rect 16853 11775 16911 11781
rect 16758 11744 16764 11756
rect 16408 11716 16764 11744
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 17236 11744 17264 11840
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17236 11716 17693 11744
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17862 11704 17868 11756
rect 17920 11704 17926 11756
rect 20088 11753 20116 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 21634 11880 21640 11892
rect 20680 11852 21640 11880
rect 20680 11840 20686 11852
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 22189 11883 22247 11889
rect 22189 11849 22201 11883
rect 22235 11880 22247 11883
rect 22278 11880 22284 11892
rect 22235 11852 22284 11880
rect 22235 11849 22247 11852
rect 22189 11843 22247 11849
rect 22278 11840 22284 11852
rect 22336 11880 22342 11892
rect 25958 11880 25964 11892
rect 22336 11852 25964 11880
rect 22336 11840 22342 11852
rect 25958 11840 25964 11852
rect 26016 11840 26022 11892
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 28537 11883 28595 11889
rect 28537 11880 28549 11883
rect 28500 11852 28549 11880
rect 28500 11840 28506 11852
rect 28537 11849 28549 11852
rect 28583 11849 28595 11883
rect 28537 11843 28595 11849
rect 29362 11840 29368 11892
rect 29420 11880 29426 11892
rect 29917 11883 29975 11889
rect 29917 11880 29929 11883
rect 29420 11852 29929 11880
rect 29420 11840 29426 11852
rect 29917 11849 29929 11852
rect 29963 11849 29975 11883
rect 29917 11843 29975 11849
rect 30006 11840 30012 11892
rect 30064 11880 30070 11892
rect 30064 11852 39988 11880
rect 30064 11840 30070 11852
rect 20162 11772 20168 11824
rect 20220 11772 20226 11824
rect 24486 11812 24492 11824
rect 20272 11784 24492 11812
rect 20272 11753 20300 11784
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 25590 11772 25596 11824
rect 25648 11812 25654 11824
rect 30282 11812 30288 11824
rect 25648 11784 25912 11812
rect 25648 11772 25654 11784
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11713 20315 11747
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 20257 11707 20315 11713
rect 21468 11716 22017 11744
rect 7892 11648 9904 11676
rect 7892 11636 7898 11648
rect 9950 11636 9956 11688
rect 10008 11636 10014 11688
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 20272 11676 20300 11707
rect 14240 11648 20300 11676
rect 20717 11679 20775 11685
rect 14240 11636 14246 11648
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 21358 11676 21364 11688
rect 20763 11648 21364 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 5261 11611 5319 11617
rect 5261 11577 5273 11611
rect 5307 11608 5319 11611
rect 5534 11608 5540 11620
rect 5307 11580 5540 11608
rect 5307 11577 5319 11580
rect 5261 11571 5319 11577
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 20990 11608 20996 11620
rect 10376 11580 20996 11608
rect 10376 11568 10382 11580
rect 20990 11568 20996 11580
rect 21048 11568 21054 11620
rect 21468 11608 21496 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 25884 11753 25912 11784
rect 27172 11784 30288 11812
rect 25869 11747 25927 11753
rect 25869 11713 25881 11747
rect 25915 11713 25927 11747
rect 25869 11707 25927 11713
rect 27172 11688 27200 11784
rect 30282 11772 30288 11784
rect 30340 11772 30346 11824
rect 39022 11772 39028 11824
rect 39080 11812 39086 11824
rect 39761 11815 39819 11821
rect 39761 11812 39773 11815
rect 39080 11784 39773 11812
rect 39080 11772 39086 11784
rect 39761 11781 39773 11784
rect 39807 11781 39819 11815
rect 39761 11775 39819 11781
rect 39850 11772 39856 11824
rect 39908 11772 39914 11824
rect 39960 11812 39988 11852
rect 40126 11840 40132 11892
rect 40184 11840 40190 11892
rect 55950 11812 55956 11824
rect 39960 11784 55956 11812
rect 55950 11772 55956 11784
rect 56008 11772 56014 11824
rect 27246 11704 27252 11756
rect 27304 11744 27310 11756
rect 27413 11747 27471 11753
rect 27413 11744 27425 11747
rect 27304 11716 27425 11744
rect 27304 11704 27310 11716
rect 27413 11713 27425 11716
rect 27459 11713 27471 11747
rect 27413 11707 27471 11713
rect 28534 11704 28540 11756
rect 28592 11744 28598 11756
rect 28994 11744 29000 11756
rect 28592 11716 29000 11744
rect 28592 11704 28598 11716
rect 28994 11704 29000 11716
rect 29052 11744 29058 11756
rect 29454 11744 29460 11756
rect 29052 11716 29460 11744
rect 29052 11704 29058 11716
rect 29454 11704 29460 11716
rect 29512 11704 29518 11756
rect 29730 11704 29736 11756
rect 29788 11704 29794 11756
rect 30009 11747 30067 11753
rect 30009 11713 30021 11747
rect 30055 11744 30067 11747
rect 32858 11744 32864 11756
rect 30055 11716 32864 11744
rect 30055 11713 30067 11716
rect 30009 11707 30067 11713
rect 32858 11704 32864 11716
rect 32916 11704 32922 11756
rect 33318 11704 33324 11756
rect 33376 11744 33382 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 33376 11716 37841 11744
rect 33376 11704 33382 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 38562 11704 38568 11756
rect 38620 11704 38626 11756
rect 38749 11747 38807 11753
rect 38749 11713 38761 11747
rect 38795 11713 38807 11747
rect 38749 11707 38807 11713
rect 21634 11636 21640 11688
rect 21692 11676 21698 11688
rect 25501 11679 25559 11685
rect 25501 11676 25513 11679
rect 21692 11648 25513 11676
rect 21692 11636 21698 11648
rect 25501 11645 25513 11648
rect 25547 11645 25559 11679
rect 25501 11639 25559 11645
rect 25682 11636 25688 11688
rect 25740 11636 25746 11688
rect 25777 11679 25835 11685
rect 25777 11645 25789 11679
rect 25823 11676 25835 11679
rect 25823 11648 25912 11676
rect 25823 11645 25835 11648
rect 25777 11639 25835 11645
rect 21100 11580 21496 11608
rect 2280 11512 4384 11540
rect 2280 11500 2286 11512
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8110 11540 8116 11552
rect 7524 11512 8116 11540
rect 7524 11500 7530 11512
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9548 11512 9873 11540
rect 9548 11500 9554 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 9861 11503 9919 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 17037 11543 17095 11549
rect 17037 11540 17049 11543
rect 16724 11512 17049 11540
rect 16724 11500 16730 11512
rect 17037 11509 17049 11512
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 17681 11543 17739 11549
rect 17681 11509 17693 11543
rect 17727 11540 17739 11543
rect 18598 11540 18604 11552
rect 17727 11512 18604 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 21100 11540 21128 11580
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 25590 11608 25596 11620
rect 21600 11580 25596 11608
rect 21600 11568 21606 11580
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 20036 11512 21128 11540
rect 25884 11540 25912 11648
rect 25958 11636 25964 11688
rect 26016 11636 26022 11688
rect 27154 11636 27160 11688
rect 27212 11636 27218 11688
rect 30374 11636 30380 11688
rect 30432 11676 30438 11688
rect 38764 11676 38792 11707
rect 38838 11704 38844 11756
rect 38896 11704 38902 11756
rect 39577 11747 39635 11753
rect 39577 11713 39589 11747
rect 39623 11713 39635 11747
rect 39577 11707 39635 11713
rect 30432 11648 38792 11676
rect 30432 11636 30438 11648
rect 39114 11636 39120 11688
rect 39172 11676 39178 11688
rect 39592 11676 39620 11707
rect 39942 11704 39948 11756
rect 40000 11704 40006 11756
rect 42426 11676 42432 11688
rect 39172 11648 42432 11676
rect 39172 11636 39178 11648
rect 42426 11636 42432 11648
rect 42484 11636 42490 11688
rect 38565 11611 38623 11617
rect 38565 11577 38577 11611
rect 38611 11608 38623 11611
rect 40034 11608 40040 11620
rect 38611 11580 40040 11608
rect 38611 11577 38623 11580
rect 38565 11571 38623 11577
rect 40034 11568 40040 11580
rect 40092 11568 40098 11620
rect 28074 11540 28080 11552
rect 25884 11512 28080 11540
rect 20036 11500 20042 11512
rect 28074 11500 28080 11512
rect 28132 11500 28138 11552
rect 29733 11543 29791 11549
rect 29733 11509 29745 11543
rect 29779 11540 29791 11543
rect 31478 11540 31484 11552
rect 29779 11512 31484 11540
rect 29779 11509 29791 11512
rect 29733 11503 29791 11509
rect 31478 11500 31484 11512
rect 31536 11500 31542 11552
rect 37918 11500 37924 11552
rect 37976 11540 37982 11552
rect 38013 11543 38071 11549
rect 38013 11540 38025 11543
rect 37976 11512 38025 11540
rect 37976 11500 37982 11512
rect 38013 11509 38025 11512
rect 38059 11509 38071 11543
rect 38013 11503 38071 11509
rect 38654 11500 38660 11552
rect 38712 11540 38718 11552
rect 43254 11540 43260 11552
rect 38712 11512 43260 11540
rect 38712 11500 38718 11512
rect 43254 11500 43260 11512
rect 43312 11500 43318 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 4982 11296 4988 11348
rect 5040 11296 5046 11348
rect 5258 11296 5264 11348
rect 5316 11296 5322 11348
rect 8294 11336 8300 11348
rect 7852 11308 8300 11336
rect 3050 11228 3056 11280
rect 3108 11228 3114 11280
rect 3694 11228 3700 11280
rect 3752 11268 3758 11280
rect 6454 11268 6460 11280
rect 3752 11240 6460 11268
rect 3752 11228 3758 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 3936 11172 4997 11200
rect 3936 11160 3942 11172
rect 4985 11169 4997 11172
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 7852 11209 7880 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 12989 11339 13047 11345
rect 12989 11336 13001 11339
rect 12952 11308 13001 11336
rect 12952 11296 12958 11308
rect 12989 11305 13001 11308
rect 13035 11305 13047 11339
rect 12989 11299 13047 11305
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 17862 11336 17868 11348
rect 16356 11308 17868 11336
rect 16356 11296 16362 11308
rect 17862 11296 17868 11308
rect 17920 11336 17926 11348
rect 19334 11336 19340 11348
rect 17920 11308 19340 11336
rect 17920 11296 17926 11308
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 21358 11296 21364 11348
rect 21416 11336 21422 11348
rect 23658 11336 23664 11348
rect 21416 11308 23664 11336
rect 21416 11296 21422 11308
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 27706 11296 27712 11348
rect 27764 11336 27770 11348
rect 28626 11336 28632 11348
rect 27764 11308 28632 11336
rect 27764 11296 27770 11308
rect 28626 11296 28632 11308
rect 28684 11296 28690 11348
rect 29730 11296 29736 11348
rect 29788 11336 29794 11348
rect 30377 11339 30435 11345
rect 30377 11336 30389 11339
rect 29788 11308 30389 11336
rect 29788 11296 29794 11308
rect 30377 11305 30389 11308
rect 30423 11305 30435 11339
rect 30377 11299 30435 11305
rect 38562 11296 38568 11348
rect 38620 11336 38626 11348
rect 39393 11339 39451 11345
rect 39393 11336 39405 11339
rect 38620 11308 39405 11336
rect 38620 11296 38626 11308
rect 39393 11305 39405 11308
rect 39439 11305 39451 11339
rect 39393 11299 39451 11305
rect 8386 11268 8392 11280
rect 8220 11240 8392 11268
rect 8220 11209 8248 11240
rect 8386 11228 8392 11240
rect 8444 11268 8450 11280
rect 8444 11240 9076 11268
rect 8444 11228 8450 11240
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 5408 11172 7849 11200
rect 5408 11160 5414 11172
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11200 8355 11203
rect 8754 11200 8760 11212
rect 8343 11172 8760 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9048 11200 9076 11240
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 10321 11271 10379 11277
rect 10321 11268 10333 11271
rect 10192 11240 10333 11268
rect 10192 11228 10198 11240
rect 10321 11237 10333 11240
rect 10367 11237 10379 11271
rect 10321 11231 10379 11237
rect 9490 11200 9496 11212
rect 9048 11172 9496 11200
rect 9490 11160 9496 11172
rect 9548 11200 9554 11212
rect 10336 11200 10364 11231
rect 24670 11228 24676 11280
rect 24728 11268 24734 11280
rect 32585 11271 32643 11277
rect 24728 11240 31754 11268
rect 24728 11228 24734 11240
rect 10962 11200 10968 11212
rect 9548 11172 10088 11200
rect 10336 11172 10968 11200
rect 9548 11160 9554 11172
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 3970 11132 3976 11144
rect 1719 11104 3976 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7282 11132 7288 11144
rect 7147 11104 7288 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7926 11132 7932 11144
rect 7392 11104 7932 11132
rect 1946 11073 1952 11076
rect 1940 11027 1952 11073
rect 1946 11024 1952 11027
rect 2004 11024 2010 11076
rect 4908 11064 4936 11092
rect 5258 11064 5264 11076
rect 4908 11036 5264 11064
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 6932 11064 6960 11092
rect 7392 11064 7420 11104
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 8076 11104 8401 11132
rect 8076 11092 8082 11104
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 9950 11132 9956 11144
rect 9723 11104 9956 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 6932 11036 7420 11064
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 9692 11064 9720 11095
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10060 11141 10088 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 15841 11203 15899 11209
rect 15841 11200 15853 11203
rect 13872 11172 15853 11200
rect 13872 11160 13878 11172
rect 15841 11169 15853 11172
rect 15887 11169 15899 11203
rect 15841 11163 15899 11169
rect 16025 11203 16083 11209
rect 16025 11169 16037 11203
rect 16071 11200 16083 11203
rect 16574 11200 16580 11212
rect 16071 11172 16580 11200
rect 16071 11169 16083 11172
rect 16025 11163 16083 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 22373 11203 22431 11209
rect 22373 11200 22385 11203
rect 21652 11172 22385 11200
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 10502 11132 10508 11144
rect 10459 11104 10508 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 14182 11132 14188 11144
rect 11716 11104 14188 11132
rect 7616 11036 9720 11064
rect 7616 11024 7622 11036
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 11716 11064 11744 11104
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 15102 11132 15108 11144
rect 14516 11104 15108 11132
rect 14516 11092 14522 11104
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 9916 11036 11744 11064
rect 11876 11067 11934 11073
rect 9916 11024 9922 11036
rect 11876 11033 11888 11067
rect 11922 11064 11934 11067
rect 12250 11064 12256 11076
rect 11922 11036 12256 11064
rect 11922 11033 11934 11036
rect 11876 11027 11934 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15197 11067 15255 11073
rect 15197 11064 15209 11067
rect 15068 11036 15209 11064
rect 15068 11024 15074 11036
rect 15197 11033 15209 11036
rect 15243 11033 15255 11067
rect 16132 11064 16160 11095
rect 16206 11092 16212 11144
rect 16264 11092 16270 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 17126 11132 17132 11144
rect 16347 11104 17132 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18598 11092 18604 11144
rect 18656 11092 18662 11144
rect 21358 11092 21364 11144
rect 21416 11092 21422 11144
rect 21652 11141 21680 11172
rect 22373 11169 22385 11172
rect 22419 11200 22431 11203
rect 22419 11172 25084 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 25056 11144 25084 11172
rect 30006 11160 30012 11212
rect 30064 11200 30070 11212
rect 31726 11200 31754 11240
rect 32585 11237 32597 11271
rect 32631 11268 32643 11271
rect 33962 11268 33968 11280
rect 32631 11240 33968 11268
rect 32631 11237 32643 11240
rect 32585 11231 32643 11237
rect 33962 11228 33968 11240
rect 34020 11228 34026 11280
rect 38930 11268 38936 11280
rect 35360 11240 38936 11268
rect 35360 11200 35388 11240
rect 38930 11228 38936 11240
rect 38988 11228 38994 11280
rect 42705 11271 42763 11277
rect 42705 11237 42717 11271
rect 42751 11268 42763 11271
rect 42751 11240 43392 11268
rect 42751 11237 42763 11240
rect 42705 11231 42763 11237
rect 30064 11172 30236 11200
rect 31726 11172 35388 11200
rect 30064 11160 30070 11172
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 18046 11064 18052 11076
rect 16132 11036 18052 11064
rect 15197 11027 15255 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 21545 11067 21603 11073
rect 21545 11033 21557 11067
rect 21591 11064 21603 11067
rect 22278 11064 22284 11076
rect 21591 11036 22284 11064
rect 21591 11033 21603 11036
rect 21545 11027 21603 11033
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 24964 11064 24992 11095
rect 25038 11092 25044 11144
rect 25096 11132 25102 11144
rect 25225 11135 25283 11141
rect 25225 11132 25237 11135
rect 25096 11104 25237 11132
rect 25096 11092 25102 11104
rect 25225 11101 25237 11104
rect 25271 11132 25283 11135
rect 26602 11132 26608 11144
rect 25271 11104 26608 11132
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 28258 11092 28264 11144
rect 28316 11132 28322 11144
rect 28902 11132 28908 11144
rect 28316 11104 28908 11132
rect 28316 11092 28322 11104
rect 28902 11092 28908 11104
rect 28960 11132 28966 11144
rect 30208 11141 30236 11172
rect 38010 11160 38016 11212
rect 38068 11200 38074 11212
rect 38105 11203 38163 11209
rect 38105 11200 38117 11203
rect 38068 11172 38117 11200
rect 38068 11160 38074 11172
rect 38105 11169 38117 11172
rect 38151 11169 38163 11203
rect 38105 11163 38163 11169
rect 38856 11172 41460 11200
rect 29825 11135 29883 11141
rect 29825 11132 29837 11135
rect 28960 11104 29837 11132
rect 28960 11092 28966 11104
rect 29825 11101 29837 11104
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 30193 11135 30251 11141
rect 30193 11101 30205 11135
rect 30239 11101 30251 11135
rect 30193 11095 30251 11101
rect 32766 11092 32772 11144
rect 32824 11092 32830 11144
rect 32858 11092 32864 11144
rect 32916 11092 32922 11144
rect 37642 11092 37648 11144
rect 37700 11092 37706 11144
rect 37829 11135 37887 11141
rect 37829 11101 37841 11135
rect 37875 11132 37887 11135
rect 38746 11132 38752 11144
rect 37875 11104 38752 11132
rect 37875 11101 37887 11104
rect 37829 11095 37887 11101
rect 38746 11092 38752 11104
rect 38804 11092 38810 11144
rect 38856 11141 38884 11172
rect 38841 11135 38899 11141
rect 38841 11101 38853 11135
rect 38887 11101 38899 11135
rect 38841 11095 38899 11101
rect 39114 11092 39120 11144
rect 39172 11092 39178 11144
rect 39209 11135 39267 11141
rect 39209 11101 39221 11135
rect 39255 11132 39267 11135
rect 39298 11132 39304 11144
rect 39255 11104 39304 11132
rect 39255 11101 39267 11104
rect 39209 11095 39267 11101
rect 39298 11092 39304 11104
rect 39356 11132 39362 11144
rect 39942 11132 39948 11144
rect 39356 11104 39948 11132
rect 39356 11092 39362 11104
rect 39942 11092 39948 11104
rect 40000 11092 40006 11144
rect 40678 11092 40684 11144
rect 40736 11132 40742 11144
rect 41322 11132 41328 11144
rect 40736 11104 41328 11132
rect 40736 11092 40742 11104
rect 41322 11092 41328 11104
rect 41380 11092 41386 11144
rect 41432 11132 41460 11172
rect 42720 11132 42748 11231
rect 43364 11144 43392 11240
rect 44266 11160 44272 11212
rect 44324 11160 44330 11212
rect 41432 11104 42748 11132
rect 43346 11092 43352 11144
rect 43404 11132 43410 11144
rect 44085 11135 44143 11141
rect 44085 11132 44097 11135
rect 43404 11104 44097 11132
rect 43404 11092 43410 11104
rect 44085 11101 44097 11104
rect 44131 11101 44143 11135
rect 44085 11095 44143 11101
rect 25314 11064 25320 11076
rect 24964 11036 25320 11064
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 29914 11024 29920 11076
rect 29972 11064 29978 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 29972 11036 30021 11064
rect 29972 11024 29978 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 30101 11067 30159 11073
rect 30101 11033 30113 11067
rect 30147 11033 30159 11067
rect 30101 11027 30159 11033
rect 7009 10999 7067 11005
rect 7009 10965 7021 10999
rect 7055 10996 7067 10999
rect 7374 10996 7380 11008
rect 7055 10968 7380 10996
rect 7055 10965 7067 10968
rect 7009 10959 7067 10965
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 17954 10996 17960 11008
rect 9824 10968 17960 10996
rect 9824 10956 9830 10968
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 18509 10999 18567 11005
rect 18509 10965 18521 10999
rect 18555 10996 18567 10999
rect 18874 10996 18880 11008
rect 18555 10968 18880 10996
rect 18555 10965 18567 10968
rect 18509 10959 18567 10965
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 21177 10999 21235 11005
rect 21177 10965 21189 10999
rect 21223 10996 21235 10999
rect 21266 10996 21272 11008
rect 21223 10968 21272 10996
rect 21223 10965 21235 10968
rect 21177 10959 21235 10965
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 24762 10956 24768 11008
rect 24820 10956 24826 11008
rect 25130 10956 25136 11008
rect 25188 10956 25194 11008
rect 29638 10956 29644 11008
rect 29696 10996 29702 11008
rect 30116 10996 30144 11027
rect 32582 11024 32588 11076
rect 32640 11024 32646 11076
rect 33226 11024 33232 11076
rect 33284 11064 33290 11076
rect 35434 11064 35440 11076
rect 33284 11036 35440 11064
rect 33284 11024 33290 11036
rect 35434 11024 35440 11036
rect 35492 11024 35498 11076
rect 35526 11024 35532 11076
rect 35584 11064 35590 11076
rect 37737 11067 37795 11073
rect 37737 11064 37749 11067
rect 35584 11036 37749 11064
rect 35584 11024 35590 11036
rect 37737 11033 37749 11036
rect 37783 11033 37795 11067
rect 37737 11027 37795 11033
rect 37918 11024 37924 11076
rect 37976 11073 37982 11076
rect 37976 11067 38005 11073
rect 37993 11064 38005 11067
rect 38102 11064 38108 11076
rect 37993 11036 38108 11064
rect 37993 11033 38005 11036
rect 37976 11027 38005 11033
rect 37976 11024 37982 11027
rect 38102 11024 38108 11036
rect 38160 11024 38166 11076
rect 38470 11024 38476 11076
rect 38528 11064 38534 11076
rect 38930 11064 38936 11076
rect 38528 11036 38936 11064
rect 38528 11024 38534 11036
rect 38930 11024 38936 11036
rect 38988 11024 38994 11076
rect 39022 11024 39028 11076
rect 39080 11024 39086 11076
rect 41592 11067 41650 11073
rect 41592 11033 41604 11067
rect 41638 11064 41650 11067
rect 42978 11064 42984 11076
rect 41638 11036 42984 11064
rect 41638 11033 41650 11036
rect 41592 11027 41650 11033
rect 42978 11024 42984 11036
rect 43036 11024 43042 11076
rect 43530 11024 43536 11076
rect 43588 11064 43594 11076
rect 44177 11067 44235 11073
rect 44177 11064 44189 11067
rect 43588 11036 44189 11064
rect 43588 11024 43594 11036
rect 44177 11033 44189 11036
rect 44223 11033 44235 11067
rect 44177 11027 44235 11033
rect 29696 10968 30144 10996
rect 29696 10956 29702 10968
rect 31018 10956 31024 11008
rect 31076 10996 31082 11008
rect 36722 10996 36728 11008
rect 31076 10968 36728 10996
rect 31076 10956 31082 10968
rect 36722 10956 36728 10968
rect 36780 10956 36786 11008
rect 37458 10956 37464 11008
rect 37516 10956 37522 11008
rect 43162 10956 43168 11008
rect 43220 10996 43226 11008
rect 43717 10999 43775 11005
rect 43717 10996 43729 10999
rect 43220 10968 43729 10996
rect 43220 10956 43226 10968
rect 43717 10965 43729 10968
rect 43763 10965 43775 10999
rect 43717 10959 43775 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1946 10752 1952 10804
rect 2004 10752 2010 10804
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 3050 10792 3056 10804
rect 2363 10764 3056 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 5994 10792 6000 10804
rect 5828 10764 6000 10792
rect 2409 10727 2467 10733
rect 2409 10693 2421 10727
rect 2455 10724 2467 10727
rect 2498 10724 2504 10736
rect 2455 10696 2504 10724
rect 2455 10693 2467 10696
rect 2409 10687 2467 10693
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 5828 10733 5856 10764
rect 5994 10752 6000 10764
rect 6052 10792 6058 10804
rect 9766 10792 9772 10804
rect 6052 10764 9772 10792
rect 6052 10752 6058 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 12250 10752 12256 10804
rect 12308 10752 12314 10804
rect 12621 10795 12679 10801
rect 12621 10761 12633 10795
rect 12667 10792 12679 10795
rect 12894 10792 12900 10804
rect 12667 10764 12900 10792
rect 12667 10761 12679 10764
rect 12621 10755 12679 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 18230 10792 18236 10804
rect 15344 10764 18236 10792
rect 15344 10752 15350 10764
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19521 10795 19579 10801
rect 19521 10792 19533 10795
rect 19392 10764 19533 10792
rect 19392 10752 19398 10764
rect 19521 10761 19533 10764
rect 19567 10761 19579 10795
rect 19521 10755 19579 10761
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 22612 10764 24900 10792
rect 22612 10752 22618 10764
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10693 5871 10727
rect 5813 10687 5871 10693
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 7834 10724 7840 10736
rect 7340 10696 7840 10724
rect 7340 10684 7346 10696
rect 7834 10684 7840 10696
rect 7892 10684 7898 10736
rect 8021 10727 8079 10733
rect 8021 10693 8033 10727
rect 8067 10724 8079 10727
rect 9401 10727 9459 10733
rect 9401 10724 9413 10727
rect 8067 10696 9413 10724
rect 8067 10693 8079 10696
rect 8021 10687 8079 10693
rect 9401 10693 9413 10696
rect 9447 10724 9459 10727
rect 9447 10696 14136 10724
rect 9447 10693 9459 10696
rect 9401 10687 9459 10693
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 2424 10628 3249 10656
rect 934 10548 940 10600
rect 992 10588 998 10600
rect 2424 10588 2452 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 992 10560 2452 10588
rect 2501 10591 2559 10597
rect 992 10548 998 10560
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3050 10588 3056 10600
rect 2547 10560 3056 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2406 10480 2412 10532
rect 2464 10520 2470 10532
rect 2516 10520 2544 10551
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 5736 10588 5764 10619
rect 6822 10616 6828 10668
rect 6880 10656 6886 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 6880 10628 10149 10656
rect 6880 10616 6886 10628
rect 10137 10625 10149 10628
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 7098 10588 7104 10600
rect 5736 10560 7104 10588
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 7282 10548 7288 10600
rect 7340 10548 7346 10600
rect 7374 10548 7380 10600
rect 7432 10548 7438 10600
rect 7466 10548 7472 10600
rect 7524 10548 7530 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 12452 10588 12480 10619
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 14108 10656 14136 10696
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 14424 10696 15209 10724
rect 14424 10684 14430 10696
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 15197 10687 15255 10693
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 16482 10724 16488 10736
rect 15896 10696 16488 10724
rect 15896 10684 15902 10696
rect 16482 10684 16488 10696
rect 16540 10724 16546 10736
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 16540 10696 17141 10724
rect 16540 10684 16546 10696
rect 17129 10693 17141 10696
rect 17175 10724 17187 10727
rect 18322 10724 18328 10736
rect 17175 10696 18328 10724
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 24112 10727 24170 10733
rect 24112 10693 24124 10727
rect 24158 10724 24170 10727
rect 24762 10724 24768 10736
rect 24158 10696 24768 10724
rect 24158 10693 24170 10696
rect 24112 10687 24170 10693
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 24872 10724 24900 10764
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25225 10795 25283 10801
rect 25225 10792 25237 10795
rect 25188 10764 25237 10792
rect 25188 10752 25194 10764
rect 25225 10761 25237 10764
rect 25271 10761 25283 10795
rect 25225 10755 25283 10761
rect 25682 10752 25688 10804
rect 25740 10752 25746 10804
rect 29914 10752 29920 10804
rect 29972 10792 29978 10804
rect 30374 10792 30380 10804
rect 29972 10764 30380 10792
rect 29972 10752 29978 10764
rect 30116 10733 30144 10764
rect 30374 10752 30380 10764
rect 30432 10752 30438 10804
rect 30469 10795 30527 10801
rect 30469 10761 30481 10795
rect 30515 10792 30527 10795
rect 32582 10792 32588 10804
rect 30515 10764 32588 10792
rect 30515 10761 30527 10764
rect 30469 10755 30527 10761
rect 32582 10752 32588 10764
rect 32640 10752 32646 10804
rect 37642 10752 37648 10804
rect 37700 10792 37706 10804
rect 37737 10795 37795 10801
rect 37737 10792 37749 10795
rect 37700 10764 37749 10792
rect 37700 10752 37706 10764
rect 37737 10761 37749 10764
rect 37783 10761 37795 10795
rect 37737 10755 37795 10761
rect 42978 10752 42984 10804
rect 43036 10752 43042 10804
rect 44266 10752 44272 10804
rect 44324 10752 44330 10804
rect 30101 10727 30159 10733
rect 24872 10696 26188 10724
rect 14458 10656 14464 10668
rect 12768 10628 13952 10656
rect 14108 10628 14464 10656
rect 12768 10616 12774 10628
rect 13814 10588 13820 10600
rect 12452 10560 13820 10588
rect 8757 10551 8815 10557
rect 2464 10492 2544 10520
rect 2464 10480 2470 10492
rect 2682 10480 2688 10532
rect 2740 10520 2746 10532
rect 4062 10520 4068 10532
rect 2740 10492 4068 10520
rect 2740 10480 2746 10492
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 8772 10520 8800 10551
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 13924 10588 13952 10628
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 16850 10616 16856 10668
rect 16908 10616 16914 10668
rect 18414 10665 18420 10668
rect 18408 10619 18420 10665
rect 18414 10616 18420 10619
rect 18472 10616 18478 10668
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 23845 10659 23903 10665
rect 23845 10656 23857 10659
rect 23532 10628 23857 10656
rect 23532 10616 23538 10628
rect 23845 10625 23857 10628
rect 23891 10625 23903 10659
rect 23845 10619 23903 10625
rect 24670 10616 24676 10668
rect 24728 10656 24734 10668
rect 24728 10628 24900 10656
rect 24728 10616 24734 10628
rect 14918 10588 14924 10600
rect 13924 10560 14924 10588
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 17920 10560 18153 10588
rect 17920 10548 17926 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 24872 10588 24900 10628
rect 25130 10616 25136 10668
rect 25188 10656 25194 10668
rect 26160 10665 26188 10696
rect 30101 10693 30113 10727
rect 30147 10693 30159 10727
rect 30101 10687 30159 10693
rect 30193 10727 30251 10733
rect 30193 10693 30205 10727
rect 30239 10724 30251 10727
rect 31018 10724 31024 10736
rect 30239 10696 31024 10724
rect 30239 10693 30251 10696
rect 30193 10687 30251 10693
rect 31018 10684 31024 10696
rect 31076 10684 31082 10736
rect 31205 10727 31263 10733
rect 31205 10693 31217 10727
rect 31251 10724 31263 10727
rect 35526 10724 35532 10736
rect 31251 10696 32260 10724
rect 31251 10693 31263 10696
rect 31205 10687 31263 10693
rect 26053 10659 26111 10665
rect 26053 10656 26065 10659
rect 25188 10628 26065 10656
rect 25188 10616 25194 10628
rect 26053 10625 26065 10628
rect 26099 10625 26111 10659
rect 26053 10619 26111 10625
rect 26145 10659 26203 10665
rect 26145 10625 26157 10659
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 29638 10616 29644 10668
rect 29696 10656 29702 10668
rect 29917 10659 29975 10665
rect 29917 10656 29929 10659
rect 29696 10628 29929 10656
rect 29696 10616 29702 10628
rect 29917 10625 29929 10628
rect 29963 10625 29975 10659
rect 29917 10619 29975 10625
rect 30285 10659 30343 10665
rect 30285 10625 30297 10659
rect 30331 10625 30343 10659
rect 30285 10619 30343 10625
rect 31113 10659 31171 10665
rect 31113 10625 31125 10659
rect 31159 10625 31171 10659
rect 31113 10619 31171 10625
rect 25869 10591 25927 10597
rect 25869 10588 25881 10591
rect 24872 10560 25881 10588
rect 18141 10551 18199 10557
rect 25869 10557 25881 10560
rect 25915 10557 25927 10591
rect 25869 10551 25927 10557
rect 25961 10591 26019 10597
rect 25961 10557 25973 10591
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 4672 10492 8800 10520
rect 4672 10480 4678 10492
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3329 10455 3387 10461
rect 3329 10452 3341 10455
rect 3016 10424 3341 10452
rect 3016 10412 3022 10424
rect 3329 10421 3341 10424
rect 3375 10421 3387 10455
rect 3329 10415 3387 10421
rect 7101 10455 7159 10461
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 7466 10452 7472 10464
rect 7147 10424 7472 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10594 10452 10600 10464
rect 9824 10424 10600 10452
rect 9824 10412 9830 10424
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 24578 10412 24584 10464
rect 24636 10452 24642 10464
rect 25976 10452 26004 10551
rect 30006 10548 30012 10600
rect 30064 10588 30070 10600
rect 30300 10588 30328 10619
rect 30064 10560 30328 10588
rect 30064 10548 30070 10560
rect 31128 10520 31156 10619
rect 31294 10616 31300 10668
rect 31352 10616 31358 10668
rect 31435 10659 31493 10665
rect 31435 10625 31447 10659
rect 31481 10656 31493 10659
rect 31662 10656 31668 10668
rect 31481 10628 31668 10656
rect 31481 10625 31493 10628
rect 31435 10619 31493 10625
rect 31662 10616 31668 10628
rect 31720 10616 31726 10668
rect 31202 10548 31208 10600
rect 31260 10588 31266 10600
rect 31573 10591 31631 10597
rect 31573 10588 31585 10591
rect 31260 10560 31585 10588
rect 31260 10548 31266 10560
rect 31573 10557 31585 10560
rect 31619 10557 31631 10591
rect 32232 10588 32260 10696
rect 32324 10696 35532 10724
rect 32324 10665 32352 10696
rect 35526 10684 35532 10696
rect 35584 10684 35590 10736
rect 35986 10684 35992 10736
rect 36044 10724 36050 10736
rect 36044 10696 38240 10724
rect 36044 10684 36050 10696
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 33962 10616 33968 10668
rect 34020 10616 34026 10668
rect 34149 10659 34207 10665
rect 34149 10625 34161 10659
rect 34195 10656 34207 10659
rect 34514 10656 34520 10668
rect 34195 10628 34520 10656
rect 34195 10625 34207 10628
rect 34149 10619 34207 10625
rect 34514 10616 34520 10628
rect 34572 10616 34578 10668
rect 38010 10616 38016 10668
rect 38068 10656 38074 10668
rect 38105 10659 38163 10665
rect 38105 10656 38117 10659
rect 38068 10628 38117 10656
rect 38068 10616 38074 10628
rect 38105 10625 38117 10628
rect 38151 10625 38163 10659
rect 38212 10656 38240 10696
rect 40402 10684 40408 10736
rect 40460 10724 40466 10736
rect 40926 10727 40984 10733
rect 40926 10724 40938 10727
rect 40460 10696 40938 10724
rect 40460 10684 40466 10696
rect 40926 10693 40938 10696
rect 40972 10693 40984 10727
rect 40926 10687 40984 10693
rect 42334 10684 42340 10736
rect 42392 10724 42398 10736
rect 43349 10727 43407 10733
rect 43349 10724 43361 10727
rect 42392 10696 43361 10724
rect 42392 10684 42398 10696
rect 43349 10693 43361 10696
rect 43395 10693 43407 10727
rect 43349 10687 43407 10693
rect 38212 10628 42564 10656
rect 38105 10619 38163 10625
rect 32490 10588 32496 10600
rect 32232 10560 32496 10588
rect 31573 10551 31631 10557
rect 32490 10548 32496 10560
rect 32548 10548 32554 10600
rect 36722 10548 36728 10600
rect 36780 10588 36786 10600
rect 38197 10591 38255 10597
rect 38197 10588 38209 10591
rect 36780 10560 38209 10588
rect 36780 10548 36786 10560
rect 38197 10557 38209 10560
rect 38243 10557 38255 10591
rect 38197 10551 38255 10557
rect 38378 10548 38384 10600
rect 38436 10548 38442 10600
rect 40678 10548 40684 10600
rect 40736 10548 40742 10600
rect 42536 10588 42564 10628
rect 43162 10616 43168 10668
rect 43220 10616 43226 10668
rect 43254 10616 43260 10668
rect 43312 10616 43318 10668
rect 43438 10616 43444 10668
rect 43496 10665 43502 10668
rect 43496 10659 43525 10665
rect 43513 10625 43525 10659
rect 43496 10619 43525 10625
rect 44177 10659 44235 10665
rect 44177 10625 44189 10659
rect 44223 10625 44235 10659
rect 44177 10619 44235 10625
rect 43496 10616 43502 10619
rect 43625 10591 43683 10597
rect 43625 10588 43637 10591
rect 42536 10560 43637 10588
rect 43625 10557 43637 10560
rect 43671 10557 43683 10591
rect 43625 10551 43683 10557
rect 33042 10520 33048 10532
rect 31128 10492 33048 10520
rect 33042 10480 33048 10492
rect 33100 10480 33106 10532
rect 44192 10520 44220 10619
rect 41984 10492 44220 10520
rect 24636 10424 26004 10452
rect 30929 10455 30987 10461
rect 24636 10412 24642 10424
rect 30929 10421 30941 10455
rect 30975 10452 30987 10455
rect 31938 10452 31944 10464
rect 30975 10424 31944 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 31938 10412 31944 10424
rect 31996 10412 32002 10464
rect 33962 10412 33968 10464
rect 34020 10412 34026 10464
rect 37090 10412 37096 10464
rect 37148 10452 37154 10464
rect 41984 10452 42012 10492
rect 37148 10424 42012 10452
rect 42061 10455 42119 10461
rect 37148 10412 37154 10424
rect 42061 10421 42073 10455
rect 42107 10452 42119 10455
rect 42518 10452 42524 10464
rect 42107 10424 42524 10452
rect 42107 10421 42119 10424
rect 42061 10415 42119 10421
rect 42518 10412 42524 10424
rect 42576 10412 42582 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 2746 10220 22094 10248
rect 2590 10140 2596 10192
rect 2648 10180 2654 10192
rect 2746 10180 2774 10220
rect 2648 10152 2774 10180
rect 2648 10140 2654 10152
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 11054 10180 11060 10192
rect 4120 10152 11060 10180
rect 4120 10140 4126 10152
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 16574 10140 16580 10192
rect 16632 10140 16638 10192
rect 18414 10140 18420 10192
rect 18472 10140 18478 10192
rect 22066 10180 22094 10220
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 22336 10220 22385 10248
rect 22336 10208 22342 10220
rect 22373 10217 22385 10220
rect 22419 10217 22431 10251
rect 22373 10211 22431 10217
rect 23934 10208 23940 10260
rect 23992 10248 23998 10260
rect 24578 10248 24584 10260
rect 23992 10220 24584 10248
rect 23992 10208 23998 10220
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 26694 10208 26700 10260
rect 26752 10248 26758 10260
rect 27249 10251 27307 10257
rect 27249 10248 27261 10251
rect 26752 10220 27261 10248
rect 26752 10208 26758 10220
rect 27249 10217 27261 10220
rect 27295 10217 27307 10251
rect 27249 10211 27307 10217
rect 28445 10251 28503 10257
rect 28445 10217 28457 10251
rect 28491 10248 28503 10251
rect 35986 10248 35992 10260
rect 28491 10220 35992 10248
rect 28491 10217 28503 10220
rect 28445 10211 28503 10217
rect 27893 10183 27951 10189
rect 27893 10180 27905 10183
rect 22066 10152 27905 10180
rect 27893 10149 27905 10152
rect 27939 10180 27951 10183
rect 28460 10180 28488 10211
rect 35986 10208 35992 10220
rect 36044 10208 36050 10260
rect 36722 10208 36728 10260
rect 36780 10208 36786 10260
rect 40218 10208 40224 10260
rect 40276 10248 40282 10260
rect 43165 10251 43223 10257
rect 43165 10248 43177 10251
rect 40276 10220 43177 10248
rect 40276 10208 40282 10220
rect 43165 10217 43177 10220
rect 43211 10217 43223 10251
rect 43165 10211 43223 10217
rect 27939 10152 28488 10180
rect 28629 10183 28687 10189
rect 27939 10149 27951 10152
rect 27893 10143 27951 10149
rect 28629 10149 28641 10183
rect 28675 10149 28687 10183
rect 31294 10180 31300 10192
rect 28629 10143 28687 10149
rect 28920 10152 31300 10180
rect 2958 10072 2964 10124
rect 3016 10072 3022 10124
rect 3050 10072 3056 10124
rect 3108 10072 3114 10124
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 7558 10112 7564 10124
rect 7515 10084 7564 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 9858 10112 9864 10124
rect 9508 10084 9864 10112
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 5902 10044 5908 10056
rect 1627 10016 5908 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 5994 10004 6000 10056
rect 6052 10004 6058 10056
rect 7098 10004 7104 10056
rect 7156 10004 7162 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8202 10044 8208 10056
rect 7883 10016 8208 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9508 10053 9536 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 11664 10084 12357 10112
rect 11664 10072 11670 10084
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 16482 10072 16488 10124
rect 16540 10112 16546 10124
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 16540 10084 16773 10112
rect 16540 10072 16546 10084
rect 16761 10081 16773 10084
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10112 17003 10115
rect 17126 10112 17132 10124
rect 16991 10084 17132 10112
rect 16991 10081 17003 10084
rect 16945 10075 17003 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 20993 10115 21051 10121
rect 20993 10112 21005 10115
rect 17920 10084 21005 10112
rect 17920 10072 17926 10084
rect 20993 10081 21005 10084
rect 21039 10081 21051 10115
rect 20993 10075 21051 10081
rect 25314 10072 25320 10124
rect 25372 10112 25378 10124
rect 28644 10112 28672 10143
rect 25372 10084 28672 10112
rect 25372 10072 25378 10084
rect 28920 10056 28948 10152
rect 31294 10140 31300 10152
rect 31352 10140 31358 10192
rect 39025 10183 39083 10189
rect 39025 10149 39037 10183
rect 39071 10180 39083 10183
rect 39850 10180 39856 10192
rect 39071 10152 39856 10180
rect 39071 10149 39083 10152
rect 39025 10143 39083 10149
rect 39850 10140 39856 10152
rect 39908 10140 39914 10192
rect 30282 10072 30288 10124
rect 30340 10112 30346 10124
rect 30837 10115 30895 10121
rect 30837 10112 30849 10115
rect 30340 10084 30849 10112
rect 30340 10072 30346 10084
rect 30837 10081 30849 10084
rect 30883 10112 30895 10115
rect 31754 10112 31760 10124
rect 30883 10084 31760 10112
rect 30883 10081 30895 10084
rect 30837 10075 30895 10081
rect 31754 10072 31760 10084
rect 31812 10112 31818 10124
rect 32033 10115 32091 10121
rect 32033 10112 32045 10115
rect 31812 10084 32045 10112
rect 31812 10072 31818 10084
rect 32033 10081 32045 10084
rect 32079 10081 32091 10115
rect 32033 10075 32091 10081
rect 35342 10072 35348 10124
rect 35400 10072 35406 10124
rect 38378 10072 38384 10124
rect 38436 10112 38442 10124
rect 43717 10115 43775 10121
rect 43717 10112 43729 10115
rect 38436 10084 43729 10112
rect 38436 10072 38442 10084
rect 43717 10081 43729 10084
rect 43763 10081 43775 10115
rect 43717 10075 43775 10081
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 10505 10047 10563 10053
rect 10505 10044 10517 10047
rect 9493 10007 9551 10013
rect 9600 10016 10517 10044
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 992 9948 1869 9976
rect 992 9936 998 9948
rect 1857 9945 1869 9948
rect 1903 9945 1915 9979
rect 1857 9939 1915 9945
rect 6549 9979 6607 9985
rect 6549 9945 6561 9979
rect 6595 9945 6607 9979
rect 6549 9939 6607 9945
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 2501 9911 2559 9917
rect 2501 9908 2513 9911
rect 2464 9880 2513 9908
rect 2464 9868 2470 9880
rect 2501 9877 2513 9880
rect 2547 9877 2559 9911
rect 2501 9871 2559 9877
rect 2866 9868 2872 9920
rect 2924 9868 2930 9920
rect 6564 9908 6592 9939
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 9600 9976 9628 10016
rect 10505 10013 10517 10016
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10044 11023 10047
rect 11790 10044 11796 10056
rect 11011 10016 11796 10044
rect 11011 10013 11023 10016
rect 10965 10007 11023 10013
rect 8352 9948 9628 9976
rect 8352 9936 8358 9948
rect 9766 9936 9772 9988
rect 9824 9936 9830 9988
rect 10318 9936 10324 9988
rect 10376 9976 10382 9988
rect 10980 9976 11008 10007
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 14918 10044 14924 10056
rect 14783 10016 14924 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 10376 9948 11008 9976
rect 11808 9976 11836 10004
rect 12342 9976 12348 9988
rect 11808 9948 12348 9976
rect 10376 9936 10382 9948
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 12612 9979 12670 9985
rect 12612 9945 12624 9979
rect 12658 9976 12670 9979
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 12658 9948 14289 9976
rect 12658 9945 12670 9948
rect 12612 9939 12670 9945
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 14476 9976 14504 10007
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 16666 9976 16672 9988
rect 14476 9948 16672 9976
rect 14277 9939 14335 9945
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 16868 9976 16896 10007
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17310 10044 17316 10056
rect 17092 10016 17316 10044
rect 17092 10004 17098 10016
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10013 18659 10047
rect 18601 10007 18659 10013
rect 17770 9976 17776 9988
rect 16868 9948 17776 9976
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 18616 9976 18644 10007
rect 18874 10004 18880 10056
rect 18932 10004 18938 10056
rect 21266 10053 21272 10056
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 21260 10044 21272 10053
rect 19475 10016 21128 10044
rect 21227 10016 21272 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 19242 9976 19248 9988
rect 18616 9948 19248 9976
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9945 19763 9979
rect 21100 9976 21128 10016
rect 21260 10007 21272 10016
rect 21266 10004 21272 10007
rect 21324 10004 21330 10056
rect 24670 10004 24676 10056
rect 24728 10044 24734 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 24728 10016 24777 10044
rect 24728 10004 24734 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 24857 10047 24915 10053
rect 24857 10013 24869 10047
rect 24903 10044 24915 10047
rect 26142 10044 26148 10056
rect 24903 10016 26148 10044
rect 24903 10013 24915 10016
rect 24857 10007 24915 10013
rect 22094 9976 22100 9988
rect 21100 9948 22100 9976
rect 19705 9939 19763 9945
rect 6638 9908 6644 9920
rect 6564 9880 6644 9908
rect 6638 9868 6644 9880
rect 6696 9908 6702 9920
rect 9674 9908 9680 9920
rect 6696 9880 9680 9908
rect 6696 9868 6702 9880
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 10008 9880 13737 9908
rect 10008 9868 10014 9880
rect 13725 9877 13737 9880
rect 13771 9908 13783 9911
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 13771 9880 14657 9908
rect 13771 9877 13783 9880
rect 13725 9871 13783 9877
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 16816 9880 18797 9908
rect 16816 9868 16822 9880
rect 18785 9877 18797 9880
rect 18831 9908 18843 9911
rect 19720 9908 19748 9939
rect 22094 9936 22100 9948
rect 22152 9936 22158 9988
rect 20070 9908 20076 9920
rect 18831 9880 20076 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 20990 9868 20996 9920
rect 21048 9908 21054 9920
rect 24872 9908 24900 10007
rect 26142 10004 26148 10016
rect 26200 10004 26206 10056
rect 27062 10004 27068 10056
rect 27120 10044 27126 10056
rect 27157 10047 27215 10053
rect 27157 10044 27169 10047
rect 27120 10016 27169 10044
rect 27120 10004 27126 10016
rect 27157 10013 27169 10016
rect 27203 10013 27215 10047
rect 27157 10007 27215 10013
rect 27338 10004 27344 10056
rect 27396 10004 27402 10056
rect 28902 10044 28908 10056
rect 28276 10016 28908 10044
rect 25038 9936 25044 9988
rect 25096 9976 25102 9988
rect 25317 9979 25375 9985
rect 25317 9976 25329 9979
rect 25096 9948 25329 9976
rect 25096 9936 25102 9948
rect 25317 9945 25329 9948
rect 25363 9976 25375 9979
rect 27706 9976 27712 9988
rect 25363 9948 27712 9976
rect 25363 9945 25375 9948
rect 25317 9939 25375 9945
rect 27706 9936 27712 9948
rect 27764 9936 27770 9988
rect 28276 9985 28304 10016
rect 28902 10004 28908 10016
rect 28960 10004 28966 10056
rect 30098 10004 30104 10056
rect 30156 10004 30162 10056
rect 31938 10004 31944 10056
rect 31996 10044 32002 10056
rect 32289 10047 32347 10053
rect 32289 10044 32301 10047
rect 31996 10016 32301 10044
rect 31996 10004 32002 10016
rect 32289 10013 32301 10016
rect 32335 10013 32347 10047
rect 34514 10044 34520 10056
rect 32289 10007 32347 10013
rect 33060 10016 34520 10044
rect 28261 9979 28319 9985
rect 28261 9945 28273 9979
rect 28307 9945 28319 9979
rect 28261 9939 28319 9945
rect 28477 9979 28535 9985
rect 28477 9945 28489 9979
rect 28523 9976 28535 9979
rect 28994 9976 29000 9988
rect 28523 9948 29000 9976
rect 28523 9945 28535 9948
rect 28477 9939 28535 9945
rect 28994 9936 29000 9948
rect 29052 9936 29058 9988
rect 21048 9880 24900 9908
rect 21048 9868 21054 9880
rect 26326 9868 26332 9920
rect 26384 9908 26390 9920
rect 31570 9908 31576 9920
rect 26384 9880 31576 9908
rect 26384 9868 26390 9880
rect 31570 9868 31576 9880
rect 31628 9908 31634 9920
rect 31754 9908 31760 9920
rect 31628 9880 31760 9908
rect 31628 9868 31634 9880
rect 31754 9868 31760 9880
rect 31812 9908 31818 9920
rect 33060 9908 33088 10016
rect 34514 10004 34520 10016
rect 34572 10004 34578 10056
rect 35360 10044 35388 10072
rect 37182 10044 37188 10056
rect 35360 10016 37188 10044
rect 37182 10004 37188 10016
rect 37240 10004 37246 10056
rect 37458 10053 37464 10056
rect 37452 10044 37464 10053
rect 37419 10016 37464 10044
rect 37452 10007 37464 10016
rect 37458 10004 37464 10007
rect 37516 10004 37522 10056
rect 38838 10004 38844 10056
rect 38896 10044 38902 10056
rect 39301 10047 39359 10053
rect 39301 10044 39313 10047
rect 38896 10016 39313 10044
rect 38896 10004 38902 10016
rect 39301 10013 39313 10016
rect 39347 10013 39359 10047
rect 39301 10007 39359 10013
rect 33962 9936 33968 9988
rect 34020 9976 34026 9988
rect 35590 9979 35648 9985
rect 35590 9976 35602 9979
rect 34020 9948 35602 9976
rect 34020 9936 34026 9948
rect 35590 9945 35602 9948
rect 35636 9945 35648 9979
rect 35590 9939 35648 9945
rect 39022 9936 39028 9988
rect 39080 9936 39086 9988
rect 39206 9936 39212 9988
rect 39264 9936 39270 9988
rect 31812 9880 33088 9908
rect 33413 9911 33471 9917
rect 31812 9868 31818 9880
rect 33413 9877 33425 9911
rect 33459 9908 33471 9911
rect 33686 9908 33692 9920
rect 33459 9880 33692 9908
rect 33459 9877 33471 9880
rect 33413 9871 33471 9877
rect 33686 9868 33692 9880
rect 33744 9868 33750 9920
rect 33870 9868 33876 9920
rect 33928 9908 33934 9920
rect 38010 9908 38016 9920
rect 33928 9880 38016 9908
rect 33928 9868 33934 9880
rect 38010 9868 38016 9880
rect 38068 9908 38074 9920
rect 38565 9911 38623 9917
rect 38565 9908 38577 9911
rect 38068 9880 38577 9908
rect 38068 9868 38074 9880
rect 38565 9877 38577 9880
rect 38611 9877 38623 9911
rect 38565 9871 38623 9877
rect 42518 9868 42524 9920
rect 42576 9908 42582 9920
rect 43530 9908 43536 9920
rect 42576 9880 43536 9908
rect 42576 9868 42582 9880
rect 43530 9868 43536 9880
rect 43588 9868 43594 9920
rect 43622 9868 43628 9920
rect 43680 9868 43686 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 8205 9707 8263 9713
rect 6512 9676 8156 9704
rect 6512 9664 6518 9676
rect 2148 9608 2774 9636
rect 2148 9577 2176 9608
rect 2406 9577 2412 9580
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2400 9568 2412 9577
rect 2367 9540 2412 9568
rect 2133 9531 2191 9537
rect 2400 9531 2412 9540
rect 2406 9528 2412 9531
rect 2464 9528 2470 9580
rect 2746 9568 2774 9608
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 6604 9608 7021 9636
rect 6604 9596 6610 9608
rect 7009 9605 7021 9608
rect 7055 9605 7067 9639
rect 8128 9636 8156 9676
rect 8205 9673 8217 9707
rect 8251 9704 8263 9707
rect 8294 9704 8300 9716
rect 8251 9676 8300 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 9950 9704 9956 9716
rect 8404 9676 9956 9704
rect 8404 9636 8432 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 17678 9704 17684 9716
rect 16632 9676 17684 9704
rect 16632 9664 16638 9676
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 26418 9704 26424 9716
rect 26344 9676 26424 9704
rect 8128 9608 8432 9636
rect 9401 9639 9459 9645
rect 7009 9599 7067 9605
rect 9401 9605 9413 9639
rect 9447 9636 9459 9639
rect 9490 9636 9496 9648
rect 9447 9608 9496 9636
rect 9447 9605 9459 9608
rect 9401 9599 9459 9605
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 9606 9639 9664 9645
rect 9606 9605 9618 9639
rect 9652 9636 9664 9639
rect 9652 9605 9674 9636
rect 9606 9599 9674 9605
rect 4614 9568 4620 9580
rect 2746 9540 4620 9568
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4884 9571 4942 9577
rect 4884 9537 4896 9571
rect 4930 9568 4942 9571
rect 5442 9568 5448 9580
rect 4930 9540 5448 9568
rect 4930 9537 4942 9540
rect 4884 9531 4942 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7892 9540 8125 9568
rect 7892 9528 7898 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8481 9571 8539 9577
rect 8481 9568 8493 9571
rect 8260 9540 8493 9568
rect 8260 9528 8266 9540
rect 8481 9537 8493 9540
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 8297 9503 8355 9509
rect 8297 9469 8309 9503
rect 8343 9500 8355 9503
rect 8386 9500 8392 9512
rect 8343 9472 8392 9500
rect 8343 9469 8355 9472
rect 8297 9463 8355 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 5997 9435 6055 9441
rect 5997 9432 6009 9435
rect 5960 9404 6009 9432
rect 5960 9392 5966 9404
rect 5997 9401 6009 9404
rect 6043 9401 6055 9435
rect 8478 9432 8484 9444
rect 5997 9395 6055 9401
rect 6104 9404 8484 9432
rect 2866 9324 2872 9376
rect 2924 9364 2930 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 2924 9336 3525 9364
rect 2924 9324 2930 9336
rect 3513 9333 3525 9336
rect 3559 9364 3571 9367
rect 3878 9364 3884 9376
rect 3559 9336 3884 9364
rect 3559 9333 3571 9336
rect 3513 9327 3571 9333
rect 3878 9324 3884 9336
rect 3936 9364 3942 9376
rect 6104 9364 6132 9404
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 9646 9432 9674 9599
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 9916 9608 10701 9636
rect 9916 9596 9922 9608
rect 10689 9605 10701 9608
rect 10735 9605 10747 9639
rect 10689 9599 10747 9605
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11112 9608 12434 9636
rect 11112 9596 11118 9608
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 10560 9540 12173 9568
rect 10560 9528 10566 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12406 9568 12434 9608
rect 16942 9596 16948 9648
rect 17000 9636 17006 9648
rect 17098 9639 17156 9645
rect 17098 9636 17110 9639
rect 17000 9608 17110 9636
rect 17000 9596 17006 9608
rect 17098 9605 17110 9608
rect 17144 9605 17156 9639
rect 17098 9599 17156 9605
rect 18322 9596 18328 9648
rect 18380 9636 18386 9648
rect 20901 9639 20959 9645
rect 20901 9636 20913 9639
rect 18380 9608 20913 9636
rect 18380 9596 18386 9608
rect 20901 9605 20913 9608
rect 20947 9636 20959 9639
rect 21082 9636 21088 9648
rect 20947 9608 21088 9636
rect 20947 9605 20959 9608
rect 20901 9599 20959 9605
rect 21082 9596 21088 9608
rect 21140 9636 21146 9648
rect 21140 9608 22094 9636
rect 21140 9596 21146 9608
rect 15194 9568 15200 9580
rect 12406 9540 15200 9568
rect 12253 9531 12311 9537
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 12268 9500 12296 9531
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15286 9528 15292 9580
rect 15344 9528 15350 9580
rect 15470 9528 15476 9580
rect 15528 9528 15534 9580
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 19978 9568 19984 9580
rect 17460 9540 19984 9568
rect 17460 9528 17466 9540
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20990 9528 20996 9580
rect 21048 9528 21054 9580
rect 15304 9500 15332 9528
rect 10652 9472 15332 9500
rect 16853 9503 16911 9509
rect 10652 9460 10658 9472
rect 16853 9469 16865 9503
rect 16899 9469 16911 9503
rect 22066 9500 22094 9608
rect 22278 9596 22284 9648
rect 22336 9596 22342 9648
rect 25133 9639 25191 9645
rect 25133 9605 25145 9639
rect 25179 9636 25191 9639
rect 25961 9639 26019 9645
rect 25961 9636 25973 9639
rect 25179 9608 25973 9636
rect 25179 9605 25191 9608
rect 25133 9599 25191 9605
rect 25961 9605 25973 9608
rect 26007 9605 26019 9639
rect 25961 9599 26019 9605
rect 22296 9568 22324 9596
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 22296 9540 22385 9568
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9568 22523 9571
rect 22554 9568 22560 9580
rect 22511 9540 22560 9568
rect 22511 9537 22523 9540
rect 22465 9531 22523 9537
rect 22554 9528 22560 9540
rect 22612 9528 22618 9580
rect 25314 9528 25320 9580
rect 25372 9528 25378 9580
rect 26234 9528 26240 9580
rect 26292 9528 26298 9580
rect 26344 9577 26372 9676
rect 26418 9664 26424 9676
rect 26476 9704 26482 9716
rect 27062 9704 27068 9716
rect 26476 9676 27068 9704
rect 26476 9664 26482 9676
rect 27062 9664 27068 9676
rect 27120 9664 27126 9716
rect 30006 9664 30012 9716
rect 30064 9704 30070 9716
rect 31846 9704 31852 9716
rect 30064 9676 31852 9704
rect 30064 9664 30070 9676
rect 31846 9664 31852 9676
rect 31904 9664 31910 9716
rect 39022 9664 39028 9716
rect 39080 9704 39086 9716
rect 39393 9707 39451 9713
rect 39393 9704 39405 9707
rect 39080 9676 39405 9704
rect 39080 9664 39086 9676
rect 39393 9673 39405 9676
rect 39439 9673 39451 9707
rect 39393 9667 39451 9673
rect 43254 9664 43260 9716
rect 43312 9704 43318 9716
rect 43990 9704 43996 9716
rect 43312 9676 43996 9704
rect 43312 9664 43318 9676
rect 43990 9664 43996 9676
rect 44048 9664 44054 9716
rect 26694 9636 26700 9648
rect 26436 9608 26700 9636
rect 26436 9577 26464 9608
rect 26694 9596 26700 9608
rect 26752 9596 26758 9648
rect 28350 9636 28356 9648
rect 27448 9608 28356 9636
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 26602 9528 26608 9580
rect 26660 9528 26666 9580
rect 27448 9577 27476 9608
rect 28350 9596 28356 9608
rect 28408 9596 28414 9648
rect 28810 9636 28816 9648
rect 28552 9608 28816 9636
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27526 9571 27584 9577
rect 27526 9537 27538 9571
rect 27572 9537 27584 9571
rect 27526 9531 27584 9537
rect 22189 9503 22247 9509
rect 22189 9500 22201 9503
rect 22066 9472 22201 9500
rect 16853 9463 16911 9469
rect 22189 9469 22201 9472
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 11054 9432 11060 9444
rect 9646 9404 11060 9432
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 16482 9432 16488 9444
rect 15160 9404 16488 9432
rect 15160 9392 15166 9404
rect 16482 9392 16488 9404
rect 16540 9432 16546 9444
rect 16868 9432 16896 9463
rect 16540 9404 16896 9432
rect 22204 9432 22232 9463
rect 22278 9460 22284 9512
rect 22336 9460 22342 9512
rect 26252 9500 26280 9528
rect 27338 9500 27344 9512
rect 26252 9472 27344 9500
rect 27338 9460 27344 9472
rect 27396 9500 27402 9512
rect 27540 9500 27568 9531
rect 27706 9528 27712 9580
rect 27764 9528 27770 9580
rect 27798 9528 27804 9580
rect 27856 9528 27862 9580
rect 27939 9571 27997 9577
rect 27939 9537 27951 9571
rect 27985 9568 27997 9571
rect 28552 9568 28580 9608
rect 28810 9596 28816 9608
rect 28868 9596 28874 9648
rect 28994 9596 29000 9648
rect 29052 9596 29058 9648
rect 30098 9596 30104 9648
rect 30156 9636 30162 9648
rect 35989 9639 36047 9645
rect 35989 9636 36001 9639
rect 30156 9608 36001 9636
rect 30156 9596 30162 9608
rect 35989 9605 36001 9608
rect 36035 9636 36047 9639
rect 36446 9636 36452 9648
rect 36035 9608 36452 9636
rect 36035 9605 36047 9608
rect 35989 9599 36047 9605
rect 36446 9596 36452 9608
rect 36504 9596 36510 9648
rect 37182 9596 37188 9648
rect 37240 9636 37246 9648
rect 39945 9639 40003 9645
rect 37240 9608 39344 9636
rect 37240 9596 37246 9608
rect 27985 9540 28580 9568
rect 27985 9537 27997 9540
rect 27939 9531 27997 9537
rect 28626 9528 28632 9580
rect 28684 9528 28690 9580
rect 29012 9568 29040 9596
rect 30834 9568 30840 9580
rect 29012 9540 30840 9568
rect 30834 9528 30840 9540
rect 30892 9528 30898 9580
rect 31478 9528 31484 9580
rect 31536 9528 31542 9580
rect 31665 9571 31723 9577
rect 31665 9537 31677 9571
rect 31711 9568 31723 9571
rect 31754 9568 31760 9580
rect 31711 9540 31760 9568
rect 31711 9537 31723 9540
rect 31665 9531 31723 9537
rect 31754 9528 31760 9540
rect 31812 9528 31818 9580
rect 32122 9528 32128 9580
rect 32180 9568 32186 9580
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 32180 9540 32321 9568
rect 32180 9528 32186 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9537 32551 9571
rect 32493 9531 32551 9537
rect 27396 9472 27568 9500
rect 30929 9503 30987 9509
rect 27396 9460 27402 9472
rect 30929 9469 30941 9503
rect 30975 9500 30987 9503
rect 31938 9500 31944 9512
rect 30975 9472 31944 9500
rect 30975 9469 30987 9472
rect 30929 9463 30987 9469
rect 31938 9460 31944 9472
rect 31996 9460 32002 9512
rect 32214 9460 32220 9512
rect 32272 9500 32278 9512
rect 32508 9500 32536 9531
rect 33686 9528 33692 9580
rect 33744 9568 33750 9580
rect 33781 9571 33839 9577
rect 33781 9568 33793 9571
rect 33744 9540 33793 9568
rect 33744 9528 33750 9540
rect 33781 9537 33793 9540
rect 33827 9537 33839 9571
rect 33781 9531 33839 9537
rect 38654 9528 38660 9580
rect 38712 9568 38718 9580
rect 38841 9571 38899 9577
rect 38841 9568 38853 9571
rect 38712 9540 38853 9568
rect 38712 9528 38718 9540
rect 38841 9537 38853 9540
rect 38887 9537 38899 9571
rect 38841 9531 38899 9537
rect 39022 9528 39028 9580
rect 39080 9528 39086 9580
rect 39117 9571 39175 9577
rect 39117 9537 39129 9571
rect 39163 9537 39175 9571
rect 39117 9531 39175 9537
rect 32272 9472 32536 9500
rect 33873 9503 33931 9509
rect 32272 9460 32278 9472
rect 33873 9469 33885 9503
rect 33919 9500 33931 9503
rect 33962 9500 33968 9512
rect 33919 9472 33968 9500
rect 33919 9469 33931 9472
rect 33873 9463 33931 9469
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 34054 9460 34060 9512
rect 34112 9460 34118 9512
rect 36078 9460 36084 9512
rect 36136 9500 36142 9512
rect 36725 9503 36783 9509
rect 36725 9500 36737 9503
rect 36136 9472 36737 9500
rect 36136 9460 36142 9472
rect 36725 9469 36737 9472
rect 36771 9469 36783 9503
rect 36725 9463 36783 9469
rect 23474 9432 23480 9444
rect 22204 9404 23480 9432
rect 16540 9392 16546 9404
rect 23474 9392 23480 9404
rect 23532 9432 23538 9444
rect 24670 9432 24676 9444
rect 23532 9404 24676 9432
rect 23532 9392 23538 9404
rect 24670 9392 24676 9404
rect 24728 9392 24734 9444
rect 28074 9392 28080 9444
rect 28132 9392 28138 9444
rect 28626 9392 28632 9444
rect 28684 9432 28690 9444
rect 36538 9432 36544 9444
rect 28684 9404 36544 9432
rect 28684 9392 28690 9404
rect 36538 9392 36544 9404
rect 36596 9392 36602 9444
rect 3936 9336 6132 9364
rect 3936 9324 3942 9336
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 8168 9336 8401 9364
rect 8168 9324 8174 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 8904 9336 9597 9364
rect 8904 9324 8910 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11756 9336 11989 9364
rect 11756 9324 11762 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 11977 9327 12035 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12894 9364 12900 9376
rect 12483 9336 12900 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 15381 9367 15439 9373
rect 15381 9333 15393 9367
rect 15427 9364 15439 9367
rect 16022 9364 16028 9376
rect 15427 9336 16028 9364
rect 15427 9333 15439 9336
rect 15381 9327 15439 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 17184 9336 18245 9364
rect 17184 9324 17190 9336
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 21177 9367 21235 9373
rect 21177 9333 21189 9367
rect 21223 9364 21235 9367
rect 21266 9364 21272 9376
rect 21223 9336 21272 9364
rect 21223 9333 21235 9336
rect 21177 9327 21235 9333
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21450 9324 21456 9376
rect 21508 9364 21514 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21508 9336 22017 9364
rect 21508 9324 21514 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 25406 9324 25412 9376
rect 25464 9364 25470 9376
rect 25501 9367 25559 9373
rect 25501 9364 25513 9367
rect 25464 9336 25513 9364
rect 25464 9324 25470 9336
rect 25501 9333 25513 9336
rect 25547 9333 25559 9367
rect 25501 9327 25559 9333
rect 31478 9324 31484 9376
rect 31536 9324 31542 9376
rect 32309 9367 32367 9373
rect 32309 9333 32321 9367
rect 32355 9364 32367 9367
rect 32950 9364 32956 9376
rect 32355 9336 32956 9364
rect 32355 9333 32367 9336
rect 32309 9327 32367 9333
rect 32950 9324 32956 9336
rect 33008 9324 33014 9376
rect 33042 9324 33048 9376
rect 33100 9364 33106 9376
rect 33413 9367 33471 9373
rect 33413 9364 33425 9367
rect 33100 9336 33425 9364
rect 33100 9324 33106 9336
rect 33413 9333 33425 9336
rect 33459 9333 33471 9367
rect 39132 9364 39160 9531
rect 39206 9528 39212 9580
rect 39264 9528 39270 9580
rect 39316 9500 39344 9608
rect 39945 9605 39957 9639
rect 39991 9636 40003 9639
rect 40926 9639 40984 9645
rect 40926 9636 40938 9639
rect 39991 9608 40938 9636
rect 39991 9605 40003 9608
rect 39945 9599 40003 9605
rect 40926 9605 40938 9608
rect 40972 9605 40984 9639
rect 40926 9599 40984 9605
rect 39850 9528 39856 9580
rect 39908 9528 39914 9580
rect 40037 9571 40095 9577
rect 40037 9537 40049 9571
rect 40083 9568 40095 9571
rect 40770 9568 40776 9580
rect 40083 9540 40776 9568
rect 40083 9537 40095 9540
rect 40037 9531 40095 9537
rect 40770 9528 40776 9540
rect 40828 9528 40834 9580
rect 40678 9500 40684 9512
rect 39316 9472 40684 9500
rect 40678 9460 40684 9472
rect 40736 9460 40742 9512
rect 42061 9435 42119 9441
rect 42061 9401 42073 9435
rect 42107 9432 42119 9435
rect 43622 9432 43628 9444
rect 42107 9404 43628 9432
rect 42107 9401 42119 9404
rect 42061 9395 42119 9401
rect 40954 9364 40960 9376
rect 39132 9336 40960 9364
rect 33413 9327 33471 9333
rect 40954 9324 40960 9336
rect 41012 9364 41018 9376
rect 42076 9364 42104 9395
rect 43622 9392 43628 9404
rect 43680 9392 43686 9444
rect 41012 9336 42104 9364
rect 41012 9324 41018 9336
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 2498 9120 2504 9172
rect 2556 9120 2562 9172
rect 3234 9120 3240 9172
rect 3292 9120 3298 9172
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7156 9132 7481 9160
rect 7156 9120 7162 9132
rect 7469 9129 7481 9132
rect 7515 9160 7527 9163
rect 8110 9160 8116 9172
rect 7515 9132 8116 9160
rect 7515 9129 7527 9132
rect 7469 9123 7527 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 9582 9160 9588 9172
rect 8352 9132 9588 9160
rect 8352 9120 8358 9132
rect 9582 9120 9588 9132
rect 9640 9160 9646 9172
rect 12158 9160 12164 9172
rect 9640 9132 12164 9160
rect 9640 9120 9646 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 28626 9160 28632 9172
rect 12400 9132 28632 9160
rect 12400 9120 12406 9132
rect 28626 9120 28632 9132
rect 28684 9120 28690 9172
rect 30650 9160 30656 9172
rect 29748 9132 30656 9160
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 10502 9092 10508 9104
rect 1903 9064 10508 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 12805 9095 12863 9101
rect 12805 9061 12817 9095
rect 12851 9092 12863 9095
rect 14274 9092 14280 9104
rect 12851 9064 14280 9092
rect 12851 9061 12863 9064
rect 12805 9055 12863 9061
rect 1118 8984 1124 9036
rect 1176 9024 1182 9036
rect 1176 8996 2774 9024
rect 1176 8984 1182 8996
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 2409 8959 2467 8965
rect 2409 8956 2421 8959
rect 992 8928 2421 8956
rect 992 8916 998 8928
rect 2409 8925 2421 8928
rect 2455 8925 2467 8959
rect 2746 8956 2774 8996
rect 5644 8996 9076 9024
rect 5644 8965 5672 8996
rect 3145 8959 3203 8965
rect 3145 8956 3157 8959
rect 2746 8928 3157 8956
rect 2409 8919 2467 8925
rect 3145 8925 3157 8928
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5776 8928 5917 8956
rect 5776 8916 5782 8928
rect 5905 8925 5917 8928
rect 5951 8956 5963 8959
rect 6546 8956 6552 8968
rect 5951 8928 6552 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6546 8916 6552 8928
rect 6604 8956 6610 8968
rect 6604 8928 7696 8956
rect 6604 8916 6610 8928
rect 1026 8848 1032 8900
rect 1084 8888 1090 8900
rect 1673 8891 1731 8897
rect 1673 8888 1685 8891
rect 1084 8860 1685 8888
rect 1084 8848 1090 8860
rect 1673 8857 1685 8860
rect 1719 8857 1731 8891
rect 1673 8851 1731 8857
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7285 8891 7343 8897
rect 7285 8888 7297 8891
rect 7248 8860 7297 8888
rect 7248 8848 7254 8860
rect 7285 8857 7297 8860
rect 7331 8857 7343 8891
rect 7285 8851 7343 8857
rect 7466 8848 7472 8900
rect 7524 8897 7530 8900
rect 7524 8891 7543 8897
rect 7531 8857 7543 8891
rect 7668 8888 7696 8928
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7800 8928 8125 8956
rect 7800 8916 7806 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8662 8888 8668 8900
rect 7668 8860 8668 8888
rect 7524 8851 7543 8857
rect 7524 8848 7530 8851
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 5813 8823 5871 8829
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 5902 8820 5908 8832
rect 5859 8792 5908 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 8294 8820 8300 8832
rect 7699 8792 8300 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 9048 8820 9076 8996
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10008 8996 10180 9024
rect 10008 8984 10014 8996
rect 9858 8916 9864 8968
rect 9916 8916 9922 8968
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10152 8965 10180 8996
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 11514 8956 11520 8968
rect 11471 8928 11520 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12820 8956 12848 9055
rect 14274 9052 14280 9064
rect 14332 9052 14338 9104
rect 16393 9095 16451 9101
rect 16393 9061 16405 9095
rect 16439 9092 16451 9095
rect 16942 9092 16948 9104
rect 16439 9064 16948 9092
rect 16439 9061 16451 9064
rect 16393 9055 16451 9061
rect 16942 9052 16948 9064
rect 17000 9052 17006 9104
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 17494 9092 17500 9104
rect 17276 9064 17500 9092
rect 17276 9052 17282 9064
rect 17494 9052 17500 9064
rect 17552 9092 17558 9104
rect 17773 9095 17831 9101
rect 17773 9092 17785 9095
rect 17552 9064 17785 9092
rect 17552 9052 17558 9064
rect 17773 9061 17785 9064
rect 17819 9061 17831 9095
rect 17773 9055 17831 9061
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 17788 9024 17816 9055
rect 19150 9052 19156 9104
rect 19208 9092 19214 9104
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 19208 9064 21281 9092
rect 19208 9052 19214 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 29748 9092 29776 9132
rect 30650 9120 30656 9132
rect 30708 9120 30714 9172
rect 36538 9120 36544 9172
rect 36596 9160 36602 9172
rect 42242 9160 42248 9172
rect 36596 9132 42248 9160
rect 36596 9120 36602 9132
rect 42242 9120 42248 9132
rect 42300 9120 42306 9172
rect 21269 9055 21327 9061
rect 21376 9064 21772 9092
rect 20346 9024 20352 9036
rect 12952 8996 17264 9024
rect 17788 8996 20352 9024
rect 12952 8984 12958 8996
rect 11624 8928 12848 8956
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11624 8888 11652 8928
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 16574 8956 16580 8968
rect 16172 8928 16580 8956
rect 16172 8916 16178 8928
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16669 8959 16727 8965
rect 16669 8925 16681 8959
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8956 17003 8959
rect 17126 8956 17132 8968
rect 16991 8928 17132 8956
rect 16991 8925 17003 8928
rect 16945 8919 17003 8925
rect 11020 8860 11652 8888
rect 11692 8891 11750 8897
rect 11020 8848 11026 8860
rect 11692 8857 11704 8891
rect 11738 8888 11750 8891
rect 12066 8888 12072 8900
rect 11738 8860 12072 8888
rect 11738 8857 11750 8860
rect 11692 8851 11750 8857
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 16022 8848 16028 8900
rect 16080 8888 16086 8900
rect 16684 8888 16712 8919
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17236 8956 17264 8996
rect 20346 8984 20352 8996
rect 20404 9024 20410 9036
rect 21376 9024 21404 9064
rect 20404 8996 21404 9024
rect 20404 8984 20410 8996
rect 21450 8984 21456 9036
rect 21508 8984 21514 9036
rect 21634 8984 21640 9036
rect 21692 8984 21698 9036
rect 19150 8956 19156 8968
rect 17236 8928 19156 8956
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19260 8928 19441 8956
rect 16080 8860 16712 8888
rect 16080 8848 16086 8860
rect 16758 8848 16764 8900
rect 16816 8888 16822 8900
rect 17037 8891 17095 8897
rect 17037 8888 17049 8891
rect 16816 8860 17049 8888
rect 16816 8848 16822 8860
rect 17037 8857 17049 8860
rect 17083 8857 17095 8891
rect 17037 8851 17095 8857
rect 17589 8891 17647 8897
rect 17589 8857 17601 8891
rect 17635 8857 17647 8891
rect 17589 8851 17647 8857
rect 12158 8820 12164 8832
rect 9048 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12526 8820 12532 8832
rect 12308 8792 12532 8820
rect 12308 8780 12314 8792
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 17604 8820 17632 8851
rect 17678 8848 17684 8900
rect 17736 8888 17742 8900
rect 19260 8888 19288 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 21542 8916 21548 8968
rect 21600 8916 21606 8968
rect 21744 8965 21772 9064
rect 28368 9064 29776 9092
rect 25314 8984 25320 9036
rect 25372 9024 25378 9036
rect 26602 9024 26608 9036
rect 25372 8996 26608 9024
rect 25372 8984 25378 8996
rect 21729 8959 21787 8965
rect 21729 8925 21741 8959
rect 21775 8956 21787 8959
rect 25958 8956 25964 8968
rect 21775 8928 25964 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 26528 8965 26556 8996
rect 26602 8984 26608 8996
rect 26660 8984 26666 9036
rect 28368 8965 28396 9064
rect 32858 9052 32864 9104
rect 32916 9092 32922 9104
rect 36630 9092 36636 9104
rect 32916 9064 36636 9092
rect 32916 9052 32922 9064
rect 36630 9052 36636 9064
rect 36688 9092 36694 9104
rect 38838 9092 38844 9104
rect 36688 9064 38844 9092
rect 36688 9052 36694 9064
rect 38838 9052 38844 9064
rect 38896 9092 38902 9104
rect 38896 9064 40264 9092
rect 38896 9052 38902 9064
rect 37182 8984 37188 9036
rect 37240 8984 37246 9036
rect 40236 9033 40264 9064
rect 40221 9027 40279 9033
rect 40221 8993 40233 9027
rect 40267 8993 40279 9027
rect 40221 8987 40279 8993
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8925 26295 8959
rect 26237 8919 26295 8925
rect 26513 8959 26571 8965
rect 26513 8925 26525 8959
rect 26559 8925 26571 8959
rect 26513 8919 26571 8925
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 17736 8860 19288 8888
rect 17736 8848 17742 8860
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 19705 8891 19763 8897
rect 19705 8888 19717 8891
rect 19392 8860 19717 8888
rect 19392 8848 19398 8860
rect 19705 8857 19717 8860
rect 19751 8888 19763 8891
rect 22094 8888 22100 8900
rect 19751 8860 22100 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 22094 8848 22100 8860
rect 22152 8888 22158 8900
rect 22554 8888 22560 8900
rect 22152 8860 22560 8888
rect 22152 8848 22158 8860
rect 22554 8848 22560 8860
rect 22612 8848 22618 8900
rect 26252 8888 26280 8919
rect 29730 8916 29736 8968
rect 29788 8956 29794 8968
rect 30282 8956 30288 8968
rect 29788 8928 30288 8956
rect 29788 8916 29794 8928
rect 30282 8916 30288 8928
rect 30340 8916 30346 8968
rect 31386 8916 31392 8968
rect 31444 8956 31450 8968
rect 31941 8959 31999 8965
rect 31941 8956 31953 8959
rect 31444 8928 31953 8956
rect 31444 8916 31450 8928
rect 31941 8925 31953 8928
rect 31987 8925 31999 8959
rect 31941 8919 31999 8925
rect 32858 8916 32864 8968
rect 32916 8956 32922 8968
rect 32916 8928 36400 8956
rect 32916 8916 32922 8928
rect 26602 8888 26608 8900
rect 26252 8860 26608 8888
rect 26602 8848 26608 8860
rect 26660 8848 26666 8900
rect 28629 8891 28687 8897
rect 28629 8857 28641 8891
rect 28675 8888 28687 8891
rect 28902 8888 28908 8900
rect 28675 8860 28908 8888
rect 28675 8857 28687 8860
rect 28629 8851 28687 8857
rect 28902 8848 28908 8860
rect 28960 8888 28966 8900
rect 29270 8888 29276 8900
rect 28960 8860 29276 8888
rect 28960 8848 28966 8860
rect 29270 8848 29276 8860
rect 29328 8848 29334 8900
rect 30000 8891 30058 8897
rect 30000 8857 30012 8891
rect 30046 8888 30058 8891
rect 31478 8888 31484 8900
rect 30046 8860 31484 8888
rect 30046 8857 30058 8860
rect 30000 8851 30058 8857
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 31573 8891 31631 8897
rect 31573 8857 31585 8891
rect 31619 8857 31631 8891
rect 31573 8851 31631 8857
rect 31757 8891 31815 8897
rect 31757 8857 31769 8891
rect 31803 8888 31815 8891
rect 32214 8888 32220 8900
rect 31803 8860 32220 8888
rect 31803 8857 31815 8860
rect 31757 8851 31815 8857
rect 12676 8792 17632 8820
rect 26053 8823 26111 8829
rect 12676 8780 12682 8792
rect 26053 8789 26065 8823
rect 26099 8820 26111 8823
rect 26142 8820 26148 8832
rect 26099 8792 26148 8820
rect 26099 8789 26111 8792
rect 26053 8783 26111 8789
rect 26142 8780 26148 8792
rect 26200 8780 26206 8832
rect 26234 8780 26240 8832
rect 26292 8820 26298 8832
rect 26421 8823 26479 8829
rect 26421 8820 26433 8823
rect 26292 8792 26433 8820
rect 26292 8780 26298 8792
rect 26421 8789 26433 8792
rect 26467 8789 26479 8823
rect 26421 8783 26479 8789
rect 29638 8780 29644 8832
rect 29696 8820 29702 8832
rect 31113 8823 31171 8829
rect 31113 8820 31125 8823
rect 29696 8792 31125 8820
rect 29696 8780 29702 8792
rect 31113 8789 31125 8792
rect 31159 8789 31171 8823
rect 31588 8820 31616 8851
rect 32214 8848 32220 8860
rect 32272 8848 32278 8900
rect 33226 8848 33232 8900
rect 33284 8888 33290 8900
rect 35621 8891 35679 8897
rect 35621 8888 35633 8891
rect 33284 8860 35633 8888
rect 33284 8848 33290 8860
rect 35621 8857 35633 8860
rect 35667 8857 35679 8891
rect 36372 8888 36400 8928
rect 36446 8916 36452 8968
rect 36504 8916 36510 8968
rect 37550 8916 37556 8968
rect 37608 8956 37614 8968
rect 40037 8959 40095 8965
rect 40037 8956 40049 8959
rect 37608 8928 40049 8956
rect 37608 8916 37614 8928
rect 40037 8925 40049 8928
rect 40083 8956 40095 8959
rect 40126 8956 40132 8968
rect 40083 8928 40132 8956
rect 40083 8925 40095 8928
rect 40037 8919 40095 8925
rect 40126 8916 40132 8928
rect 40184 8916 40190 8968
rect 39206 8888 39212 8900
rect 36372 8860 39212 8888
rect 35621 8851 35679 8857
rect 39206 8848 39212 8860
rect 39264 8888 39270 8900
rect 40310 8888 40316 8900
rect 39264 8860 40316 8888
rect 39264 8848 39270 8860
rect 40310 8848 40316 8860
rect 40368 8848 40374 8900
rect 32122 8820 32128 8832
rect 31588 8792 32128 8820
rect 31113 8783 31171 8789
rect 32122 8780 32128 8792
rect 32180 8780 32186 8832
rect 34606 8780 34612 8832
rect 34664 8820 34670 8832
rect 34790 8820 34796 8832
rect 34664 8792 34796 8820
rect 34664 8780 34670 8792
rect 34790 8780 34796 8792
rect 34848 8780 34854 8832
rect 35897 8823 35955 8829
rect 35897 8789 35909 8823
rect 35943 8820 35955 8823
rect 37550 8820 37556 8832
rect 35943 8792 37556 8820
rect 35943 8789 35955 8792
rect 35897 8783 35955 8789
rect 37550 8780 37556 8792
rect 37608 8780 37614 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 7800 8588 8769 8616
rect 7800 8576 7806 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 9548 8588 10609 8616
rect 9548 8576 9554 8588
rect 10597 8585 10609 8588
rect 10643 8616 10655 8619
rect 10962 8616 10968 8628
rect 10643 8588 10968 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 12066 8576 12072 8628
rect 12124 8576 12130 8628
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 12216 8588 13829 8616
rect 12216 8576 12222 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16724 8588 17049 8616
rect 16724 8576 16730 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17678 8616 17684 8628
rect 17184 8588 17684 8616
rect 17184 8576 17190 8588
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19484 8588 19901 8616
rect 19484 8576 19490 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 19889 8579 19947 8585
rect 20272 8588 20484 8616
rect 1026 8508 1032 8560
rect 1084 8548 1090 8560
rect 2593 8551 2651 8557
rect 2593 8548 2605 8551
rect 1084 8520 2605 8548
rect 1084 8508 1090 8520
rect 2593 8517 2605 8520
rect 2639 8517 2651 8551
rect 2593 8511 2651 8517
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8548 2835 8551
rect 2823 8520 10180 8548
rect 2823 8517 2835 8520
rect 2777 8511 2835 8517
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 5166 8480 5172 8492
rect 1627 8452 5172 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5626 8480 5632 8492
rect 5307 8452 5632 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 7190 8440 7196 8492
rect 7248 8480 7254 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 7248 8452 7297 8480
rect 7248 8440 7254 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 8966 8483 9024 8489
rect 8966 8480 8978 8483
rect 7852 8452 8978 8480
rect 934 8372 940 8424
rect 992 8412 998 8424
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 992 8384 1777 8412
rect 992 8372 998 8384
rect 1765 8381 1777 8384
rect 1811 8381 1823 8415
rect 1765 8375 1823 8381
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 7852 8412 7880 8452
rect 8966 8449 8978 8452
rect 9012 8449 9024 8483
rect 10152 8480 10180 8520
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 12621 8551 12679 8557
rect 10376 8520 11928 8548
rect 10376 8508 10382 8520
rect 11238 8480 11244 8492
rect 10152 8452 11244 8480
rect 8966 8443 9024 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11900 8489 11928 8520
rect 12621 8517 12633 8551
rect 12667 8548 12679 8551
rect 20272 8548 20300 8588
rect 12667 8520 14872 8548
rect 12667 8517 12679 8520
rect 12621 8511 12679 8517
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12710 8440 12716 8492
rect 12768 8440 12774 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13780 8452 14105 8480
rect 13780 8440 13786 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 14844 8489 14872 8520
rect 17236 8520 20300 8548
rect 20456 8548 20484 8588
rect 22370 8576 22376 8628
rect 22428 8616 22434 8628
rect 22922 8616 22928 8628
rect 22428 8588 22928 8616
rect 22428 8576 22434 8588
rect 22922 8576 22928 8588
rect 22980 8616 22986 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 22980 8588 24041 8616
rect 22980 8576 22986 8588
rect 24029 8585 24041 8588
rect 24075 8585 24087 8619
rect 34790 8616 34796 8628
rect 24029 8579 24087 8585
rect 33612 8588 34796 8616
rect 22554 8548 22560 8560
rect 20456 8520 22560 8548
rect 14829 8483 14887 8489
rect 14240 8452 14780 8480
rect 14240 8440 14246 8452
rect 7524 8384 7880 8412
rect 7524 8372 7530 8384
rect 7926 8372 7932 8424
rect 7984 8372 7990 8424
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 8481 8415 8539 8421
rect 8481 8412 8493 8415
rect 8168 8384 8493 8412
rect 8168 8372 8174 8384
rect 8481 8381 8493 8384
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8846 8372 8852 8424
rect 8904 8372 8910 8424
rect 8956 8384 10364 8412
rect 5442 8304 5448 8356
rect 5500 8304 5506 8356
rect 8386 8304 8392 8356
rect 8444 8344 8450 8356
rect 8864 8344 8892 8372
rect 8956 8356 8984 8384
rect 8444 8316 8892 8344
rect 8444 8304 8450 8316
rect 8938 8304 8944 8356
rect 8996 8304 9002 8356
rect 9125 8347 9183 8353
rect 9125 8313 9137 8347
rect 9171 8344 9183 8347
rect 9950 8344 9956 8356
rect 9171 8316 9956 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9950 8304 9956 8316
rect 10008 8304 10014 8356
rect 10336 8344 10364 8384
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10560 8384 10701 8412
rect 10560 8372 10566 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 10962 8412 10968 8424
rect 10919 8384 10968 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 12728 8344 12756 8440
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 10336 8316 12756 8344
rect 14016 8344 14044 8375
rect 14274 8372 14280 8424
rect 14332 8372 14338 8424
rect 14752 8412 14780 8452
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 17236 8489 17264 8520
rect 22554 8508 22560 8520
rect 22612 8508 22618 8560
rect 22664 8520 25912 8548
rect 17221 8483 17279 8489
rect 14976 8452 16712 8480
rect 14976 8440 14982 8452
rect 15105 8415 15163 8421
rect 15105 8412 15117 8415
rect 14752 8384 15117 8412
rect 15105 8381 15117 8384
rect 15151 8412 15163 8415
rect 16206 8412 16212 8424
rect 15151 8384 16212 8412
rect 15151 8381 15163 8384
rect 15105 8375 15163 8381
rect 16206 8372 16212 8384
rect 16264 8412 16270 8424
rect 16684 8412 16712 8452
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17310 8440 17316 8492
rect 17368 8440 17374 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 19886 8480 19892 8492
rect 18371 8452 19892 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 20346 8440 20352 8492
rect 20404 8440 20410 8492
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 22370 8480 22376 8492
rect 21315 8452 22376 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 22664 8489 22692 8520
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 18156 8412 18184 8440
rect 16264 8384 16620 8412
rect 16684 8384 18184 8412
rect 18785 8415 18843 8421
rect 16264 8372 16270 8384
rect 16482 8344 16488 8356
rect 14016 8316 16488 8344
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 16592 8344 16620 8384
rect 18785 8381 18797 8415
rect 18831 8412 18843 8415
rect 19978 8412 19984 8424
rect 18831 8384 19984 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 17402 8344 17408 8356
rect 16592 8316 17408 8344
rect 17402 8304 17408 8316
rect 17460 8344 17466 8356
rect 20088 8344 20116 8375
rect 20162 8372 20168 8424
rect 20220 8372 20226 8424
rect 20257 8415 20315 8421
rect 20257 8381 20269 8415
rect 20303 8412 20315 8415
rect 20303 8384 21036 8412
rect 20303 8381 20315 8384
rect 20257 8375 20315 8381
rect 20901 8347 20959 8353
rect 20901 8344 20913 8347
rect 17460 8316 20024 8344
rect 20088 8316 20913 8344
rect 17460 8304 17466 8316
rect 10229 8279 10287 8285
rect 10229 8245 10241 8279
rect 10275 8276 10287 8279
rect 10318 8276 10324 8288
rect 10275 8248 10324 8276
rect 10275 8245 10287 8248
rect 10229 8239 10287 8245
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 13998 8276 14004 8288
rect 11756 8248 14004 8276
rect 11756 8236 11762 8248
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 19996 8276 20024 8316
rect 20901 8313 20913 8316
rect 20947 8313 20959 8347
rect 20901 8307 20959 8313
rect 20806 8276 20812 8288
rect 19996 8248 20812 8276
rect 20806 8236 20812 8248
rect 20864 8236 20870 8288
rect 21008 8276 21036 8384
rect 21174 8372 21180 8424
rect 21232 8372 21238 8424
rect 21361 8415 21419 8421
rect 21361 8381 21373 8415
rect 21407 8381 21419 8415
rect 21361 8375 21419 8381
rect 21376 8344 21404 8375
rect 22002 8372 22008 8424
rect 22060 8412 22066 8424
rect 22664 8412 22692 8443
rect 22738 8440 22744 8492
rect 22796 8480 22802 8492
rect 25148 8489 25176 8520
rect 25884 8492 25912 8520
rect 31846 8508 31852 8560
rect 31904 8548 31910 8560
rect 32858 8548 32864 8560
rect 31904 8520 32864 8548
rect 31904 8508 31910 8520
rect 32858 8508 32864 8520
rect 32916 8508 32922 8560
rect 33042 8508 33048 8560
rect 33100 8548 33106 8560
rect 33612 8557 33640 8588
rect 34790 8576 34796 8588
rect 34848 8616 34854 8628
rect 34848 8588 38056 8616
rect 34848 8576 34854 8588
rect 33597 8551 33655 8557
rect 33597 8548 33609 8551
rect 33100 8520 33609 8548
rect 33100 8508 33106 8520
rect 33597 8517 33609 8520
rect 33643 8517 33655 8551
rect 35894 8548 35900 8560
rect 33597 8511 33655 8517
rect 33704 8520 35900 8548
rect 25406 8489 25412 8492
rect 22905 8483 22963 8489
rect 22905 8480 22917 8483
rect 22796 8452 22917 8480
rect 22796 8440 22802 8452
rect 22905 8449 22917 8452
rect 22951 8449 22963 8483
rect 22905 8443 22963 8449
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25400 8480 25412 8489
rect 25367 8452 25412 8480
rect 25133 8443 25191 8449
rect 25400 8443 25412 8452
rect 25406 8440 25412 8443
rect 25464 8440 25470 8492
rect 25866 8440 25872 8492
rect 25924 8480 25930 8492
rect 31938 8480 31944 8492
rect 25924 8452 31944 8480
rect 25924 8440 25930 8452
rect 31938 8440 31944 8452
rect 31996 8440 32002 8492
rect 32122 8440 32128 8492
rect 32180 8480 32186 8492
rect 32401 8483 32459 8489
rect 32401 8480 32413 8483
rect 32180 8452 32413 8480
rect 32180 8440 32186 8452
rect 32401 8449 32413 8452
rect 32447 8480 32459 8483
rect 32447 8452 32812 8480
rect 32447 8449 32459 8452
rect 32401 8443 32459 8449
rect 32784 8424 32812 8452
rect 33318 8440 33324 8492
rect 33376 8440 33382 8492
rect 22060 8384 22692 8412
rect 22060 8372 22066 8384
rect 31754 8372 31760 8424
rect 31812 8412 31818 8424
rect 32309 8415 32367 8421
rect 32309 8412 32321 8415
rect 31812 8384 32321 8412
rect 31812 8372 31818 8384
rect 32309 8381 32321 8384
rect 32355 8412 32367 8415
rect 32490 8412 32496 8424
rect 32355 8384 32496 8412
rect 32355 8381 32367 8384
rect 32309 8375 32367 8381
rect 32490 8372 32496 8384
rect 32548 8372 32554 8424
rect 32766 8372 32772 8424
rect 32824 8412 32830 8424
rect 33704 8412 33732 8520
rect 35434 8440 35440 8492
rect 35492 8440 35498 8492
rect 35544 8489 35572 8520
rect 35894 8508 35900 8520
rect 35952 8508 35958 8560
rect 35986 8508 35992 8560
rect 36044 8548 36050 8560
rect 36449 8551 36507 8557
rect 36044 8520 36400 8548
rect 36044 8508 36050 8520
rect 35529 8483 35587 8489
rect 35529 8449 35541 8483
rect 35575 8449 35587 8483
rect 35529 8443 35587 8449
rect 35621 8483 35679 8489
rect 35621 8449 35633 8483
rect 35667 8480 35679 8483
rect 35710 8480 35716 8492
rect 35667 8452 35716 8480
rect 35667 8449 35679 8452
rect 35621 8443 35679 8449
rect 35710 8440 35716 8452
rect 35768 8440 35774 8492
rect 35805 8483 35863 8489
rect 35805 8449 35817 8483
rect 35851 8480 35863 8483
rect 36265 8483 36323 8489
rect 36265 8480 36277 8483
rect 35851 8452 36277 8480
rect 35851 8449 35863 8452
rect 35805 8443 35863 8449
rect 36265 8449 36277 8452
rect 36311 8449 36323 8483
rect 36372 8480 36400 8520
rect 36449 8517 36461 8551
rect 36495 8548 36507 8551
rect 37734 8548 37740 8560
rect 36495 8520 37740 8548
rect 36495 8517 36507 8520
rect 36449 8511 36507 8517
rect 37734 8508 37740 8520
rect 37792 8508 37798 8560
rect 36541 8483 36599 8489
rect 36541 8480 36553 8483
rect 36372 8452 36553 8480
rect 36265 8443 36323 8449
rect 36541 8449 36553 8452
rect 36587 8449 36599 8483
rect 36541 8443 36599 8449
rect 35820 8412 35848 8443
rect 36630 8440 36636 8492
rect 36688 8440 36694 8492
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 32824 8384 33732 8412
rect 33888 8384 35848 8412
rect 32824 8372 32830 8384
rect 22094 8344 22100 8356
rect 21376 8316 22100 8344
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 26326 8304 26332 8356
rect 26384 8344 26390 8356
rect 26513 8347 26571 8353
rect 26513 8344 26525 8347
rect 26384 8316 26525 8344
rect 26384 8304 26390 8316
rect 26513 8313 26525 8316
rect 26559 8313 26571 8347
rect 32508 8344 32536 8372
rect 33888 8344 33916 8384
rect 35894 8372 35900 8424
rect 35952 8412 35958 8424
rect 36170 8412 36176 8424
rect 35952 8384 36176 8412
rect 35952 8372 35958 8384
rect 36170 8372 36176 8384
rect 36228 8412 36234 8424
rect 36722 8412 36728 8424
rect 36228 8384 36728 8412
rect 36228 8372 36234 8384
rect 36722 8372 36728 8384
rect 36780 8372 36786 8424
rect 37461 8415 37519 8421
rect 37461 8381 37473 8415
rect 37507 8412 37519 8415
rect 37550 8412 37556 8424
rect 37507 8384 37556 8412
rect 37507 8381 37519 8384
rect 37461 8375 37519 8381
rect 37550 8372 37556 8384
rect 37608 8372 37614 8424
rect 32508 8316 33916 8344
rect 26513 8307 26571 8313
rect 33888 8288 33916 8316
rect 36817 8347 36875 8353
rect 36817 8313 36829 8347
rect 36863 8344 36875 8347
rect 37660 8344 37688 8443
rect 38028 8424 38056 8588
rect 39482 8576 39488 8628
rect 39540 8576 39546 8628
rect 43438 8616 43444 8628
rect 40696 8588 43444 8616
rect 39301 8551 39359 8557
rect 39301 8517 39313 8551
rect 39347 8548 39359 8551
rect 40402 8548 40408 8560
rect 39347 8520 40408 8548
rect 39347 8517 39359 8520
rect 39301 8511 39359 8517
rect 40402 8508 40408 8520
rect 40460 8508 40466 8560
rect 38838 8440 38844 8492
rect 38896 8480 38902 8492
rect 39577 8483 39635 8489
rect 39577 8480 39589 8483
rect 38896 8452 39589 8480
rect 38896 8440 38902 8452
rect 39577 8449 39589 8452
rect 39623 8449 39635 8483
rect 40221 8483 40279 8489
rect 40221 8480 40233 8483
rect 39577 8443 39635 8449
rect 39960 8452 40233 8480
rect 38010 8372 38016 8424
rect 38068 8412 38074 8424
rect 39960 8412 39988 8452
rect 40221 8449 40233 8452
rect 40267 8480 40279 8483
rect 40696 8480 40724 8588
rect 43438 8576 43444 8588
rect 43496 8576 43502 8628
rect 40770 8508 40776 8560
rect 40828 8548 40834 8560
rect 40828 8520 41092 8548
rect 40828 8508 40834 8520
rect 40267 8452 40724 8480
rect 40267 8449 40279 8452
rect 40221 8443 40279 8449
rect 40862 8440 40868 8492
rect 40920 8440 40926 8492
rect 41064 8489 41092 8520
rect 41049 8483 41107 8489
rect 41049 8449 41061 8483
rect 41095 8449 41107 8483
rect 41049 8443 41107 8449
rect 38068 8384 39988 8412
rect 38068 8372 38074 8384
rect 40034 8372 40040 8424
rect 40092 8372 40098 8424
rect 40126 8372 40132 8424
rect 40184 8412 40190 8424
rect 40405 8415 40463 8421
rect 40405 8412 40417 8415
rect 40184 8384 40417 8412
rect 40184 8372 40190 8384
rect 40405 8381 40417 8384
rect 40451 8381 40463 8415
rect 40405 8375 40463 8381
rect 40957 8415 41015 8421
rect 40957 8381 40969 8415
rect 41003 8412 41015 8415
rect 41506 8412 41512 8424
rect 41003 8384 41512 8412
rect 41003 8381 41015 8384
rect 40957 8375 41015 8381
rect 41506 8372 41512 8384
rect 41564 8372 41570 8424
rect 36863 8316 37688 8344
rect 39301 8347 39359 8353
rect 36863 8313 36875 8316
rect 36817 8307 36875 8313
rect 39301 8313 39313 8347
rect 39347 8344 39359 8347
rect 40678 8344 40684 8356
rect 39347 8316 40684 8344
rect 39347 8313 39359 8316
rect 39301 8307 39359 8313
rect 40678 8304 40684 8316
rect 40736 8304 40742 8356
rect 21634 8276 21640 8288
rect 21008 8248 21640 8276
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 25774 8276 25780 8288
rect 22244 8248 25780 8276
rect 22244 8236 22250 8248
rect 25774 8236 25780 8248
rect 25832 8236 25838 8288
rect 33870 8236 33876 8288
rect 33928 8236 33934 8288
rect 35161 8279 35219 8285
rect 35161 8245 35173 8279
rect 35207 8276 35219 8279
rect 35342 8276 35348 8288
rect 35207 8248 35348 8276
rect 35207 8245 35219 8248
rect 35161 8239 35219 8245
rect 35342 8236 35348 8248
rect 35400 8236 35406 8288
rect 37826 8236 37832 8288
rect 37884 8236 37890 8288
rect 40586 8236 40592 8288
rect 40644 8276 40650 8288
rect 54110 8276 54116 8288
rect 40644 8248 54116 8276
rect 40644 8236 40650 8248
rect 54110 8236 54116 8248
rect 54168 8236 54174 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 3053 8075 3111 8081
rect 3053 8072 3065 8075
rect 2372 8044 3065 8072
rect 2372 8032 2378 8044
rect 3053 8041 3065 8044
rect 3099 8072 3111 8075
rect 5074 8072 5080 8084
rect 3099 8044 5080 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 5224 8044 5365 8072
rect 5224 8032 5230 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10962 8072 10968 8084
rect 10008 8044 10968 8072
rect 10008 8032 10014 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12342 8072 12348 8084
rect 11112 8044 12348 8072
rect 11112 8032 11118 8044
rect 12342 8032 12348 8044
rect 12400 8072 12406 8084
rect 15010 8072 15016 8084
rect 12400 8044 15016 8072
rect 12400 8032 12406 8044
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 16540 8044 18337 8072
rect 16540 8032 16546 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 20714 8072 20720 8084
rect 18325 8035 18383 8041
rect 19444 8044 20720 8072
rect 10226 7964 10232 8016
rect 10284 7964 10290 8016
rect 10594 7964 10600 8016
rect 10652 8004 10658 8016
rect 13538 8004 13544 8016
rect 10652 7976 13544 8004
rect 10652 7964 10658 7976
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 14274 8004 14280 8016
rect 13648 7976 14280 8004
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 1762 7868 1768 7880
rect 1719 7840 1768 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 1762 7828 1768 7840
rect 1820 7868 1826 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 1820 7840 3985 7868
rect 1820 7828 1826 7840
rect 3973 7837 3985 7840
rect 4019 7868 4031 7871
rect 4614 7868 4620 7880
rect 4019 7840 4620 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7248 7840 8033 7868
rect 7248 7828 7254 7840
rect 8021 7837 8033 7840
rect 8067 7868 8079 7871
rect 8110 7868 8116 7880
rect 8067 7840 8116 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 10042 7868 10048 7880
rect 8251 7840 10048 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10244 7868 10272 7964
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 11606 7936 11612 7948
rect 11204 7908 11612 7936
rect 11204 7896 11210 7908
rect 11606 7896 11612 7908
rect 11664 7936 11670 7948
rect 13648 7945 13676 7976
rect 14274 7964 14280 7976
rect 14332 7964 14338 8016
rect 17770 7964 17776 8016
rect 17828 8004 17834 8016
rect 19444 8004 19472 8044
rect 20714 8032 20720 8044
rect 20772 8072 20778 8084
rect 21174 8072 21180 8084
rect 20772 8044 21180 8072
rect 20772 8032 20778 8044
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 21634 8032 21640 8084
rect 21692 8032 21698 8084
rect 22373 8075 22431 8081
rect 22373 8041 22385 8075
rect 22419 8072 22431 8075
rect 22738 8072 22744 8084
rect 22419 8044 22744 8072
rect 22419 8041 22431 8044
rect 22373 8035 22431 8041
rect 22738 8032 22744 8044
rect 22796 8032 22802 8084
rect 26234 8072 26240 8084
rect 23676 8044 26240 8072
rect 17828 7976 19472 8004
rect 17828 7964 17834 7976
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 11664 7908 13645 7936
rect 11664 7896 11670 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14918 7936 14924 7948
rect 14056 7908 14924 7936
rect 14056 7896 14062 7908
rect 10962 7868 10968 7880
rect 10244 7840 10968 7868
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 14182 7868 14188 7880
rect 13587 7840 14188 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14384 7877 14412 7908
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 19426 7936 19432 7948
rect 17920 7908 19432 7936
rect 17920 7896 17926 7908
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 21192 7936 21220 8032
rect 22554 7964 22560 8016
rect 22612 8004 22618 8016
rect 23293 8007 23351 8013
rect 23293 8004 23305 8007
rect 22612 7976 23305 8004
rect 22612 7964 22618 7976
rect 23293 7973 23305 7976
rect 23339 7973 23351 8007
rect 23293 7967 23351 7973
rect 23676 7945 23704 8044
rect 26234 8032 26240 8044
rect 26292 8072 26298 8084
rect 27249 8075 27307 8081
rect 27249 8072 27261 8075
rect 26292 8044 27261 8072
rect 26292 8032 26298 8044
rect 27249 8041 27261 8044
rect 27295 8041 27307 8075
rect 27249 8035 27307 8041
rect 27338 8032 27344 8084
rect 27396 8072 27402 8084
rect 40586 8072 40592 8084
rect 27396 8044 40592 8072
rect 27396 8032 27402 8044
rect 40586 8032 40592 8044
rect 40644 8032 40650 8084
rect 30742 7964 30748 8016
rect 30800 8004 30806 8016
rect 31757 8007 31815 8013
rect 31757 8004 31769 8007
rect 30800 7976 31769 8004
rect 30800 7964 30806 7976
rect 31757 7973 31769 7976
rect 31803 7973 31815 8007
rect 33226 8004 33232 8016
rect 31757 7967 31815 7973
rect 32324 7976 33232 8004
rect 23569 7939 23627 7945
rect 23569 7936 23581 7939
rect 21192 7908 23581 7936
rect 23569 7905 23581 7908
rect 23615 7905 23627 7939
rect 23569 7899 23627 7905
rect 23661 7939 23719 7945
rect 23661 7905 23673 7939
rect 23707 7905 23719 7939
rect 23661 7899 23719 7905
rect 25866 7896 25872 7948
rect 25924 7896 25930 7948
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15286 7868 15292 7880
rect 14599 7840 15292 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 1946 7809 1952 7812
rect 1940 7763 1952 7809
rect 1946 7760 1952 7763
rect 2004 7760 2010 7812
rect 4240 7803 4298 7809
rect 4240 7769 4252 7803
rect 4286 7800 4298 7803
rect 4522 7800 4528 7812
rect 4286 7772 4528 7800
rect 4286 7769 4298 7772
rect 4240 7763 4298 7769
rect 4522 7760 4528 7772
rect 4580 7760 4586 7812
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7742 7800 7748 7812
rect 7156 7772 7748 7800
rect 7156 7760 7162 7772
rect 7742 7760 7748 7772
rect 7800 7800 7806 7812
rect 7837 7803 7895 7809
rect 7837 7800 7849 7803
rect 7800 7772 7849 7800
rect 7800 7760 7806 7772
rect 7837 7769 7849 7772
rect 7883 7769 7895 7803
rect 7837 7763 7895 7769
rect 11238 7760 11244 7812
rect 11296 7800 11302 7812
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 11296 7772 14473 7800
rect 11296 7760 11302 7772
rect 14461 7769 14473 7772
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 8846 7732 8852 7744
rect 4764 7704 8852 7732
rect 4764 7692 4770 7704
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 11204 7704 13185 7732
rect 11204 7692 11210 7704
rect 13173 7701 13185 7704
rect 13219 7701 13231 7735
rect 13173 7695 13231 7701
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14568 7732 14596 7831
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 18509 7871 18567 7877
rect 18509 7868 18521 7871
rect 18380 7840 18521 7868
rect 18380 7828 18386 7840
rect 18509 7837 18521 7840
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 19334 7868 19340 7880
rect 18831 7840 19340 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 15013 7803 15071 7809
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 15746 7800 15752 7812
rect 15059 7772 15752 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15746 7760 15752 7772
rect 15804 7800 15810 7812
rect 17402 7800 17408 7812
rect 15804 7772 17408 7800
rect 15804 7760 15810 7772
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 18616 7800 18644 7831
rect 17828 7772 18644 7800
rect 17828 7760 17834 7772
rect 14148 7704 14596 7732
rect 18708 7732 18736 7831
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 22554 7868 22560 7880
rect 20036 7840 22560 7868
rect 20036 7828 20042 7840
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 23106 7868 23112 7880
rect 22879 7840 23112 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 23106 7828 23112 7840
rect 23164 7828 23170 7880
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 26142 7877 26148 7880
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7837 23811 7871
rect 26136 7868 26148 7877
rect 26103 7840 26148 7868
rect 23753 7831 23811 7837
rect 26136 7831 26148 7840
rect 19150 7760 19156 7812
rect 19208 7800 19214 7812
rect 19674 7803 19732 7809
rect 19674 7800 19686 7803
rect 19208 7772 19686 7800
rect 19208 7760 19214 7772
rect 19674 7769 19686 7772
rect 19720 7769 19732 7803
rect 19674 7763 19732 7769
rect 20898 7760 20904 7812
rect 20956 7800 20962 7812
rect 21361 7803 21419 7809
rect 21361 7800 21373 7803
rect 20956 7772 21373 7800
rect 20956 7760 20962 7772
rect 21361 7769 21373 7772
rect 21407 7769 21419 7803
rect 21361 7763 21419 7769
rect 22741 7803 22799 7809
rect 22741 7769 22753 7803
rect 22787 7800 22799 7803
rect 22922 7800 22928 7812
rect 22787 7772 22928 7800
rect 22787 7769 22799 7772
rect 22741 7763 22799 7769
rect 22922 7760 22928 7772
rect 22980 7760 22986 7812
rect 20806 7732 20812 7744
rect 18708 7704 20812 7732
rect 14148 7692 14154 7704
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 23768 7732 23796 7831
rect 26142 7828 26148 7831
rect 26200 7828 26206 7880
rect 31570 7828 31576 7880
rect 31628 7828 31634 7880
rect 31662 7828 31668 7880
rect 31720 7868 31726 7880
rect 32324 7877 32352 7976
rect 33226 7964 33232 7976
rect 33284 8004 33290 8016
rect 33594 8004 33600 8016
rect 33284 7976 33600 8004
rect 33284 7964 33290 7976
rect 33594 7964 33600 7976
rect 33652 7964 33658 8016
rect 35176 7976 35940 8004
rect 32398 7896 32404 7948
rect 32456 7896 32462 7948
rect 32858 7896 32864 7948
rect 32916 7936 32922 7948
rect 35176 7945 35204 7976
rect 35161 7939 35219 7945
rect 35161 7936 35173 7939
rect 32916 7908 35173 7936
rect 32916 7896 32922 7908
rect 35161 7905 35173 7908
rect 35207 7905 35219 7939
rect 35161 7899 35219 7905
rect 35342 7896 35348 7948
rect 35400 7896 35406 7948
rect 32309 7871 32367 7877
rect 31720 7828 31754 7868
rect 32309 7837 32321 7871
rect 32355 7837 32367 7871
rect 32416 7868 32444 7896
rect 32585 7871 32643 7877
rect 32585 7868 32597 7871
rect 32416 7840 32597 7868
rect 32309 7831 32367 7837
rect 32585 7837 32597 7840
rect 32631 7837 32643 7871
rect 32585 7831 32643 7837
rect 32677 7871 32735 7877
rect 32677 7837 32689 7871
rect 32723 7868 32735 7871
rect 33042 7868 33048 7880
rect 32723 7840 33048 7868
rect 32723 7837 32735 7840
rect 32677 7831 32735 7837
rect 22152 7704 23796 7732
rect 31726 7732 31754 7828
rect 32398 7760 32404 7812
rect 32456 7800 32462 7812
rect 32493 7803 32551 7809
rect 32493 7800 32505 7803
rect 32456 7772 32505 7800
rect 32456 7760 32462 7772
rect 32493 7769 32505 7772
rect 32539 7769 32551 7803
rect 32493 7763 32551 7769
rect 32692 7732 32720 7831
rect 33042 7828 33048 7840
rect 33100 7828 33106 7880
rect 33134 7828 33140 7880
rect 33192 7868 33198 7880
rect 33321 7871 33379 7877
rect 33321 7868 33333 7871
rect 33192 7840 33333 7868
rect 33192 7828 33198 7840
rect 33321 7837 33333 7840
rect 33367 7868 33379 7871
rect 34054 7868 34060 7880
rect 33367 7840 34060 7868
rect 33367 7837 33379 7840
rect 33321 7831 33379 7837
rect 34054 7828 34060 7840
rect 34112 7828 34118 7880
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 35069 7871 35127 7877
rect 35069 7868 35081 7871
rect 34848 7840 35081 7868
rect 34848 7828 34854 7840
rect 35069 7837 35081 7840
rect 35115 7837 35127 7871
rect 35069 7831 35127 7837
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7837 35311 7871
rect 35253 7831 35311 7837
rect 33226 7760 33232 7812
rect 33284 7800 33290 7812
rect 33597 7803 33655 7809
rect 33597 7800 33609 7803
rect 33284 7772 33609 7800
rect 33284 7760 33290 7772
rect 33597 7769 33609 7772
rect 33643 7769 33655 7803
rect 33597 7763 33655 7769
rect 33778 7760 33784 7812
rect 33836 7800 33842 7812
rect 35268 7800 35296 7831
rect 33836 7772 35296 7800
rect 35912 7800 35940 7976
rect 40310 7896 40316 7948
rect 40368 7936 40374 7948
rect 40368 7908 40448 7936
rect 40368 7896 40374 7908
rect 35986 7828 35992 7880
rect 36044 7828 36050 7880
rect 36256 7871 36314 7877
rect 36256 7837 36268 7871
rect 36302 7868 36314 7871
rect 37826 7868 37832 7880
rect 36302 7840 37832 7868
rect 36302 7837 36314 7840
rect 36256 7831 36314 7837
rect 37826 7828 37832 7840
rect 37884 7828 37890 7880
rect 40034 7828 40040 7880
rect 40092 7828 40098 7880
rect 40420 7877 40448 7908
rect 40405 7871 40463 7877
rect 40405 7837 40417 7871
rect 40451 7837 40463 7871
rect 40405 7831 40463 7837
rect 41046 7828 41052 7880
rect 41104 7868 41110 7880
rect 41506 7877 41512 7880
rect 41233 7871 41291 7877
rect 41233 7868 41245 7871
rect 41104 7840 41245 7868
rect 41104 7828 41110 7840
rect 41233 7837 41245 7840
rect 41279 7837 41291 7871
rect 41233 7831 41291 7837
rect 41500 7831 41512 7877
rect 41506 7828 41512 7831
rect 41564 7828 41570 7880
rect 40126 7800 40132 7812
rect 35912 7772 40132 7800
rect 33836 7760 33842 7772
rect 40126 7760 40132 7772
rect 40184 7760 40190 7812
rect 40218 7760 40224 7812
rect 40276 7760 40282 7812
rect 40313 7803 40371 7809
rect 40313 7769 40325 7803
rect 40359 7800 40371 7803
rect 40359 7772 42656 7800
rect 40359 7769 40371 7772
rect 40313 7763 40371 7769
rect 31726 7704 32720 7732
rect 32861 7735 32919 7741
rect 22152 7692 22158 7704
rect 32861 7701 32873 7735
rect 32907 7732 32919 7735
rect 33134 7732 33140 7744
rect 32907 7704 33140 7732
rect 32907 7701 32919 7704
rect 32861 7695 32919 7701
rect 33134 7692 33140 7704
rect 33192 7692 33198 7744
rect 33410 7692 33416 7744
rect 33468 7732 33474 7744
rect 34330 7732 34336 7744
rect 33468 7704 34336 7732
rect 33468 7692 33474 7704
rect 34330 7692 34336 7704
rect 34388 7692 34394 7744
rect 34885 7735 34943 7741
rect 34885 7701 34897 7735
rect 34931 7732 34943 7735
rect 35618 7732 35624 7744
rect 34931 7704 35624 7732
rect 34931 7701 34943 7704
rect 34885 7695 34943 7701
rect 35618 7692 35624 7704
rect 35676 7692 35682 7744
rect 37369 7735 37427 7741
rect 37369 7701 37381 7735
rect 37415 7732 37427 7735
rect 38654 7732 38660 7744
rect 37415 7704 38660 7732
rect 37415 7701 37427 7704
rect 37369 7695 37427 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 40402 7692 40408 7744
rect 40460 7732 40466 7744
rect 42628 7741 42656 7772
rect 40589 7735 40647 7741
rect 40589 7732 40601 7735
rect 40460 7704 40601 7732
rect 40460 7692 40466 7704
rect 40589 7701 40601 7704
rect 40635 7701 40647 7735
rect 40589 7695 40647 7701
rect 42613 7735 42671 7741
rect 42613 7701 42625 7735
rect 42659 7732 42671 7735
rect 43254 7732 43260 7744
rect 42659 7704 43260 7732
rect 42659 7701 42671 7704
rect 42613 7695 42671 7701
rect 43254 7692 43260 7704
rect 43312 7692 43318 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 1946 7488 1952 7540
rect 2004 7488 2010 7540
rect 2314 7488 2320 7540
rect 2372 7488 2378 7540
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 2455 7500 3341 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 4522 7488 4528 7540
rect 4580 7488 4586 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5166 7528 5172 7540
rect 4939 7500 5172 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9766 7528 9772 7540
rect 9447 7500 9772 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 13412 7500 14841 7528
rect 13412 7488 13418 7500
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 14829 7491 14887 7497
rect 19150 7488 19156 7540
rect 19208 7488 19214 7540
rect 19521 7531 19579 7537
rect 19521 7497 19533 7531
rect 19567 7528 19579 7531
rect 20806 7528 20812 7540
rect 19567 7500 20812 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 27338 7528 27344 7540
rect 22066 7500 27344 7528
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 3237 7463 3295 7469
rect 3237 7460 3249 7463
rect 992 7432 3249 7460
rect 992 7420 998 7432
rect 3237 7429 3249 7432
rect 3283 7429 3295 7463
rect 11146 7460 11152 7472
rect 3237 7423 3295 7429
rect 4724 7432 11152 7460
rect 4724 7401 4752 7432
rect 11146 7420 11152 7432
rect 11204 7420 11210 7472
rect 11698 7420 11704 7472
rect 11756 7420 11762 7472
rect 11917 7463 11975 7469
rect 11917 7429 11929 7463
rect 11963 7460 11975 7463
rect 14090 7460 14096 7472
rect 11963 7432 14096 7460
rect 11963 7429 11975 7432
rect 11917 7423 11975 7429
rect 14090 7420 14096 7432
rect 14148 7420 14154 7472
rect 17770 7460 17776 7472
rect 15120 7432 17776 7460
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5718 7392 5724 7404
rect 5031 7364 5724 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7392 7067 7395
rect 7190 7392 7196 7404
rect 7055 7364 7196 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 10318 7392 10324 7404
rect 9355 7364 10324 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10686 7352 10692 7404
rect 10744 7352 10750 7404
rect 12406 7364 14964 7392
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 2464 7296 2513 7324
rect 2464 7284 2470 7296
rect 2501 7293 2513 7296
rect 2547 7324 2559 7327
rect 2590 7324 2596 7336
rect 2547 7296 2596 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 7098 7284 7104 7336
rect 7156 7284 7162 7336
rect 9582 7284 9588 7336
rect 9640 7284 9646 7336
rect 10870 7284 10876 7336
rect 10928 7284 10934 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 12066 7324 12072 7336
rect 11112 7296 12072 7324
rect 11112 7284 11118 7296
rect 12066 7284 12072 7296
rect 12124 7324 12130 7336
rect 12406 7324 12434 7364
rect 12124 7296 12434 7324
rect 14936 7324 14964 7364
rect 15010 7352 15016 7404
rect 15068 7352 15074 7404
rect 15120 7333 15148 7432
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 20254 7420 20260 7472
rect 20312 7460 20318 7472
rect 22066 7460 22094 7500
rect 27338 7488 27344 7500
rect 27396 7488 27402 7540
rect 32398 7488 32404 7540
rect 32456 7488 32462 7540
rect 32508 7500 32720 7528
rect 20312 7432 22094 7460
rect 20312 7420 20318 7432
rect 22554 7420 22560 7472
rect 22612 7460 22618 7472
rect 32508 7460 32536 7500
rect 22612 7432 32536 7460
rect 32692 7460 32720 7500
rect 33318 7488 33324 7540
rect 33376 7528 33382 7540
rect 33505 7531 33563 7537
rect 33505 7528 33517 7531
rect 33376 7500 33517 7528
rect 33376 7488 33382 7500
rect 33505 7497 33517 7500
rect 33551 7497 33563 7531
rect 33505 7491 33563 7497
rect 37734 7488 37740 7540
rect 37792 7488 37798 7540
rect 42610 7460 42616 7472
rect 32692 7432 42616 7460
rect 22612 7420 22618 7432
rect 42610 7420 42616 7432
rect 42668 7420 42674 7472
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 16666 7392 16672 7404
rect 15243 7364 16672 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 19610 7352 19616 7404
rect 19668 7392 19674 7404
rect 20070 7392 20076 7404
rect 19668 7364 20076 7392
rect 19668 7352 19674 7364
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 24670 7392 24676 7404
rect 22971 7364 24676 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 30374 7352 30380 7404
rect 30432 7392 30438 7404
rect 31294 7392 31300 7404
rect 30432 7364 31300 7392
rect 30432 7352 30438 7364
rect 31294 7352 31300 7364
rect 31352 7392 31358 7404
rect 32398 7392 32404 7404
rect 31352 7364 32404 7392
rect 31352 7352 31358 7364
rect 32398 7352 32404 7364
rect 32456 7392 32462 7404
rect 32585 7395 32643 7401
rect 32585 7392 32597 7395
rect 32456 7364 32597 7392
rect 32456 7352 32462 7364
rect 32585 7361 32597 7364
rect 32631 7361 32643 7395
rect 32585 7355 32643 7361
rect 32674 7352 32680 7404
rect 32732 7352 32738 7404
rect 32953 7395 33011 7401
rect 32953 7361 32965 7395
rect 32999 7361 33011 7395
rect 32953 7355 33011 7361
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14936 7296 15117 7324
rect 12124 7284 12130 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7324 15347 7327
rect 17034 7324 17040 7336
rect 15335 7296 17040 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 23014 7284 23020 7336
rect 23072 7284 23078 7336
rect 23106 7284 23112 7336
rect 23164 7284 23170 7336
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7293 23259 7327
rect 23201 7287 23259 7293
rect 17218 7256 17224 7268
rect 11900 7228 17224 7256
rect 7282 7148 7288 7200
rect 7340 7148 7346 7200
rect 8938 7148 8944 7200
rect 8996 7148 9002 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10502 7188 10508 7200
rect 10284 7160 10508 7188
rect 10284 7148 10290 7160
rect 10502 7148 10508 7160
rect 10560 7188 10566 7200
rect 11900 7197 11928 7228
rect 17218 7216 17224 7228
rect 17276 7216 17282 7268
rect 23216 7256 23244 7287
rect 30834 7284 30840 7336
rect 30892 7324 30898 7336
rect 32858 7324 32864 7336
rect 30892 7296 32864 7324
rect 30892 7284 30898 7296
rect 32858 7284 32864 7296
rect 32916 7284 32922 7336
rect 32968 7324 32996 7355
rect 33410 7352 33416 7404
rect 33468 7352 33474 7404
rect 33597 7395 33655 7401
rect 33597 7361 33609 7395
rect 33643 7392 33655 7395
rect 33870 7392 33876 7404
rect 33643 7364 33876 7392
rect 33643 7361 33655 7364
rect 33597 7355 33655 7361
rect 33870 7352 33876 7364
rect 33928 7392 33934 7404
rect 34330 7392 34336 7404
rect 33928 7364 34336 7392
rect 33928 7352 33934 7364
rect 34330 7352 34336 7364
rect 34388 7352 34394 7404
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7392 38163 7395
rect 38654 7392 38660 7404
rect 38151 7364 38660 7392
rect 38151 7361 38163 7364
rect 38105 7355 38163 7361
rect 38654 7352 38660 7364
rect 38712 7392 38718 7404
rect 39206 7392 39212 7404
rect 38712 7364 39212 7392
rect 38712 7352 38718 7364
rect 39206 7352 39212 7364
rect 39264 7352 39270 7404
rect 42794 7352 42800 7404
rect 42852 7352 42858 7404
rect 33686 7324 33692 7336
rect 32968 7296 33692 7324
rect 33686 7284 33692 7296
rect 33744 7284 33750 7336
rect 38194 7284 38200 7336
rect 38252 7284 38258 7336
rect 38378 7284 38384 7336
rect 38436 7284 38442 7336
rect 41690 7284 41696 7336
rect 41748 7324 41754 7336
rect 42613 7327 42671 7333
rect 42613 7324 42625 7327
rect 41748 7296 42625 7324
rect 41748 7284 41754 7296
rect 42613 7293 42625 7296
rect 42659 7293 42671 7327
rect 42613 7287 42671 7293
rect 33042 7256 33048 7268
rect 22066 7228 33048 7256
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 10560 7160 11897 7188
rect 10560 7148 10566 7160
rect 11885 7157 11897 7160
rect 11931 7157 11943 7191
rect 11885 7151 11943 7157
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 12032 7160 12081 7188
rect 12032 7148 12038 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 22066 7188 22094 7228
rect 33042 7216 33048 7228
rect 33100 7216 33106 7268
rect 33226 7216 33232 7268
rect 33284 7256 33290 7268
rect 39022 7256 39028 7268
rect 33284 7228 39028 7256
rect 33284 7216 33290 7228
rect 39022 7216 39028 7228
rect 39080 7256 39086 7268
rect 40218 7256 40224 7268
rect 39080 7228 40224 7256
rect 39080 7216 39086 7228
rect 40218 7216 40224 7228
rect 40276 7216 40282 7268
rect 14608 7160 22094 7188
rect 14608 7148 14614 7160
rect 22738 7148 22744 7200
rect 22796 7148 22802 7200
rect 32030 7148 32036 7200
rect 32088 7188 32094 7200
rect 32766 7188 32772 7200
rect 32088 7160 32772 7188
rect 32088 7148 32094 7160
rect 32766 7148 32772 7160
rect 32824 7188 32830 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32824 7160 32873 7188
rect 32824 7148 32830 7160
rect 32861 7157 32873 7160
rect 32907 7157 32919 7191
rect 32861 7151 32919 7157
rect 32950 7148 32956 7200
rect 33008 7188 33014 7200
rect 33410 7188 33416 7200
rect 33008 7160 33416 7188
rect 33008 7148 33014 7160
rect 33410 7148 33416 7160
rect 33468 7148 33474 7200
rect 42978 7148 42984 7200
rect 43036 7148 43042 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13446 6984 13452 6996
rect 12492 6956 13452 6984
rect 12492 6944 12498 6956
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 16666 6944 16672 6996
rect 16724 6944 16730 6996
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 33778 6984 33784 6996
rect 17276 6956 33784 6984
rect 17276 6944 17282 6956
rect 33778 6944 33784 6956
rect 33836 6944 33842 6996
rect 11054 6916 11060 6928
rect 10796 6888 11060 6916
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 2685 6851 2743 6857
rect 2685 6848 2697 6851
rect 2648 6820 2697 6848
rect 2648 6808 2654 6820
rect 2685 6817 2697 6820
rect 2731 6817 2743 6851
rect 2685 6811 2743 6817
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4798 6848 4804 6860
rect 4295 6820 4804 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 10796 6848 10824 6888
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 32858 6916 32864 6928
rect 31588 6888 32864 6916
rect 8444 6820 10824 6848
rect 8444 6808 8450 6820
rect 10870 6808 10876 6860
rect 10928 6808 10934 6860
rect 22002 6808 22008 6860
rect 22060 6808 22066 6860
rect 24670 6808 24676 6860
rect 24728 6808 24734 6860
rect 30006 6808 30012 6860
rect 30064 6848 30070 6860
rect 30929 6851 30987 6857
rect 30929 6848 30941 6851
rect 30064 6820 30941 6848
rect 30064 6808 30070 6820
rect 30929 6817 30941 6820
rect 30975 6817 30987 6851
rect 30929 6811 30987 6817
rect 31297 6851 31355 6857
rect 31297 6817 31309 6851
rect 31343 6848 31355 6851
rect 31588 6848 31616 6888
rect 32858 6876 32864 6888
rect 32916 6876 32922 6928
rect 31754 6848 31760 6860
rect 31343 6820 31616 6848
rect 31680 6820 31760 6848
rect 31343 6817 31355 6820
rect 31297 6811 31355 6817
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 992 6752 4077 6780
rect 992 6740 998 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 8076 6752 8125 6780
rect 8076 6740 8082 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 10888 6780 10916 6808
rect 10183 6752 10916 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 13446 6780 13452 6792
rect 11572 6752 13452 6780
rect 11572 6740 11578 6752
rect 13446 6740 13452 6752
rect 13504 6780 13510 6792
rect 15102 6780 15108 6792
rect 13504 6752 15108 6780
rect 13504 6740 13510 6752
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15160 6752 15301 6780
rect 15160 6740 15166 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6780 17371 6783
rect 17402 6780 17408 6792
rect 17359 6752 17408 6780
rect 17359 6749 17371 6752
rect 17313 6743 17371 6749
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17552 6752 17601 6780
rect 17552 6740 17558 6752
rect 17589 6749 17601 6752
rect 17635 6780 17647 6783
rect 19242 6780 19248 6792
rect 17635 6752 19248 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 19242 6740 19248 6752
rect 19300 6780 19306 6792
rect 19610 6780 19616 6792
rect 19300 6752 19616 6780
rect 19300 6740 19306 6752
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 22272 6783 22330 6789
rect 22272 6749 22284 6783
rect 22318 6780 22330 6783
rect 22738 6780 22744 6792
rect 22318 6752 22744 6780
rect 22318 6749 22330 6752
rect 22272 6743 22330 6749
rect 22738 6740 22744 6752
rect 22796 6740 22802 6792
rect 24486 6740 24492 6792
rect 24544 6780 24550 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 24544 6752 24593 6780
rect 24544 6740 24550 6752
rect 24581 6749 24593 6752
rect 24627 6780 24639 6783
rect 26418 6780 26424 6792
rect 24627 6752 26424 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 29328 6752 29745 6780
rect 29328 6740 29334 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 29914 6740 29920 6792
rect 29972 6740 29978 6792
rect 30098 6740 30104 6792
rect 30156 6740 30162 6792
rect 30282 6740 30288 6792
rect 30340 6740 30346 6792
rect 30834 6740 30840 6792
rect 30892 6780 30898 6792
rect 31113 6783 31171 6789
rect 31113 6780 31125 6783
rect 30892 6752 31125 6780
rect 30892 6740 30898 6752
rect 31113 6749 31125 6752
rect 31159 6749 31171 6783
rect 31113 6743 31171 6749
rect 31202 6740 31208 6792
rect 31260 6740 31266 6792
rect 31386 6740 31392 6792
rect 31444 6740 31450 6792
rect 31680 6780 31708 6820
rect 31754 6808 31760 6820
rect 31812 6808 31818 6860
rect 31864 6820 32996 6848
rect 31588 6752 31708 6780
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 8389 6715 8447 6721
rect 8389 6712 8401 6715
rect 8352 6684 8401 6712
rect 8352 6672 8358 6684
rect 8389 6681 8401 6684
rect 8435 6712 8447 6715
rect 9030 6712 9036 6724
rect 8435 6684 9036 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 10870 6672 10876 6724
rect 10928 6672 10934 6724
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11606 6712 11612 6724
rect 11112 6684 11612 6712
rect 11112 6672 11118 6684
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 11790 6721 11796 6724
rect 11784 6675 11796 6721
rect 11790 6672 11796 6675
rect 11848 6672 11854 6724
rect 15556 6715 15614 6721
rect 15556 6681 15568 6715
rect 15602 6712 15614 6715
rect 17129 6715 17187 6721
rect 17129 6712 17141 6715
rect 15602 6684 17141 6712
rect 15602 6681 15614 6684
rect 15556 6675 15614 6681
rect 17129 6681 17141 6684
rect 17175 6681 17187 6715
rect 17129 6675 17187 6681
rect 17218 6672 17224 6724
rect 17276 6712 17282 6724
rect 31220 6712 31248 6740
rect 31588 6712 31616 6752
rect 17276 6684 31156 6712
rect 31220 6684 31616 6712
rect 17276 6672 17282 6684
rect 2130 6604 2136 6656
rect 2188 6604 2194 6656
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 2593 6647 2651 6653
rect 2593 6613 2605 6647
rect 2639 6644 2651 6647
rect 3418 6644 3424 6656
rect 2639 6616 3424 6644
rect 2639 6613 2651 6616
rect 2593 6607 2651 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 11698 6644 11704 6656
rect 9916 6616 11704 6644
rect 9916 6604 9922 6616
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12216 6616 12909 6644
rect 12216 6604 12222 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 16724 6616 17509 6644
rect 16724 6604 16730 6616
rect 17497 6613 17509 6616
rect 17543 6613 17555 6647
rect 17497 6607 17555 6613
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 23385 6647 23443 6653
rect 23385 6644 23397 6647
rect 22152 6616 23397 6644
rect 22152 6604 22158 6616
rect 23385 6613 23397 6616
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 30466 6604 30472 6656
rect 30524 6604 30530 6656
rect 31128 6644 31156 6684
rect 31864 6644 31892 6820
rect 32030 6740 32036 6792
rect 32088 6740 32094 6792
rect 32217 6783 32275 6789
rect 32217 6749 32229 6783
rect 32263 6780 32275 6783
rect 32490 6780 32496 6792
rect 32263 6752 32496 6780
rect 32263 6749 32275 6752
rect 32217 6743 32275 6749
rect 32490 6740 32496 6752
rect 32548 6740 32554 6792
rect 32861 6783 32919 6789
rect 32861 6749 32873 6783
rect 32907 6749 32919 6783
rect 32861 6743 32919 6749
rect 32306 6672 32312 6724
rect 32364 6672 32370 6724
rect 31128 6616 31892 6644
rect 31938 6604 31944 6656
rect 31996 6644 32002 6656
rect 32876 6644 32904 6743
rect 32968 6712 32996 6820
rect 35710 6808 35716 6860
rect 35768 6848 35774 6860
rect 36633 6851 36691 6857
rect 36633 6848 36645 6851
rect 35768 6820 36645 6848
rect 35768 6808 35774 6820
rect 36633 6817 36645 6820
rect 36679 6817 36691 6851
rect 36633 6811 36691 6817
rect 44008 6820 44496 6848
rect 33134 6789 33140 6792
rect 33128 6780 33140 6789
rect 33095 6752 33140 6780
rect 33128 6743 33140 6752
rect 33134 6740 33140 6743
rect 33192 6740 33198 6792
rect 35526 6740 35532 6792
rect 35584 6740 35590 6792
rect 35618 6740 35624 6792
rect 35676 6740 35682 6792
rect 35728 6752 38654 6780
rect 35728 6712 35756 6752
rect 32968 6684 35756 6712
rect 36265 6715 36323 6721
rect 36265 6681 36277 6715
rect 36311 6681 36323 6715
rect 36265 6675 36323 6681
rect 31996 6616 32904 6644
rect 34241 6647 34299 6653
rect 31996 6604 32002 6616
rect 34241 6613 34253 6647
rect 34287 6644 34299 6647
rect 34514 6644 34520 6656
rect 34287 6616 34520 6644
rect 34287 6613 34299 6616
rect 34241 6607 34299 6613
rect 34514 6604 34520 6616
rect 34572 6604 34578 6656
rect 35802 6604 35808 6656
rect 35860 6604 35866 6656
rect 36280 6644 36308 6675
rect 36446 6672 36452 6724
rect 36504 6672 36510 6724
rect 36722 6672 36728 6724
rect 36780 6712 36786 6724
rect 38626 6712 38654 6752
rect 41046 6740 41052 6792
rect 41104 6780 41110 6792
rect 41325 6783 41383 6789
rect 41325 6780 41337 6783
rect 41104 6752 41337 6780
rect 41104 6740 41110 6752
rect 41325 6749 41337 6752
rect 41371 6749 41383 6783
rect 41325 6743 41383 6749
rect 41592 6783 41650 6789
rect 41592 6749 41604 6783
rect 41638 6780 41650 6783
rect 42978 6780 42984 6792
rect 41638 6752 42984 6780
rect 41638 6749 41650 6752
rect 41592 6743 41650 6749
rect 42978 6740 42984 6752
rect 43036 6740 43042 6792
rect 44008 6789 44036 6820
rect 43993 6783 44051 6789
rect 43993 6749 44005 6783
rect 44039 6749 44051 6783
rect 43993 6743 44051 6749
rect 44085 6783 44143 6789
rect 44085 6749 44097 6783
rect 44131 6749 44143 6783
rect 44085 6743 44143 6749
rect 44177 6783 44235 6789
rect 44177 6749 44189 6783
rect 44223 6780 44235 6783
rect 44266 6780 44272 6792
rect 44223 6752 44272 6780
rect 44223 6749 44235 6752
rect 44177 6743 44235 6749
rect 42150 6712 42156 6724
rect 36780 6684 38516 6712
rect 38626 6684 42156 6712
rect 36780 6672 36786 6684
rect 36538 6644 36544 6656
rect 36280 6616 36544 6644
rect 36538 6604 36544 6616
rect 36596 6644 36602 6656
rect 38378 6644 38384 6656
rect 36596 6616 38384 6644
rect 36596 6604 36602 6616
rect 38378 6604 38384 6616
rect 38436 6604 38442 6656
rect 38488 6644 38516 6684
rect 42150 6672 42156 6684
rect 42208 6672 42214 6724
rect 44100 6712 44128 6743
rect 44266 6740 44272 6752
rect 44324 6740 44330 6792
rect 44361 6783 44419 6789
rect 44361 6749 44373 6783
rect 44407 6749 44419 6783
rect 44361 6743 44419 6749
rect 44376 6712 44404 6743
rect 42628 6684 44128 6712
rect 44284 6684 44404 6712
rect 42628 6644 42656 6684
rect 38488 6616 42656 6644
rect 42705 6647 42763 6653
rect 42705 6613 42717 6647
rect 42751 6644 42763 6647
rect 42886 6644 42892 6656
rect 42751 6616 42892 6644
rect 42751 6613 42763 6616
rect 42705 6607 42763 6613
rect 42886 6604 42892 6616
rect 42944 6604 42950 6656
rect 43070 6604 43076 6656
rect 43128 6644 43134 6656
rect 43717 6647 43775 6653
rect 43717 6644 43729 6647
rect 43128 6616 43729 6644
rect 43128 6604 43134 6616
rect 43717 6613 43729 6616
rect 43763 6613 43775 6647
rect 43717 6607 43775 6613
rect 43990 6604 43996 6656
rect 44048 6644 44054 6656
rect 44284 6644 44312 6684
rect 44048 6616 44312 6644
rect 44048 6604 44054 6616
rect 44358 6604 44364 6656
rect 44416 6644 44422 6656
rect 44468 6644 44496 6820
rect 44416 6616 44496 6644
rect 44416 6604 44422 6616
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 8386 6440 8392 6452
rect 2556 6412 8392 6440
rect 2556 6400 2562 6412
rect 2130 6381 2136 6384
rect 2124 6335 2136 6381
rect 2130 6332 2136 6335
rect 2188 6332 2194 6384
rect 4080 6381 4108 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 8938 6440 8944 6452
rect 8527 6412 8944 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9088 6412 9904 6440
rect 9088 6400 9094 6412
rect 4065 6375 4123 6381
rect 4065 6341 4077 6375
rect 4111 6341 4123 6375
rect 4065 6335 4123 6341
rect 7282 6332 7288 6384
rect 7340 6332 7346 6384
rect 8018 6332 8024 6384
rect 8076 6372 8082 6384
rect 9876 6372 9904 6412
rect 10318 6400 10324 6452
rect 10376 6400 10382 6452
rect 11054 6440 11060 6452
rect 10428 6412 11060 6440
rect 10428 6372 10456 6412
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 11790 6400 11796 6452
rect 11848 6400 11854 6452
rect 13464 6412 14228 6440
rect 13170 6372 13176 6384
rect 8076 6344 9674 6372
rect 9876 6344 10456 6372
rect 10520 6344 13176 6372
rect 8076 6332 8082 6344
rect 3786 6264 3792 6316
rect 3844 6264 3850 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5810 6304 5816 6316
rect 5399 6276 5816 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 1857 6239 1915 6245
rect 1857 6236 1869 6239
rect 1820 6208 1869 6236
rect 1820 6196 1826 6208
rect 1857 6205 1869 6208
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 3237 6171 3295 6177
rect 3237 6137 3249 6171
rect 3283 6168 3295 6171
rect 3804 6168 3832 6264
rect 5184 6236 5212 6267
rect 5810 6264 5816 6276
rect 5868 6304 5874 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 5868 6276 7481 6304
rect 5868 6264 5874 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 7558 6304 7564 6316
rect 7515 6276 7564 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 7699 6276 9413 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9646 6304 9674 6344
rect 10520 6313 10548 6344
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9646 6276 9781 6304
rect 9401 6267 9459 6273
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 6546 6236 6552 6248
rect 5184 6208 6552 6236
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 8570 6196 8576 6248
rect 8628 6196 8634 6248
rect 8662 6196 8668 6248
rect 8720 6196 8726 6248
rect 9784 6236 9812 6267
rect 10612 6236 10640 6267
rect 10686 6264 10692 6316
rect 10744 6264 10750 6316
rect 10827 6307 10885 6313
rect 10827 6273 10839 6307
rect 10873 6304 10885 6307
rect 11330 6304 11336 6316
rect 10873 6276 11336 6304
rect 10873 6273 10885 6276
rect 10827 6267 10885 6273
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 12158 6264 12164 6316
rect 12216 6264 12222 6316
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6304 12311 6307
rect 13464 6304 13492 6412
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 13998 6372 14004 6384
rect 13955 6344 14004 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 14090 6332 14096 6384
rect 14148 6381 14154 6384
rect 14148 6375 14167 6381
rect 14155 6341 14167 6375
rect 14200 6372 14228 6412
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 34514 6440 34520 6452
rect 17460 6412 33916 6440
rect 17460 6400 17466 6412
rect 14734 6372 14740 6384
rect 14200 6344 14740 6372
rect 14148 6335 14167 6341
rect 14148 6332 14154 6335
rect 14734 6332 14740 6344
rect 14792 6372 14798 6384
rect 17494 6372 17500 6384
rect 14792 6344 17500 6372
rect 14792 6332 14798 6344
rect 17494 6332 17500 6344
rect 17552 6332 17558 6384
rect 22373 6375 22431 6381
rect 22373 6341 22385 6375
rect 22419 6372 22431 6375
rect 26142 6372 26148 6384
rect 22419 6344 26148 6372
rect 22419 6341 22431 6344
rect 22373 6335 22431 6341
rect 26142 6332 26148 6344
rect 26200 6332 26206 6384
rect 29730 6372 29736 6384
rect 28276 6344 29736 6372
rect 12299 6276 13492 6304
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 13596 6276 19349 6304
rect 13596 6264 13602 6276
rect 19337 6273 19349 6276
rect 19383 6304 19395 6307
rect 20438 6304 20444 6316
rect 19383 6276 20444 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 22002 6264 22008 6316
rect 22060 6264 22066 6316
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22554 6313 22560 6316
rect 22281 6307 22339 6313
rect 22152 6276 22197 6304
rect 22152 6264 22158 6276
rect 22281 6273 22293 6307
rect 22327 6304 22339 6307
rect 22511 6307 22560 6313
rect 22327 6276 22416 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 10965 6239 11023 6245
rect 9784 6208 10548 6236
rect 10612 6208 10732 6236
rect 9674 6168 9680 6180
rect 3283 6140 3832 6168
rect 5092 6140 9680 6168
rect 3283 6137 3295 6140
rect 3237 6131 3295 6137
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 5092 6100 5120 6140
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 10520 6168 10548 6208
rect 10704 6168 10732 6208
rect 10965 6205 10977 6239
rect 11011 6236 11023 6239
rect 12176 6236 12204 6264
rect 22388 6248 22416 6276
rect 22511 6273 22523 6307
rect 22557 6273 22560 6307
rect 22511 6267 22560 6273
rect 22554 6264 22560 6267
rect 22612 6264 22618 6316
rect 25314 6264 25320 6316
rect 25372 6264 25378 6316
rect 25406 6264 25412 6316
rect 25464 6304 25470 6316
rect 25501 6307 25559 6313
rect 25501 6304 25513 6307
rect 25464 6276 25513 6304
rect 25464 6264 25470 6276
rect 25501 6273 25513 6276
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 25590 6264 25596 6316
rect 25648 6264 25654 6316
rect 28276 6313 28304 6344
rect 29730 6332 29736 6344
rect 29788 6332 29794 6384
rect 29914 6332 29920 6384
rect 29972 6372 29978 6384
rect 32674 6372 32680 6384
rect 29972 6344 32680 6372
rect 29972 6332 29978 6344
rect 32674 6332 32680 6344
rect 32732 6332 32738 6384
rect 28261 6307 28319 6313
rect 28261 6273 28273 6307
rect 28307 6273 28319 6307
rect 28261 6267 28319 6273
rect 28528 6307 28586 6313
rect 28528 6273 28540 6307
rect 28574 6304 28586 6307
rect 30466 6304 30472 6316
rect 28574 6276 30472 6304
rect 28574 6273 28586 6276
rect 28528 6267 28586 6273
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 17218 6236 17224 6248
rect 11011 6208 12204 6236
rect 14108 6208 17224 6236
rect 11011 6205 11023 6208
rect 10965 6199 11023 6205
rect 10870 6168 10876 6180
rect 10520 6140 10640 6168
rect 10704 6140 10876 6168
rect 1636 6072 5120 6100
rect 1636 6060 1642 6072
rect 5166 6060 5172 6112
rect 5224 6060 5230 6112
rect 8110 6060 8116 6112
rect 8168 6060 8174 6112
rect 10612 6100 10640 6140
rect 10870 6128 10876 6140
rect 10928 6168 10934 6180
rect 11422 6168 11428 6180
rect 10928 6140 11428 6168
rect 10928 6128 10934 6140
rect 11422 6128 11428 6140
rect 11480 6168 11486 6180
rect 12526 6168 12532 6180
rect 11480 6140 12532 6168
rect 11480 6128 11486 6140
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12618 6100 12624 6112
rect 10612 6072 12624 6100
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14108 6109 14136 6208
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 18782 6196 18788 6248
rect 18840 6236 18846 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18840 6208 19073 6236
rect 18840 6196 18846 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 19150 6196 19156 6248
rect 19208 6196 19214 6248
rect 19242 6196 19248 6248
rect 19300 6196 19306 6248
rect 22370 6196 22376 6248
rect 22428 6196 22434 6248
rect 23106 6196 23112 6248
rect 23164 6236 23170 6248
rect 25424 6236 25452 6264
rect 23164 6208 25452 6236
rect 23164 6196 23170 6208
rect 30650 6196 30656 6248
rect 30708 6236 30714 6248
rect 33134 6236 33140 6248
rect 30708 6208 33140 6236
rect 30708 6196 30714 6208
rect 33134 6196 33140 6208
rect 33192 6236 33198 6248
rect 33594 6236 33600 6248
rect 33192 6208 33600 6236
rect 33192 6196 33198 6208
rect 33594 6196 33600 6208
rect 33652 6196 33658 6248
rect 33888 6236 33916 6412
rect 33980 6412 34520 6440
rect 33980 6313 34008 6412
rect 34514 6400 34520 6412
rect 34572 6440 34578 6452
rect 35618 6440 35624 6452
rect 34572 6412 35624 6440
rect 34572 6400 34578 6412
rect 35618 6400 35624 6412
rect 35676 6400 35682 6452
rect 38197 6443 38255 6449
rect 38197 6409 38209 6443
rect 38243 6440 38255 6443
rect 42613 6443 42671 6449
rect 38243 6412 38792 6440
rect 38243 6409 38255 6412
rect 38197 6403 38255 6409
rect 34146 6332 34152 6384
rect 34204 6372 34210 6384
rect 37921 6375 37979 6381
rect 37921 6372 37933 6375
rect 34204 6344 37933 6372
rect 34204 6332 34210 6344
rect 37921 6341 37933 6344
rect 37967 6341 37979 6375
rect 37921 6335 37979 6341
rect 33965 6307 34023 6313
rect 33965 6273 33977 6307
rect 34011 6273 34023 6307
rect 33965 6267 34023 6273
rect 34057 6307 34115 6313
rect 34057 6273 34069 6307
rect 34103 6304 34115 6307
rect 34330 6304 34336 6316
rect 34103 6276 34336 6304
rect 34103 6273 34115 6276
rect 34057 6267 34115 6273
rect 34330 6264 34336 6276
rect 34388 6264 34394 6316
rect 35526 6264 35532 6316
rect 35584 6304 35590 6316
rect 37642 6304 37648 6316
rect 35584 6276 37648 6304
rect 35584 6264 35590 6276
rect 37642 6264 37648 6276
rect 37700 6264 37706 6316
rect 37826 6264 37832 6316
rect 37884 6264 37890 6316
rect 38010 6264 38016 6316
rect 38068 6264 38074 6316
rect 38764 6304 38792 6412
rect 42613 6409 42625 6443
rect 42659 6440 42671 6443
rect 42794 6440 42800 6452
rect 42659 6412 42800 6440
rect 42659 6409 42671 6412
rect 42613 6403 42671 6409
rect 42794 6400 42800 6412
rect 42852 6400 42858 6452
rect 42886 6400 42892 6452
rect 42944 6440 42950 6452
rect 42944 6412 43208 6440
rect 42944 6400 42950 6412
rect 42150 6332 42156 6384
rect 42208 6372 42214 6384
rect 42208 6344 43024 6372
rect 42208 6332 42214 6344
rect 38913 6307 38971 6313
rect 38913 6304 38925 6307
rect 38764 6276 38925 6304
rect 38913 6273 38925 6276
rect 38959 6273 38971 6307
rect 38913 6267 38971 6273
rect 40126 6264 40132 6316
rect 40184 6304 40190 6316
rect 42996 6313 43024 6344
rect 42889 6307 42947 6313
rect 42889 6304 42901 6307
rect 40184 6276 42901 6304
rect 40184 6264 40190 6276
rect 42889 6273 42901 6276
rect 42935 6273 42947 6307
rect 42889 6267 42947 6273
rect 42981 6307 43039 6313
rect 42981 6273 42993 6307
rect 43027 6273 43039 6307
rect 42981 6267 43039 6273
rect 43070 6264 43076 6316
rect 43128 6264 43134 6316
rect 43180 6304 43208 6412
rect 44082 6400 44088 6452
rect 44140 6400 44146 6452
rect 44266 6400 44272 6452
rect 44324 6400 44330 6452
rect 43901 6375 43959 6381
rect 43901 6341 43913 6375
rect 43947 6372 43959 6375
rect 44100 6372 44128 6400
rect 43947 6344 44128 6372
rect 43947 6341 43959 6344
rect 43901 6335 43959 6341
rect 44085 6307 44143 6313
rect 44085 6304 44097 6307
rect 43180 6276 44097 6304
rect 44085 6273 44097 6276
rect 44131 6304 44143 6307
rect 45278 6304 45284 6316
rect 44131 6276 45284 6304
rect 44131 6273 44143 6276
rect 44085 6267 44143 6273
rect 45278 6264 45284 6276
rect 45336 6264 45342 6316
rect 33888 6208 34376 6236
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 22186 6168 22192 6180
rect 14884 6140 22192 6168
rect 14884 6128 14890 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 22646 6128 22652 6180
rect 22704 6128 22710 6180
rect 29196 6140 31754 6168
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 14056 6072 14105 6100
rect 14056 6060 14062 6072
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 14093 6063 14151 6069
rect 14277 6103 14335 6109
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 14458 6100 14464 6112
rect 14323 6072 14464 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 18874 6060 18880 6112
rect 18932 6060 18938 6112
rect 25130 6060 25136 6112
rect 25188 6060 25194 6112
rect 26602 6060 26608 6112
rect 26660 6100 26666 6112
rect 29196 6100 29224 6140
rect 26660 6072 29224 6100
rect 29641 6103 29699 6109
rect 26660 6060 26666 6072
rect 29641 6069 29653 6103
rect 29687 6100 29699 6103
rect 29914 6100 29920 6112
rect 29687 6072 29920 6100
rect 29687 6069 29699 6072
rect 29641 6063 29699 6069
rect 29914 6060 29920 6072
rect 29972 6100 29978 6112
rect 30282 6100 30288 6112
rect 29972 6072 30288 6100
rect 29972 6060 29978 6072
rect 30282 6060 30288 6072
rect 30340 6060 30346 6112
rect 31726 6100 31754 6140
rect 32674 6128 32680 6180
rect 32732 6168 32738 6180
rect 34241 6171 34299 6177
rect 34241 6168 34253 6171
rect 32732 6140 34253 6168
rect 32732 6128 32738 6140
rect 34241 6137 34253 6140
rect 34287 6137 34299 6171
rect 34241 6131 34299 6137
rect 34146 6100 34152 6112
rect 31726 6072 34152 6100
rect 34146 6060 34152 6072
rect 34204 6060 34210 6112
rect 34348 6100 34376 6208
rect 35986 6196 35992 6248
rect 36044 6236 36050 6248
rect 36354 6236 36360 6248
rect 36044 6208 36360 6236
rect 36044 6196 36050 6208
rect 36354 6196 36360 6208
rect 36412 6236 36418 6248
rect 38657 6239 38715 6245
rect 38657 6236 38669 6239
rect 36412 6208 38669 6236
rect 36412 6196 36418 6208
rect 38657 6205 38669 6208
rect 38703 6205 38715 6239
rect 38657 6199 38715 6205
rect 42797 6239 42855 6245
rect 42797 6205 42809 6239
rect 42843 6205 42855 6239
rect 42797 6199 42855 6205
rect 42812 6168 42840 6199
rect 43070 6168 43076 6180
rect 39960 6140 42748 6168
rect 42812 6140 43076 6168
rect 39960 6100 39988 6140
rect 34348 6072 39988 6100
rect 40034 6060 40040 6112
rect 40092 6100 40098 6112
rect 40310 6100 40316 6112
rect 40092 6072 40316 6100
rect 40092 6060 40098 6072
rect 40310 6060 40316 6072
rect 40368 6060 40374 6112
rect 42720 6100 42748 6140
rect 43070 6128 43076 6140
rect 43128 6128 43134 6180
rect 43622 6100 43628 6112
rect 42720 6072 43628 6100
rect 43622 6060 43628 6072
rect 43680 6060 43686 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 2700 5868 3372 5896
rect 934 5720 940 5772
rect 992 5760 998 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 992 5732 1777 5760
rect 992 5720 998 5732
rect 1765 5729 1777 5732
rect 1811 5729 1823 5763
rect 1765 5723 1823 5729
rect 1578 5652 1584 5704
rect 1636 5652 1642 5704
rect 2700 5701 2728 5868
rect 3344 5828 3372 5868
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 3476 5868 4169 5896
rect 3476 5856 3482 5868
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 6914 5896 6920 5908
rect 4157 5859 4215 5865
rect 4264 5868 6920 5896
rect 4264 5828 4292 5868
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7098 5896 7104 5908
rect 7055 5868 7104 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 9858 5896 9864 5908
rect 7975 5868 9864 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 11514 5856 11520 5908
rect 11572 5896 11578 5908
rect 12342 5896 12348 5908
rect 11572 5868 12348 5896
rect 11572 5856 11578 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 18782 5856 18788 5908
rect 18840 5856 18846 5908
rect 23014 5856 23020 5908
rect 23072 5856 23078 5908
rect 26602 5896 26608 5908
rect 25976 5868 26608 5896
rect 3344 5800 4292 5828
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 11238 5828 11244 5840
rect 9364 5800 11244 5828
rect 9364 5788 9370 5800
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 11974 5828 11980 5840
rect 11388 5800 11980 5828
rect 11388 5788 11394 5800
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 25976 5828 26004 5868
rect 26602 5856 26608 5868
rect 26660 5856 26666 5908
rect 29270 5856 29276 5908
rect 29328 5896 29334 5908
rect 30650 5896 30656 5908
rect 29328 5868 30656 5896
rect 29328 5856 29334 5868
rect 30650 5856 30656 5868
rect 30708 5856 30714 5908
rect 37826 5856 37832 5908
rect 37884 5896 37890 5908
rect 40589 5899 40647 5905
rect 40589 5896 40601 5899
rect 37884 5868 40601 5896
rect 37884 5856 37890 5868
rect 40589 5865 40601 5868
rect 40635 5865 40647 5899
rect 44266 5896 44272 5908
rect 40589 5859 40647 5865
rect 40696 5868 44272 5896
rect 20496 5800 26004 5828
rect 20496 5788 20502 5800
rect 33042 5788 33048 5840
rect 33100 5828 33106 5840
rect 33100 5800 33916 5828
rect 33100 5788 33106 5800
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 4212 5732 5457 5760
rect 4212 5720 4218 5732
rect 5445 5729 5457 5732
rect 5491 5760 5503 5763
rect 6914 5760 6920 5772
rect 5491 5732 6920 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 10413 5763 10471 5769
rect 8720 5732 10364 5760
rect 8720 5720 8726 5732
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7064 5664 8217 5692
rect 7064 5652 7070 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 10336 5692 10364 5732
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10870 5760 10876 5772
rect 10459 5732 10876 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 10980 5732 11565 5760
rect 10980 5692 11008 5732
rect 10336 5664 11008 5692
rect 11054 5652 11060 5704
rect 11112 5652 11118 5704
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 11422 5692 11428 5704
rect 11256 5664 11428 5692
rect 2590 5584 2596 5636
rect 2648 5624 2654 5636
rect 3053 5627 3111 5633
rect 3053 5624 3065 5627
rect 2648 5596 3065 5624
rect 2648 5584 2654 5596
rect 3053 5593 3065 5596
rect 3099 5593 3111 5627
rect 3053 5587 3111 5593
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 3476 5596 4077 5624
rect 3476 5584 3482 5596
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 4798 5584 4804 5636
rect 4856 5584 4862 5636
rect 6822 5584 6828 5636
rect 6880 5624 6886 5636
rect 7561 5627 7619 5633
rect 7561 5624 7573 5627
rect 6880 5596 7573 5624
rect 6880 5584 6886 5596
rect 7561 5593 7573 5596
rect 7607 5593 7619 5627
rect 7561 5587 7619 5593
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 11256 5624 11284 5664
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11537 5701 11565 5732
rect 19426 5720 19432 5772
rect 19484 5720 19490 5772
rect 20806 5720 20812 5772
rect 20864 5760 20870 5772
rect 22002 5760 22008 5772
rect 20864 5732 22008 5760
rect 20864 5720 20870 5732
rect 22002 5720 22008 5732
rect 22060 5760 22066 5772
rect 25498 5760 25504 5772
rect 22060 5732 25504 5760
rect 22060 5720 22066 5732
rect 25498 5720 25504 5732
rect 25556 5720 25562 5772
rect 25866 5720 25872 5772
rect 25924 5760 25930 5772
rect 33888 5769 33916 5800
rect 25961 5763 26019 5769
rect 25961 5760 25973 5763
rect 25924 5732 25973 5760
rect 25924 5720 25930 5732
rect 25961 5729 25973 5732
rect 26007 5729 26019 5763
rect 25961 5723 26019 5729
rect 33873 5763 33931 5769
rect 33873 5729 33885 5763
rect 33919 5729 33931 5763
rect 33873 5723 33931 5729
rect 35802 5720 35808 5772
rect 35860 5760 35866 5772
rect 35860 5732 36492 5760
rect 35860 5720 35866 5732
rect 11522 5695 11580 5701
rect 11522 5661 11534 5695
rect 11568 5661 11580 5695
rect 11522 5655 11580 5661
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 14734 5652 14740 5704
rect 14792 5652 14798 5704
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 18506 5692 18512 5704
rect 18463 5664 18512 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19685 5695 19743 5701
rect 19685 5692 19697 5695
rect 18932 5664 19697 5692
rect 18932 5652 18938 5664
rect 19685 5661 19697 5664
rect 19731 5661 19743 5695
rect 19685 5655 19743 5661
rect 22094 5652 22100 5704
rect 22152 5692 22158 5704
rect 22833 5695 22891 5701
rect 22833 5692 22845 5695
rect 22152 5664 22845 5692
rect 22152 5652 22158 5664
rect 22833 5661 22845 5664
rect 22879 5692 22891 5695
rect 23382 5692 23388 5704
rect 22879 5664 23388 5692
rect 22879 5661 22891 5664
rect 22833 5655 22891 5661
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 25130 5652 25136 5704
rect 25188 5692 25194 5704
rect 26217 5695 26275 5701
rect 26217 5692 26229 5695
rect 25188 5664 26229 5692
rect 25188 5652 25194 5664
rect 26217 5661 26229 5664
rect 26263 5661 26275 5695
rect 26217 5655 26275 5661
rect 30285 5695 30343 5701
rect 30285 5661 30297 5695
rect 30331 5692 30343 5695
rect 31938 5692 31944 5704
rect 30331 5664 31944 5692
rect 30331 5661 30343 5664
rect 30285 5655 30343 5661
rect 31938 5652 31944 5664
rect 31996 5652 32002 5704
rect 33413 5695 33471 5701
rect 33413 5661 33425 5695
rect 33459 5661 33471 5695
rect 33413 5655 33471 5661
rect 9732 5596 11284 5624
rect 9732 5584 9738 5596
rect 11330 5584 11336 5636
rect 11388 5584 11394 5636
rect 12066 5584 12072 5636
rect 12124 5624 12130 5636
rect 12161 5627 12219 5633
rect 12161 5624 12173 5627
rect 12124 5596 12173 5624
rect 12124 5584 12130 5596
rect 12161 5593 12173 5596
rect 12207 5593 12219 5627
rect 12161 5587 12219 5593
rect 12342 5584 12348 5636
rect 12400 5633 12406 5636
rect 12400 5627 12419 5633
rect 12407 5593 12419 5627
rect 12400 5587 12419 5593
rect 12400 5584 12406 5587
rect 14642 5584 14648 5636
rect 14700 5584 14706 5636
rect 18601 5627 18659 5633
rect 18601 5593 18613 5627
rect 18647 5624 18659 5627
rect 18690 5624 18696 5636
rect 18647 5596 18696 5624
rect 18647 5593 18659 5596
rect 18601 5587 18659 5593
rect 18690 5584 18696 5596
rect 18748 5624 18754 5636
rect 22649 5627 22707 5633
rect 18748 5596 19334 5624
rect 18748 5584 18754 5596
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 4893 5559 4951 5565
rect 4893 5556 4905 5559
rect 4764 5528 4905 5556
rect 4764 5516 4770 5528
rect 4893 5525 4905 5528
rect 4939 5525 4951 5559
rect 4893 5519 4951 5525
rect 7926 5516 7932 5568
rect 7984 5565 7990 5568
rect 7984 5556 7996 5565
rect 7984 5528 8029 5556
rect 7984 5519 7996 5528
rect 7984 5516 7990 5519
rect 10594 5516 10600 5568
rect 10652 5556 10658 5568
rect 11701 5559 11759 5565
rect 11701 5556 11713 5559
rect 10652 5528 11713 5556
rect 10652 5516 10658 5528
rect 11701 5525 11713 5528
rect 11747 5525 11759 5559
rect 11701 5519 11759 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 12032 5528 12541 5556
rect 12032 5516 12038 5528
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12529 5519 12587 5525
rect 14274 5516 14280 5568
rect 14332 5516 14338 5568
rect 19306 5556 19334 5596
rect 22649 5593 22661 5627
rect 22695 5624 22707 5627
rect 22738 5624 22744 5636
rect 22695 5596 22744 5624
rect 22695 5593 22707 5596
rect 22649 5587 22707 5593
rect 22738 5584 22744 5596
rect 22796 5584 22802 5636
rect 25314 5584 25320 5636
rect 25372 5624 25378 5636
rect 29730 5624 29736 5636
rect 25372 5596 29736 5624
rect 25372 5584 25378 5596
rect 29730 5584 29736 5596
rect 29788 5584 29794 5636
rect 30530 5627 30588 5633
rect 30530 5624 30542 5627
rect 30300 5596 30542 5624
rect 30300 5568 30328 5596
rect 30530 5593 30542 5596
rect 30576 5593 30588 5627
rect 30530 5587 30588 5593
rect 20809 5559 20867 5565
rect 20809 5556 20821 5559
rect 19306 5528 20821 5556
rect 20809 5525 20821 5528
rect 20855 5525 20867 5559
rect 20809 5519 20867 5525
rect 27338 5516 27344 5568
rect 27396 5516 27402 5568
rect 30282 5516 30288 5568
rect 30340 5516 30346 5568
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 31665 5559 31723 5565
rect 31665 5556 31677 5559
rect 30432 5528 31677 5556
rect 30432 5516 30438 5528
rect 31665 5525 31677 5528
rect 31711 5525 31723 5559
rect 31665 5519 31723 5525
rect 33226 5516 33232 5568
rect 33284 5516 33290 5568
rect 33428 5556 33456 5655
rect 33594 5652 33600 5704
rect 33652 5652 33658 5704
rect 33735 5695 33793 5701
rect 33735 5661 33747 5695
rect 33781 5692 33793 5695
rect 34790 5692 34796 5704
rect 33781 5664 34796 5692
rect 33781 5661 33793 5664
rect 33735 5655 33793 5661
rect 34790 5652 34796 5664
rect 34848 5652 34854 5704
rect 35894 5652 35900 5704
rect 35952 5692 35958 5704
rect 36354 5692 36360 5704
rect 35952 5664 36360 5692
rect 35952 5652 35958 5664
rect 36354 5652 36360 5664
rect 36412 5652 36418 5704
rect 36464 5692 36492 5732
rect 36613 5695 36671 5701
rect 36613 5692 36625 5695
rect 36464 5664 36625 5692
rect 36613 5661 36625 5664
rect 36659 5661 36671 5695
rect 36613 5655 36671 5661
rect 40034 5652 40040 5704
rect 40092 5652 40098 5704
rect 40218 5652 40224 5704
rect 40276 5652 40282 5704
rect 40402 5652 40408 5704
rect 40460 5652 40466 5704
rect 33505 5627 33563 5633
rect 33505 5593 33517 5627
rect 33551 5624 33563 5627
rect 34330 5624 34336 5636
rect 33551 5596 34336 5624
rect 33551 5593 33563 5596
rect 33505 5587 33563 5593
rect 34330 5584 34336 5596
rect 34388 5584 34394 5636
rect 40310 5584 40316 5636
rect 40368 5584 40374 5636
rect 35986 5556 35992 5568
rect 33428 5528 35992 5556
rect 35986 5516 35992 5528
rect 36044 5516 36050 5568
rect 36446 5516 36452 5568
rect 36504 5556 36510 5568
rect 37737 5559 37795 5565
rect 37737 5556 37749 5559
rect 36504 5528 37749 5556
rect 36504 5516 36510 5528
rect 37737 5525 37749 5528
rect 37783 5556 37795 5559
rect 40696 5556 40724 5868
rect 44266 5856 44272 5868
rect 44324 5856 44330 5908
rect 41046 5720 41052 5772
rect 41104 5760 41110 5772
rect 41141 5763 41199 5769
rect 41141 5760 41153 5763
rect 41104 5732 41153 5760
rect 41104 5720 41110 5732
rect 41141 5729 41153 5732
rect 41187 5729 41199 5763
rect 41141 5723 41199 5729
rect 43622 5720 43628 5772
rect 43680 5720 43686 5772
rect 42886 5652 42892 5704
rect 42944 5692 42950 5704
rect 43165 5695 43223 5701
rect 43165 5692 43177 5695
rect 42944 5664 43177 5692
rect 42944 5652 42950 5664
rect 43165 5661 43177 5664
rect 43211 5661 43223 5695
rect 43165 5655 43223 5661
rect 43438 5652 43444 5704
rect 43496 5701 43502 5704
rect 43496 5695 43525 5701
rect 43513 5661 43525 5695
rect 43496 5655 43525 5661
rect 43496 5652 43502 5655
rect 41408 5627 41466 5633
rect 41408 5593 41420 5627
rect 41454 5624 41466 5627
rect 42981 5627 43039 5633
rect 42981 5624 42993 5627
rect 41454 5596 42993 5624
rect 41454 5593 41466 5596
rect 41408 5587 41466 5593
rect 42981 5593 42993 5596
rect 43027 5593 43039 5627
rect 42981 5587 43039 5593
rect 43257 5627 43315 5633
rect 43257 5593 43269 5627
rect 43303 5593 43315 5627
rect 43257 5587 43315 5593
rect 43349 5627 43407 5633
rect 43349 5593 43361 5627
rect 43395 5624 43407 5627
rect 43622 5624 43628 5636
rect 43395 5596 43628 5624
rect 43395 5593 43407 5596
rect 43349 5587 43407 5593
rect 37783 5528 40724 5556
rect 37783 5525 37795 5528
rect 37737 5519 37795 5525
rect 41138 5516 41144 5568
rect 41196 5556 41202 5568
rect 42334 5556 42340 5568
rect 41196 5528 42340 5556
rect 41196 5516 41202 5528
rect 42334 5516 42340 5528
rect 42392 5516 42398 5568
rect 42521 5559 42579 5565
rect 42521 5525 42533 5559
rect 42567 5556 42579 5559
rect 42794 5556 42800 5568
rect 42567 5528 42800 5556
rect 42567 5525 42579 5528
rect 42521 5519 42579 5525
rect 42794 5516 42800 5528
rect 42852 5516 42858 5568
rect 43272 5556 43300 5587
rect 43622 5584 43628 5596
rect 43680 5584 43686 5636
rect 43990 5556 43996 5568
rect 43272 5528 43996 5556
rect 43990 5516 43996 5528
rect 44048 5516 44054 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 7558 5352 7564 5364
rect 6564 5324 7564 5352
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 3418 5284 3424 5296
rect 992 5256 3424 5284
rect 992 5244 998 5256
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 5534 5284 5540 5296
rect 4172 5256 5540 5284
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5185 2559 5219
rect 2501 5179 2559 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 992 5120 1777 5148
rect 992 5108 998 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 1026 5040 1032 5092
rect 1084 5080 1090 5092
rect 2516 5080 2544 5179
rect 3878 5176 3884 5228
rect 3936 5176 3942 5228
rect 4172 5225 4200 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 5905 5287 5963 5293
rect 5905 5253 5917 5287
rect 5951 5284 5963 5287
rect 6564 5284 6592 5324
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 8662 5312 8668 5364
rect 8720 5352 8726 5364
rect 8720 5324 10640 5352
rect 8720 5312 8726 5324
rect 8021 5287 8079 5293
rect 5951 5256 6592 5284
rect 6656 5256 7420 5284
rect 5951 5253 5963 5256
rect 5905 5247 5963 5253
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 4356 5148 4384 5179
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 5132 5188 5365 5216
rect 5132 5176 5138 5188
rect 5353 5185 5365 5188
rect 5399 5216 5411 5219
rect 6656 5216 6684 5256
rect 5399 5188 6684 5216
rect 6733 5219 6791 5225
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7282 5216 7288 5228
rect 6779 5188 7288 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 7392 5216 7420 5256
rect 8021 5253 8033 5287
rect 8067 5284 8079 5287
rect 8110 5284 8116 5296
rect 8067 5256 8116 5284
rect 8067 5253 8079 5256
rect 8021 5247 8079 5253
rect 8110 5244 8116 5256
rect 8168 5244 8174 5296
rect 8205 5287 8263 5293
rect 8205 5253 8217 5287
rect 8251 5284 8263 5287
rect 8294 5284 8300 5296
rect 8251 5256 8300 5284
rect 8251 5253 8263 5256
rect 8205 5247 8263 5253
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 10502 5284 10508 5296
rect 8404 5256 10508 5284
rect 8404 5216 8432 5256
rect 10502 5244 10508 5256
rect 10560 5244 10566 5296
rect 10612 5284 10640 5324
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 11882 5352 11888 5364
rect 10928 5324 11888 5352
rect 10928 5312 10934 5324
rect 11882 5312 11888 5324
rect 11940 5352 11946 5364
rect 12342 5352 12348 5364
rect 11940 5324 12348 5352
rect 11940 5312 11946 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14148 5324 14596 5352
rect 14148 5312 14154 5324
rect 10612 5256 10916 5284
rect 7392 5188 8432 5216
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 10888 5225 10916 5256
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 10652 5188 10701 5216
rect 10652 5176 10658 5188
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5216 13323 5219
rect 13354 5216 13360 5228
rect 13311 5188 13360 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 3108 5120 4384 5148
rect 3108 5108 3114 5120
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 6270 5148 6276 5160
rect 4672 5120 6276 5148
rect 4672 5108 4678 5120
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 6822 5108 6828 5160
rect 6880 5148 6886 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6880 5120 6929 5148
rect 6880 5108 6886 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5148 7067 5151
rect 7190 5148 7196 5160
rect 7055 5120 7196 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 7190 5108 7196 5120
rect 7248 5148 7254 5160
rect 7650 5148 7656 5160
rect 7248 5120 7656 5148
rect 7248 5108 7254 5120
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 10980 5148 11008 5179
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13532 5219 13590 5225
rect 13532 5185 13544 5219
rect 13578 5216 13590 5219
rect 14274 5216 14280 5228
rect 13578 5188 14280 5216
rect 13578 5185 13590 5188
rect 13532 5179 13590 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14568 5216 14596 5324
rect 14642 5312 14648 5364
rect 14700 5312 14706 5364
rect 18785 5355 18843 5361
rect 18785 5321 18797 5355
rect 18831 5352 18843 5355
rect 19150 5352 19156 5364
rect 18831 5324 19156 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 23934 5312 23940 5364
rect 23992 5352 23998 5364
rect 27338 5352 27344 5364
rect 23992 5324 27344 5352
rect 23992 5312 23998 5324
rect 27338 5312 27344 5324
rect 27396 5312 27402 5364
rect 27522 5352 27528 5364
rect 27448 5324 27528 5352
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16853 5287 16911 5293
rect 16853 5284 16865 5287
rect 16540 5256 16865 5284
rect 16540 5244 16546 5256
rect 16853 5253 16865 5256
rect 16899 5253 16911 5287
rect 16853 5247 16911 5253
rect 17069 5287 17127 5293
rect 17069 5253 17081 5287
rect 17115 5284 17127 5287
rect 17115 5256 18552 5284
rect 17115 5253 17127 5256
rect 17069 5247 17127 5253
rect 18524 5228 18552 5256
rect 18966 5244 18972 5296
rect 19024 5284 19030 5296
rect 23290 5284 23296 5296
rect 19024 5256 23296 5284
rect 19024 5244 19030 5256
rect 23290 5244 23296 5256
rect 23348 5244 23354 5296
rect 23382 5244 23388 5296
rect 23440 5284 23446 5296
rect 23753 5287 23811 5293
rect 23753 5284 23765 5287
rect 23440 5256 23765 5284
rect 23440 5244 23446 5256
rect 23753 5253 23765 5256
rect 23799 5253 23811 5287
rect 23753 5247 23811 5253
rect 23842 5244 23848 5296
rect 23900 5284 23906 5296
rect 27448 5293 27476 5324
rect 27522 5312 27528 5324
rect 27580 5312 27586 5364
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 27801 5355 27859 5361
rect 27801 5352 27813 5355
rect 27672 5324 27813 5352
rect 27672 5312 27678 5324
rect 27801 5321 27813 5324
rect 27847 5321 27859 5355
rect 27801 5315 27859 5321
rect 27890 5312 27896 5364
rect 27948 5352 27954 5364
rect 27948 5324 30144 5352
rect 27948 5312 27954 5324
rect 24121 5287 24179 5293
rect 24121 5284 24133 5287
rect 23900 5256 24133 5284
rect 23900 5244 23906 5256
rect 24121 5253 24133 5256
rect 24167 5253 24179 5287
rect 24121 5247 24179 5253
rect 27433 5287 27491 5293
rect 27433 5253 27445 5287
rect 27479 5253 27491 5287
rect 30006 5284 30012 5296
rect 27433 5247 27491 5253
rect 29932 5256 30012 5284
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 14568 5188 15761 5216
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 18564 5188 18613 5216
rect 18564 5176 18570 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 10836 5120 11008 5148
rect 15841 5151 15899 5157
rect 10836 5108 10842 5120
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 18690 5148 18696 5160
rect 15887 5120 17264 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 1084 5052 2544 5080
rect 2685 5083 2743 5089
rect 1084 5040 1090 5052
rect 2685 5049 2697 5083
rect 2731 5080 2743 5083
rect 2731 5052 10732 5080
rect 2731 5049 2743 5052
rect 2685 5043 2743 5049
rect 3694 4972 3700 5024
rect 3752 4972 3758 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 8294 5012 8300 5024
rect 3936 4984 8300 5012
rect 3936 4972 3942 4984
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8386 4972 8392 5024
rect 8444 4972 8450 5024
rect 10502 4972 10508 5024
rect 10560 4972 10566 5024
rect 10704 5012 10732 5052
rect 15930 5040 15936 5092
rect 15988 5040 15994 5092
rect 17236 5089 17264 5120
rect 18248 5120 18696 5148
rect 17221 5083 17279 5089
rect 17221 5049 17233 5083
rect 17267 5080 17279 5083
rect 17862 5080 17868 5092
rect 17267 5052 17868 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 18248 5024 18276 5120
rect 18690 5108 18696 5120
rect 18748 5148 18754 5160
rect 18800 5148 18828 5179
rect 22646 5176 22652 5228
rect 22704 5176 22710 5228
rect 22830 5176 22836 5228
rect 22888 5176 22894 5228
rect 24026 5176 24032 5228
rect 24084 5176 24090 5228
rect 24486 5176 24492 5228
rect 24544 5176 24550 5228
rect 25498 5176 25504 5228
rect 25556 5216 25562 5228
rect 27338 5225 27344 5228
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 25556 5188 27169 5216
rect 25556 5176 25562 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27305 5219 27344 5225
rect 27305 5185 27317 5219
rect 27305 5179 27344 5185
rect 27338 5176 27344 5179
rect 27396 5176 27402 5228
rect 27522 5174 27528 5226
rect 27580 5174 27586 5226
rect 27622 5219 27680 5225
rect 27622 5185 27634 5219
rect 27668 5185 27680 5219
rect 27622 5179 27680 5185
rect 18748 5120 18828 5148
rect 18748 5108 18754 5120
rect 22649 5083 22707 5089
rect 22649 5049 22661 5083
rect 22695 5080 22707 5083
rect 25590 5080 25596 5092
rect 22695 5052 25596 5080
rect 22695 5049 22707 5052
rect 22649 5043 22707 5049
rect 25590 5040 25596 5052
rect 25648 5040 25654 5092
rect 13998 5012 14004 5024
rect 10704 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14734 4972 14740 5024
rect 14792 5012 14798 5024
rect 15565 5015 15623 5021
rect 15565 5012 15577 5015
rect 14792 4984 15577 5012
rect 14792 4972 14798 4984
rect 15565 4981 15577 4984
rect 15611 4981 15623 5015
rect 15565 4975 15623 4981
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16264 4984 17049 5012
rect 16264 4972 16270 4984
rect 17037 4981 17049 4984
rect 17083 5012 17095 5015
rect 18230 5012 18236 5024
rect 17083 4984 18236 5012
rect 17083 4981 17095 4984
rect 17037 4975 17095 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 22554 5012 22560 5024
rect 22244 4984 22560 5012
rect 22244 4972 22250 4984
rect 22554 4972 22560 4984
rect 22612 5012 22618 5024
rect 27632 5012 27660 5179
rect 29270 5176 29276 5228
rect 29328 5216 29334 5228
rect 29932 5225 29960 5256
rect 30006 5244 30012 5256
rect 30064 5244 30070 5296
rect 30116 5284 30144 5324
rect 30282 5312 30288 5364
rect 30340 5352 30346 5364
rect 30469 5355 30527 5361
rect 30469 5352 30481 5355
rect 30340 5324 30481 5352
rect 30340 5312 30346 5324
rect 30469 5321 30481 5324
rect 30515 5321 30527 5355
rect 30469 5315 30527 5321
rect 33594 5312 33600 5364
rect 33652 5352 33658 5364
rect 33962 5352 33968 5364
rect 33652 5324 33968 5352
rect 33652 5312 33658 5324
rect 33962 5312 33968 5324
rect 34020 5312 34026 5364
rect 35345 5355 35403 5361
rect 35345 5321 35357 5355
rect 35391 5352 35403 5355
rect 36265 5355 36323 5361
rect 36265 5352 36277 5355
rect 35391 5324 36277 5352
rect 35391 5321 35403 5324
rect 35345 5315 35403 5321
rect 36265 5321 36277 5324
rect 36311 5352 36323 5355
rect 37826 5352 37832 5364
rect 36311 5324 37832 5352
rect 36311 5321 36323 5324
rect 36265 5315 36323 5321
rect 37826 5312 37832 5324
rect 37884 5352 37890 5364
rect 38194 5352 38200 5364
rect 37884 5324 38200 5352
rect 37884 5312 37890 5324
rect 38194 5312 38200 5324
rect 38252 5312 38258 5364
rect 38378 5312 38384 5364
rect 38436 5352 38442 5364
rect 41690 5352 41696 5364
rect 38436 5324 41696 5352
rect 38436 5312 38442 5324
rect 30116 5256 31754 5284
rect 29733 5219 29791 5225
rect 29733 5216 29745 5219
rect 29328 5188 29745 5216
rect 29328 5176 29334 5188
rect 29733 5185 29745 5188
rect 29779 5185 29791 5219
rect 29733 5179 29791 5185
rect 29917 5219 29975 5225
rect 29917 5185 29929 5219
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 30098 5176 30104 5228
rect 30156 5176 30162 5228
rect 30285 5219 30343 5225
rect 30285 5185 30297 5219
rect 30331 5216 30343 5219
rect 30374 5216 30380 5228
rect 30331 5188 30380 5216
rect 30331 5185 30343 5188
rect 30285 5179 30343 5185
rect 30374 5176 30380 5188
rect 30432 5176 30438 5228
rect 31726 5216 31754 5256
rect 33226 5244 33232 5296
rect 33284 5284 33290 5296
rect 34210 5287 34268 5293
rect 34210 5284 34222 5287
rect 33284 5256 34222 5284
rect 33284 5244 33290 5256
rect 34210 5253 34222 5256
rect 34256 5253 34268 5287
rect 41138 5284 41144 5296
rect 34210 5247 34268 5253
rect 35544 5256 41144 5284
rect 35544 5216 35572 5256
rect 41138 5244 41144 5256
rect 41196 5244 41202 5296
rect 41524 5293 41552 5324
rect 41690 5312 41696 5324
rect 41748 5312 41754 5364
rect 42794 5312 42800 5364
rect 42852 5352 42858 5364
rect 44085 5355 44143 5361
rect 44085 5352 44097 5355
rect 42852 5324 44097 5352
rect 42852 5312 42858 5324
rect 44085 5321 44097 5324
rect 44131 5352 44143 5355
rect 45189 5355 45247 5361
rect 45189 5352 45201 5355
rect 44131 5324 45201 5352
rect 44131 5321 44143 5324
rect 44085 5315 44143 5321
rect 45189 5321 45201 5324
rect 45235 5352 45247 5355
rect 49694 5352 49700 5364
rect 45235 5324 49700 5352
rect 45235 5321 45247 5324
rect 45189 5315 45247 5321
rect 49694 5312 49700 5324
rect 49752 5312 49758 5364
rect 41509 5287 41567 5293
rect 41509 5253 41521 5287
rect 41555 5253 41567 5287
rect 41509 5247 41567 5253
rect 42334 5244 42340 5296
rect 42392 5284 42398 5296
rect 56962 5284 56968 5296
rect 42392 5256 56968 5284
rect 42392 5244 42398 5256
rect 56962 5244 56968 5256
rect 57020 5244 57026 5296
rect 31726 5188 35572 5216
rect 41325 5219 41383 5225
rect 41325 5185 41337 5219
rect 41371 5185 41383 5219
rect 41325 5179 41383 5185
rect 30006 5108 30012 5160
rect 30064 5108 30070 5160
rect 33870 5108 33876 5160
rect 33928 5148 33934 5160
rect 33965 5151 34023 5157
rect 33965 5148 33977 5151
rect 33928 5120 33977 5148
rect 33928 5108 33934 5120
rect 33965 5117 33977 5120
rect 34011 5117 34023 5151
rect 33965 5111 34023 5117
rect 36354 5108 36360 5160
rect 36412 5108 36418 5160
rect 36538 5108 36544 5160
rect 36596 5108 36602 5160
rect 35897 5083 35955 5089
rect 35897 5049 35909 5083
rect 35943 5080 35955 5083
rect 35986 5080 35992 5092
rect 35943 5052 35992 5080
rect 35943 5049 35955 5052
rect 35897 5043 35955 5049
rect 35986 5040 35992 5052
rect 36044 5040 36050 5092
rect 40034 5040 40040 5092
rect 40092 5080 40098 5092
rect 41340 5080 41368 5179
rect 41414 5176 41420 5228
rect 41472 5176 41478 5228
rect 41627 5219 41685 5225
rect 41627 5185 41639 5219
rect 41673 5185 41685 5219
rect 41627 5179 41685 5185
rect 41642 5148 41670 5179
rect 41782 5176 41788 5228
rect 41840 5176 41846 5228
rect 43993 5219 44051 5225
rect 43993 5185 44005 5219
rect 44039 5185 44051 5219
rect 43993 5179 44051 5185
rect 45204 5188 45416 5216
rect 43438 5148 43444 5160
rect 41642 5120 43444 5148
rect 43438 5108 43444 5120
rect 43496 5108 43502 5160
rect 43625 5083 43683 5089
rect 43625 5080 43637 5083
rect 40092 5052 41276 5080
rect 41340 5052 43637 5080
rect 40092 5040 40098 5052
rect 22612 4984 27660 5012
rect 22612 4972 22618 4984
rect 29730 4972 29736 5024
rect 29788 5012 29794 5024
rect 38286 5012 38292 5024
rect 29788 4984 38292 5012
rect 29788 4972 29794 4984
rect 38286 4972 38292 4984
rect 38344 4972 38350 5024
rect 38746 4972 38752 5024
rect 38804 5012 38810 5024
rect 41141 5015 41199 5021
rect 41141 5012 41153 5015
rect 38804 4984 41153 5012
rect 38804 4972 38810 4984
rect 41141 4981 41153 4984
rect 41187 4981 41199 5015
rect 41248 5012 41276 5052
rect 43625 5049 43637 5052
rect 43671 5049 43683 5083
rect 43625 5043 43683 5049
rect 44008 5080 44036 5179
rect 44174 5108 44180 5160
rect 44232 5148 44238 5160
rect 44634 5148 44640 5160
rect 44232 5120 44640 5148
rect 44232 5108 44238 5120
rect 44634 5108 44640 5120
rect 44692 5148 44698 5160
rect 45204 5148 45232 5188
rect 44692 5120 45232 5148
rect 44692 5108 44698 5120
rect 45278 5108 45284 5160
rect 45336 5108 45342 5160
rect 45388 5157 45416 5188
rect 45373 5151 45431 5157
rect 45373 5117 45385 5151
rect 45419 5117 45431 5151
rect 45373 5111 45431 5117
rect 44008 5052 51074 5080
rect 44008 5012 44036 5052
rect 41248 4984 44036 5012
rect 41141 4975 41199 4981
rect 44818 4972 44824 5024
rect 44876 4972 44882 5024
rect 51046 5012 51074 5052
rect 51626 5012 51632 5024
rect 51046 4984 51632 5012
rect 51626 4972 51632 4984
rect 51684 4972 51690 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 1636 4780 2774 4808
rect 1636 4768 1642 4780
rect 2746 4740 2774 4780
rect 3050 4768 3056 4820
rect 3108 4768 3114 4820
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 5718 4808 5724 4820
rect 5123 4780 5724 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 8570 4808 8576 4820
rect 6656 4780 8576 4808
rect 6656 4740 6684 4780
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 11480 4780 11621 4808
rect 11480 4768 11486 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 16025 4811 16083 4817
rect 16025 4808 16037 4811
rect 15988 4780 16037 4808
rect 15988 4768 15994 4780
rect 16025 4777 16037 4780
rect 16071 4777 16083 4811
rect 16025 4771 16083 4777
rect 22097 4811 22155 4817
rect 22097 4777 22109 4811
rect 22143 4777 22155 4811
rect 22097 4771 22155 4777
rect 2746 4712 6684 4740
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 20070 4740 20076 4752
rect 19852 4712 20076 4740
rect 19852 4700 19858 4712
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 19705 4675 19763 4681
rect 5224 4644 5764 4672
rect 5224 4632 5230 4644
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 1762 4604 1768 4616
rect 1719 4576 1768 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 1762 4564 1768 4576
rect 1820 4604 1826 4616
rect 2498 4604 2504 4616
rect 1820 4576 2504 4604
rect 1820 4564 1826 4576
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 5350 4604 5356 4616
rect 4304 4576 5356 4604
rect 4304 4564 4310 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 1940 4539 1998 4545
rect 1940 4505 1952 4539
rect 1986 4536 1998 4539
rect 3694 4536 3700 4548
rect 1986 4508 3700 4536
rect 1986 4505 1998 4508
rect 1940 4499 1998 4505
rect 3694 4496 3700 4508
rect 3752 4496 3758 4548
rect 4062 4496 4068 4548
rect 4120 4496 4126 4548
rect 5460 4536 5488 4567
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 5736 4613 5764 4644
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 20533 4675 20591 4681
rect 20533 4672 20545 4675
rect 19751 4644 20545 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 20533 4641 20545 4644
rect 20579 4641 20591 4675
rect 22112 4672 22140 4771
rect 22646 4768 22652 4820
rect 22704 4808 22710 4820
rect 22741 4811 22799 4817
rect 22741 4808 22753 4811
rect 22704 4780 22753 4808
rect 22704 4768 22710 4780
rect 22741 4777 22753 4780
rect 22787 4777 22799 4811
rect 22741 4771 22799 4777
rect 25130 4768 25136 4820
rect 25188 4808 25194 4820
rect 27525 4811 27583 4817
rect 27525 4808 27537 4811
rect 25188 4780 27537 4808
rect 25188 4768 25194 4780
rect 27525 4777 27537 4780
rect 27571 4808 27583 4811
rect 29822 4808 29828 4820
rect 27571 4780 29828 4808
rect 27571 4777 27583 4780
rect 27525 4771 27583 4777
rect 29822 4768 29828 4780
rect 29880 4768 29886 4820
rect 30006 4768 30012 4820
rect 30064 4808 30070 4820
rect 30285 4811 30343 4817
rect 30285 4808 30297 4811
rect 30064 4780 30297 4808
rect 30064 4768 30070 4780
rect 30285 4777 30297 4780
rect 30331 4777 30343 4811
rect 30285 4771 30343 4777
rect 36538 4768 36544 4820
rect 36596 4808 36602 4820
rect 36596 4780 39344 4808
rect 36596 4768 36602 4780
rect 22281 4743 22339 4749
rect 22281 4709 22293 4743
rect 22327 4740 22339 4743
rect 22830 4740 22836 4752
rect 22327 4712 22836 4740
rect 22327 4709 22339 4712
rect 22281 4703 22339 4709
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 23658 4700 23664 4752
rect 23716 4740 23722 4752
rect 23716 4712 25820 4740
rect 23716 4700 23722 4712
rect 23750 4672 23756 4684
rect 22112 4644 23756 4672
rect 20533 4635 20591 4641
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 10502 4613 10508 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6972 4576 7205 4604
rect 6972 4564 6978 4576
rect 7193 4573 7205 4576
rect 7239 4604 7251 4607
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 7239 4576 10241 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10496 4604 10508 4613
rect 10463 4576 10508 4604
rect 10229 4567 10287 4573
rect 10496 4567 10508 4576
rect 10502 4564 10508 4567
rect 10560 4564 10566 4616
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 16206 4604 16212 4616
rect 10836 4576 16212 4604
rect 10836 4564 10842 4576
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16347 4576 18368 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 5626 4536 5632 4548
rect 5460 4508 5632 4536
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 6270 4496 6276 4548
rect 6328 4496 6334 4548
rect 7460 4539 7518 4545
rect 7460 4505 7472 4539
rect 7506 4536 7518 4539
rect 8386 4536 8392 4548
rect 7506 4508 8392 4536
rect 7506 4505 7518 4508
rect 7460 4499 7518 4505
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 16025 4539 16083 4545
rect 16025 4536 16037 4539
rect 15344 4508 16037 4536
rect 15344 4496 15350 4508
rect 16025 4505 16037 4508
rect 16071 4536 16083 4539
rect 16482 4536 16488 4548
rect 16071 4508 16488 4536
rect 16071 4505 16083 4508
rect 16025 4499 16083 4505
rect 16482 4496 16488 4508
rect 16540 4536 16546 4548
rect 17402 4536 17408 4548
rect 16540 4508 17408 4536
rect 16540 4496 16546 4508
rect 17402 4496 17408 4508
rect 17460 4536 17466 4548
rect 17460 4508 17908 4536
rect 17460 4496 17466 4508
rect 4154 4428 4160 4480
rect 4212 4428 4218 4480
rect 6362 4428 6368 4480
rect 6420 4428 6426 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 14826 4468 14832 4480
rect 7616 4440 14832 4468
rect 7616 4428 7622 4440
rect 14826 4428 14832 4440
rect 14884 4468 14890 4480
rect 16114 4468 16120 4480
rect 14884 4440 16120 4468
rect 14884 4428 14890 4440
rect 16114 4428 16120 4440
rect 16172 4428 16178 4480
rect 17880 4468 17908 4508
rect 17954 4496 17960 4548
rect 18012 4496 18018 4548
rect 18230 4496 18236 4548
rect 18288 4496 18294 4548
rect 18340 4545 18368 4576
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 19392 4576 19625 4604
rect 19392 4564 19398 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 19794 4564 19800 4616
rect 19852 4564 19858 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 19978 4604 19984 4616
rect 19935 4576 19984 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20441 4607 20499 4613
rect 20441 4573 20453 4607
rect 20487 4604 20499 4607
rect 23017 4607 23075 4613
rect 23017 4604 23029 4607
rect 20487 4576 23029 4604
rect 20487 4573 20499 4576
rect 20441 4567 20499 4573
rect 18325 4539 18383 4545
rect 18325 4505 18337 4539
rect 18371 4536 18383 4539
rect 18506 4536 18512 4548
rect 18371 4508 18512 4536
rect 18371 4505 18383 4508
rect 18325 4499 18383 4505
rect 18506 4496 18512 4508
rect 18564 4496 18570 4548
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 20456 4536 20484 4567
rect 22112 4545 22140 4576
rect 23017 4573 23029 4576
rect 23063 4604 23075 4607
rect 23842 4604 23848 4616
rect 23063 4576 23848 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 18739 4508 20484 4536
rect 21913 4539 21971 4545
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 21913 4505 21925 4539
rect 21959 4536 21971 4539
rect 22112 4539 22171 4545
rect 21959 4508 21993 4536
rect 22112 4508 22125 4539
rect 21959 4505 21971 4508
rect 21913 4499 21971 4505
rect 22113 4505 22125 4508
rect 22159 4505 22171 4539
rect 22113 4499 22171 4505
rect 22741 4539 22799 4545
rect 22741 4505 22753 4539
rect 22787 4536 22799 4539
rect 23934 4536 23940 4548
rect 22787 4508 23940 4536
rect 22787 4505 22799 4508
rect 22741 4499 22799 4505
rect 18141 4471 18199 4477
rect 18141 4468 18153 4471
rect 17880 4440 18153 4468
rect 18141 4437 18153 4440
rect 18187 4437 18199 4471
rect 18141 4431 18199 4437
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4468 19487 4471
rect 19978 4468 19984 4480
rect 19475 4440 19984 4468
rect 19475 4437 19487 4440
rect 19429 4431 19487 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 21818 4428 21824 4480
rect 21876 4468 21882 4480
rect 21928 4468 21956 4499
rect 22756 4468 22784 4499
rect 23934 4496 23940 4508
rect 23992 4496 23998 4548
rect 21876 4440 22784 4468
rect 22925 4471 22983 4477
rect 21876 4428 21882 4440
rect 22925 4437 22937 4471
rect 22971 4468 22983 4471
rect 23750 4468 23756 4480
rect 22971 4440 23756 4468
rect 22971 4437 22983 4440
rect 22925 4431 22983 4437
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 25792 4468 25820 4712
rect 37642 4700 37648 4752
rect 37700 4740 37706 4752
rect 38010 4740 38016 4752
rect 37700 4712 38016 4740
rect 37700 4700 37706 4712
rect 38010 4700 38016 4712
rect 38068 4740 38074 4752
rect 38378 4740 38384 4752
rect 38068 4712 38384 4740
rect 38068 4700 38074 4712
rect 38378 4700 38384 4712
rect 38436 4700 38442 4752
rect 38749 4743 38807 4749
rect 38749 4709 38761 4743
rect 38795 4709 38807 4743
rect 38749 4703 38807 4709
rect 25866 4632 25872 4684
rect 25924 4672 25930 4684
rect 26145 4675 26203 4681
rect 26145 4672 26157 4675
rect 25924 4644 26157 4672
rect 25924 4632 25930 4644
rect 26145 4641 26157 4644
rect 26191 4641 26203 4675
rect 26145 4635 26203 4641
rect 29914 4632 29920 4684
rect 29972 4632 29978 4684
rect 38764 4672 38792 4703
rect 39316 4681 39344 4780
rect 41414 4768 41420 4820
rect 41472 4808 41478 4820
rect 41690 4808 41696 4820
rect 41472 4780 41696 4808
rect 41472 4768 41478 4780
rect 41690 4768 41696 4780
rect 41748 4808 41754 4820
rect 42886 4808 42892 4820
rect 41748 4780 42892 4808
rect 41748 4768 41754 4780
rect 42886 4768 42892 4780
rect 42944 4808 42950 4820
rect 43990 4808 43996 4820
rect 42944 4780 43996 4808
rect 42944 4768 42950 4780
rect 43990 4768 43996 4780
rect 44048 4768 44054 4820
rect 43070 4740 43076 4752
rect 41340 4712 43076 4740
rect 37844 4644 38792 4672
rect 39301 4675 39359 4681
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4604 30159 4607
rect 31202 4604 31208 4616
rect 30147 4576 31208 4604
rect 30147 4573 30159 4576
rect 30101 4567 30159 4573
rect 31202 4564 31208 4576
rect 31260 4564 31266 4616
rect 37844 4613 37872 4644
rect 39301 4641 39313 4675
rect 39347 4641 39359 4675
rect 39301 4635 39359 4641
rect 37829 4607 37887 4613
rect 37829 4573 37841 4607
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 38010 4564 38016 4616
rect 38068 4564 38074 4616
rect 38102 4564 38108 4616
rect 38160 4613 38166 4616
rect 38160 4607 38189 4613
rect 38177 4573 38189 4607
rect 38160 4567 38189 4573
rect 38160 4564 38166 4567
rect 38286 4564 38292 4616
rect 38344 4564 38350 4616
rect 26412 4539 26470 4545
rect 26412 4505 26424 4539
rect 26458 4536 26470 4539
rect 30006 4536 30012 4548
rect 26458 4508 30012 4536
rect 26458 4505 26470 4508
rect 26412 4499 26470 4505
rect 30006 4496 30012 4508
rect 30064 4496 30070 4548
rect 36262 4496 36268 4548
rect 36320 4536 36326 4548
rect 37921 4539 37979 4545
rect 37921 4536 37933 4539
rect 36320 4508 37933 4536
rect 36320 4496 36326 4508
rect 37921 4505 37933 4508
rect 37967 4505 37979 4539
rect 38120 4536 38148 4564
rect 41340 4536 41368 4712
rect 43070 4700 43076 4712
rect 43128 4700 43134 4752
rect 43990 4672 43996 4684
rect 41616 4644 43996 4672
rect 41616 4613 41644 4644
rect 43990 4632 43996 4644
rect 44048 4632 44054 4684
rect 41601 4607 41659 4613
rect 41601 4573 41613 4607
rect 41647 4573 41659 4607
rect 41601 4567 41659 4573
rect 41690 4564 41696 4616
rect 41748 4564 41754 4616
rect 41782 4564 41788 4616
rect 41840 4564 41846 4616
rect 42058 4564 42064 4616
rect 42116 4564 42122 4616
rect 41903 4539 41961 4545
rect 41903 4536 41915 4539
rect 38120 4508 41644 4536
rect 37921 4499 37979 4505
rect 30834 4468 30840 4480
rect 25792 4440 30840 4468
rect 30834 4428 30840 4440
rect 30892 4428 30898 4480
rect 37645 4471 37703 4477
rect 37645 4437 37657 4471
rect 37691 4468 37703 4471
rect 38286 4468 38292 4480
rect 37691 4440 38292 4468
rect 37691 4437 37703 4440
rect 37645 4431 37703 4437
rect 38286 4428 38292 4440
rect 38344 4428 38350 4480
rect 39114 4428 39120 4480
rect 39172 4428 39178 4480
rect 39209 4471 39267 4477
rect 39209 4437 39221 4471
rect 39255 4468 39267 4471
rect 40218 4468 40224 4480
rect 39255 4440 40224 4468
rect 39255 4437 39267 4440
rect 39209 4431 39267 4437
rect 40218 4428 40224 4440
rect 40276 4428 40282 4480
rect 41414 4428 41420 4480
rect 41472 4428 41478 4480
rect 41616 4468 41644 4508
rect 41892 4505 41915 4536
rect 41949 4505 41961 4539
rect 41892 4499 41961 4505
rect 41892 4468 41920 4499
rect 41616 4440 41920 4468
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 3421 4267 3479 4273
rect 3421 4233 3433 4267
rect 3467 4264 3479 4267
rect 4062 4264 4068 4276
rect 3467 4236 4068 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 5276 4236 5856 4264
rect 3050 4196 3056 4208
rect 1596 4168 3056 4196
rect 1596 4137 1624 4168
rect 3050 4156 3056 4168
rect 3108 4156 3114 4208
rect 4246 4156 4252 4208
rect 4304 4156 4310 4208
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4097 1639 4131
rect 2501 4131 2559 4137
rect 2501 4128 2513 4131
rect 1581 4091 1639 4097
rect 1688 4100 2513 4128
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1688 4060 1716 4100
rect 2501 4097 2513 4100
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4128 3295 4131
rect 3602 4128 3608 4140
rect 3283 4100 3608 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 3602 4088 3608 4100
rect 3660 4128 3666 4140
rect 3970 4128 3976 4140
rect 3660 4100 3976 4128
rect 3660 4088 3666 4100
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4062 4088 4068 4140
rect 4120 4088 4126 4140
rect 4706 4088 4712 4140
rect 4764 4088 4770 4140
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 5276 4128 5304 4236
rect 5350 4156 5356 4208
rect 5408 4156 5414 4208
rect 5828 4196 5856 4236
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 17586 4264 17592 4276
rect 11756 4236 17592 4264
rect 11756 4224 11762 4236
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 29362 4224 29368 4276
rect 29420 4264 29426 4276
rect 30742 4264 30748 4276
rect 29420 4236 30748 4264
rect 29420 4224 29426 4236
rect 30742 4224 30748 4236
rect 30800 4224 30806 4276
rect 30834 4224 30840 4276
rect 30892 4264 30898 4276
rect 42058 4264 42064 4276
rect 30892 4236 42064 4264
rect 30892 4224 30898 4236
rect 42058 4224 42064 4236
rect 42116 4224 42122 4276
rect 43622 4264 43628 4276
rect 42996 4236 43628 4264
rect 5828 4168 5948 4196
rect 5092 4100 5304 4128
rect 5368 4128 5396 4156
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5368 4100 5733 4128
rect 992 4032 1716 4060
rect 1765 4063 1823 4069
rect 992 4020 998 4032
rect 1765 4029 1777 4063
rect 1811 4029 1823 4063
rect 1765 4023 1823 4029
rect 1118 3952 1124 4004
rect 1176 3992 1182 4004
rect 1780 3992 1808 4023
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 4154 4060 4160 4072
rect 2372 4032 4160 4060
rect 2372 4020 2378 4032
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 5092 4060 5120 4100
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 5920 4128 5948 4168
rect 6840 4168 7052 4196
rect 6840 4128 6868 4168
rect 5920 4100 6868 4128
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 7024 4128 7052 4168
rect 11146 4156 11152 4208
rect 11204 4196 11210 4208
rect 11204 4168 12655 4196
rect 11204 4156 11210 4168
rect 10226 4128 10232 4140
rect 7024 4100 10232 4128
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 11993 4137 12021 4168
rect 11978 4131 12036 4137
rect 11978 4097 11990 4131
rect 12024 4097 12036 4131
rect 11978 4091 12036 4097
rect 12158 4088 12164 4140
rect 12216 4088 12222 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 12391 4131 12449 4137
rect 12391 4097 12403 4131
rect 12437 4128 12449 4131
rect 12526 4128 12532 4140
rect 12437 4100 12532 4128
rect 12437 4097 12449 4100
rect 12391 4091 12449 4097
rect 4724 4032 5120 4060
rect 1176 3964 1808 3992
rect 2685 3995 2743 4001
rect 1176 3952 1182 3964
rect 2685 3961 2697 3995
rect 2731 3992 2743 3995
rect 4724 3992 4752 4032
rect 5166 4020 5172 4072
rect 5224 4060 5230 4072
rect 5353 4063 5411 4069
rect 5353 4060 5365 4063
rect 5224 4032 5365 4060
rect 5224 4020 5230 4032
rect 5353 4029 5365 4032
rect 5399 4029 5411 4063
rect 5353 4023 5411 4029
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4060 5595 4063
rect 7193 4063 7251 4069
rect 7193 4060 7205 4063
rect 5583 4032 7205 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 7193 4029 7205 4032
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 7708 4032 8309 4060
rect 7708 4020 7714 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12268 4060 12296 4091
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12124 4032 12296 4060
rect 12627 4060 12655 4168
rect 17034 4156 17040 4208
rect 17092 4196 17098 4208
rect 17221 4199 17279 4205
rect 17221 4196 17233 4199
rect 17092 4168 17233 4196
rect 17092 4156 17098 4168
rect 17221 4165 17233 4168
rect 17267 4165 17279 4199
rect 17221 4159 17279 4165
rect 17862 4156 17868 4208
rect 17920 4156 17926 4208
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 30374 4196 30380 4208
rect 24912 4168 30380 4196
rect 24912 4156 24918 4168
rect 30374 4156 30380 4168
rect 30432 4196 30438 4208
rect 31754 4196 31760 4208
rect 30432 4168 31064 4196
rect 30432 4156 30438 4168
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 14734 4128 14740 4140
rect 14691 4100 14740 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 14826 4088 14832 4140
rect 14884 4088 14890 4140
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 17954 4128 17960 4140
rect 14976 4100 17960 4128
rect 14976 4088 14982 4100
rect 17954 4088 17960 4100
rect 18012 4128 18018 4140
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 18012 4100 18061 4128
rect 18012 4088 18018 4100
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 19242 4128 19248 4140
rect 18279 4100 19248 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 20346 4088 20352 4140
rect 20404 4088 20410 4140
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 23750 4128 23756 4140
rect 20956 4100 23756 4128
rect 20956 4088 20962 4100
rect 23750 4088 23756 4100
rect 23808 4128 23814 4140
rect 23934 4128 23940 4140
rect 23808 4100 23940 4128
rect 23808 4088 23814 4100
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 29273 4131 29331 4137
rect 29273 4097 29285 4131
rect 29319 4128 29331 4131
rect 29362 4128 29368 4140
rect 29319 4100 29368 4128
rect 29319 4097 29331 4100
rect 29273 4091 29331 4097
rect 29362 4088 29368 4100
rect 29420 4088 29426 4140
rect 29454 4088 29460 4140
rect 29512 4088 29518 4140
rect 29822 4088 29828 4140
rect 29880 4088 29886 4140
rect 30006 4088 30012 4140
rect 30064 4088 30070 4140
rect 31036 4137 31064 4168
rect 31588 4168 31760 4196
rect 30929 4131 30987 4137
rect 30929 4128 30941 4131
rect 30392 4100 30941 4128
rect 15378 4060 15384 4072
rect 12627 4032 15384 4060
rect 12124 4020 12130 4032
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 20533 4063 20591 4069
rect 20533 4060 20545 4063
rect 20312 4032 20545 4060
rect 20312 4020 20318 4032
rect 20533 4029 20545 4032
rect 20579 4029 20591 4063
rect 20533 4023 20591 4029
rect 23842 4020 23848 4072
rect 23900 4020 23906 4072
rect 28902 4020 28908 4072
rect 28960 4060 28966 4072
rect 29549 4063 29607 4069
rect 29549 4060 29561 4063
rect 28960 4032 29561 4060
rect 28960 4020 28966 4032
rect 29549 4029 29561 4032
rect 29595 4029 29607 4063
rect 29549 4023 29607 4029
rect 29641 4063 29699 4069
rect 29641 4029 29653 4063
rect 29687 4060 29699 4063
rect 30098 4060 30104 4072
rect 29687 4032 30104 4060
rect 29687 4029 29699 4032
rect 29641 4023 29699 4029
rect 30098 4020 30104 4032
rect 30156 4020 30162 4072
rect 2731 3964 4752 3992
rect 4801 3995 4859 4001
rect 2731 3961 2743 3964
rect 2685 3955 2743 3961
rect 4801 3961 4813 3995
rect 4847 3992 4859 3995
rect 6822 3992 6828 4004
rect 4847 3964 6828 3992
rect 4847 3961 4859 3964
rect 4801 3955 4859 3961
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 28534 3952 28540 4004
rect 28592 3992 28598 4004
rect 30392 3992 30420 4100
rect 30929 4097 30941 4100
rect 30975 4097 30987 4131
rect 30929 4091 30987 4097
rect 31022 4131 31080 4137
rect 31022 4097 31034 4131
rect 31068 4097 31080 4131
rect 31022 4091 31080 4097
rect 28592 3964 30420 3992
rect 28592 3952 28598 3964
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 5074 3924 5080 3936
rect 2004 3896 5080 3924
rect 2004 3884 2010 3896
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 7926 3924 7932 3936
rect 5868 3896 7932 3924
rect 5868 3884 5874 3896
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 12434 3924 12440 3936
rect 8444 3896 12440 3924
rect 8444 3884 8450 3896
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 13538 3924 13544 3936
rect 12676 3896 13544 3924
rect 12676 3884 12682 3896
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 14642 3884 14648 3936
rect 14700 3884 14706 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 16632 3896 17325 3924
rect 16632 3884 16638 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 24026 3884 24032 3936
rect 24084 3924 24090 3936
rect 24121 3927 24179 3933
rect 24121 3924 24133 3927
rect 24084 3896 24133 3924
rect 24084 3884 24090 3896
rect 24121 3893 24133 3896
rect 24167 3893 24179 3927
rect 24121 3887 24179 3893
rect 27614 3884 27620 3936
rect 27672 3924 27678 3936
rect 29270 3924 29276 3936
rect 27672 3896 29276 3924
rect 27672 3884 27678 3896
rect 29270 3884 29276 3896
rect 29328 3884 29334 3936
rect 30944 3924 30972 4091
rect 31202 4088 31208 4140
rect 31260 4088 31266 4140
rect 31294 4088 31300 4140
rect 31352 4088 31358 4140
rect 31435 4131 31493 4137
rect 31435 4097 31447 4131
rect 31481 4128 31493 4131
rect 31588 4128 31616 4168
rect 31754 4156 31760 4168
rect 31812 4156 31818 4208
rect 34514 4156 34520 4208
rect 34572 4196 34578 4208
rect 34701 4199 34759 4205
rect 34701 4196 34713 4199
rect 34572 4168 34713 4196
rect 34572 4156 34578 4168
rect 34701 4165 34713 4168
rect 34747 4165 34759 4199
rect 34701 4159 34759 4165
rect 38654 4156 38660 4208
rect 38712 4196 38718 4208
rect 38841 4199 38899 4205
rect 38841 4196 38853 4199
rect 38712 4168 38853 4196
rect 38712 4156 38718 4168
rect 38841 4165 38853 4168
rect 38887 4165 38899 4199
rect 38841 4159 38899 4165
rect 41782 4156 41788 4208
rect 41840 4196 41846 4208
rect 42996 4205 43024 4236
rect 43622 4224 43628 4236
rect 43680 4224 43686 4276
rect 43990 4224 43996 4276
rect 44048 4224 44054 4276
rect 42981 4199 43039 4205
rect 42981 4196 42993 4199
rect 41840 4168 42993 4196
rect 41840 4156 41846 4168
rect 42981 4165 42993 4168
rect 43027 4165 43039 4199
rect 42981 4159 43039 4165
rect 43070 4156 43076 4208
rect 43128 4205 43134 4208
rect 43128 4199 43157 4205
rect 43145 4165 43157 4199
rect 43128 4159 43157 4165
rect 43128 4156 43134 4159
rect 44358 4156 44364 4208
rect 44416 4156 44422 4208
rect 45557 4199 45615 4205
rect 45557 4165 45569 4199
rect 45603 4196 45615 4199
rect 46842 4196 46848 4208
rect 45603 4168 46848 4196
rect 45603 4165 45615 4168
rect 45557 4159 45615 4165
rect 33045 4131 33103 4137
rect 33045 4128 33057 4131
rect 31481 4100 31616 4128
rect 31726 4100 33057 4128
rect 31481 4097 31493 4100
rect 31435 4091 31493 4097
rect 31726 4060 31754 4100
rect 33045 4097 33057 4100
rect 33091 4097 33103 4131
rect 33045 4091 33103 4097
rect 38930 4088 38936 4140
rect 38988 4128 38994 4140
rect 39025 4131 39083 4137
rect 39025 4128 39037 4131
rect 38988 4100 39037 4128
rect 38988 4088 38994 4100
rect 39025 4097 39037 4100
rect 39071 4097 39083 4131
rect 42797 4131 42855 4137
rect 42797 4128 42809 4131
rect 39025 4091 39083 4097
rect 42720 4100 42809 4128
rect 31588 4032 31754 4060
rect 32861 4063 32919 4069
rect 31588 4001 31616 4032
rect 32861 4029 32873 4063
rect 32907 4060 32919 4063
rect 33134 4060 33140 4072
rect 32907 4032 33140 4060
rect 32907 4029 32919 4032
rect 32861 4023 32919 4029
rect 33134 4020 33140 4032
rect 33192 4020 33198 4072
rect 34698 4020 34704 4072
rect 34756 4060 34762 4072
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34756 4032 34897 4060
rect 34756 4020 34762 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 34885 4023 34943 4029
rect 36354 4020 36360 4072
rect 36412 4060 36418 4072
rect 39114 4060 39120 4072
rect 36412 4032 39120 4060
rect 36412 4020 36418 4032
rect 39114 4020 39120 4032
rect 39172 4020 39178 4072
rect 31573 3995 31631 4001
rect 31573 3961 31585 3995
rect 31619 3961 31631 3995
rect 34606 3992 34612 4004
rect 31573 3955 31631 3961
rect 31726 3964 34612 3992
rect 31726 3924 31754 3964
rect 34606 3952 34612 3964
rect 34664 3952 34670 4004
rect 42720 3992 42748 4100
rect 42797 4097 42809 4100
rect 42843 4097 42855 4131
rect 42797 4091 42855 4097
rect 42886 4088 42892 4140
rect 42944 4088 42950 4140
rect 44453 4131 44511 4137
rect 44453 4097 44465 4131
rect 44499 4128 44511 4131
rect 45572 4128 45600 4159
rect 46842 4156 46848 4168
rect 46900 4156 46906 4208
rect 44499 4100 45600 4128
rect 45649 4131 45707 4137
rect 44499 4097 44511 4100
rect 44453 4091 44511 4097
rect 45649 4097 45661 4131
rect 45695 4128 45707 4131
rect 54846 4128 54852 4140
rect 45695 4100 54852 4128
rect 45695 4097 45707 4100
rect 45649 4091 45707 4097
rect 42978 4020 42984 4072
rect 43036 4060 43042 4072
rect 43257 4063 43315 4069
rect 43257 4060 43269 4063
rect 43036 4032 43269 4060
rect 43036 4020 43042 4032
rect 43257 4029 43269 4032
rect 43303 4029 43315 4063
rect 43257 4023 43315 4029
rect 43346 4020 43352 4072
rect 43404 4060 43410 4072
rect 44468 4060 44496 4091
rect 43404 4032 44496 4060
rect 43404 4020 43410 4032
rect 44634 4020 44640 4072
rect 44692 4060 44698 4072
rect 45741 4063 45799 4069
rect 44692 4032 45600 4060
rect 44692 4020 44698 4032
rect 45189 3995 45247 4001
rect 45189 3992 45201 3995
rect 42720 3964 45201 3992
rect 45189 3961 45201 3964
rect 45235 3961 45247 3995
rect 45572 3992 45600 4032
rect 45741 4029 45753 4063
rect 45787 4029 45799 4063
rect 45741 4023 45799 4029
rect 45756 3992 45784 4023
rect 45572 3964 45784 3992
rect 45189 3955 45247 3961
rect 30944 3896 31754 3924
rect 33229 3927 33287 3933
rect 33229 3893 33241 3927
rect 33275 3924 33287 3927
rect 33962 3924 33968 3936
rect 33275 3896 33968 3924
rect 33275 3893 33287 3896
rect 33229 3887 33287 3893
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 42610 3884 42616 3936
rect 42668 3884 42674 3936
rect 43254 3884 43260 3936
rect 43312 3924 43318 3936
rect 45848 3924 45876 4100
rect 54846 4088 54852 4100
rect 54904 4088 54910 4140
rect 43312 3896 45876 3924
rect 43312 3884 43318 3896
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 1946 3680 1952 3732
rect 2004 3680 2010 3732
rect 2685 3723 2743 3729
rect 2685 3689 2697 3723
rect 2731 3720 2743 3723
rect 4614 3720 4620 3732
rect 2731 3692 4620 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 4948 3692 7205 3720
rect 4948 3680 4954 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 10686 3720 10692 3732
rect 7193 3683 7251 3689
rect 8588 3692 10692 3720
rect 934 3612 940 3664
rect 992 3652 998 3664
rect 4062 3652 4068 3664
rect 992 3624 4068 3652
rect 992 3612 998 3624
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 4801 3655 4859 3661
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 5810 3652 5816 3664
rect 4847 3624 5816 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 5810 3612 5816 3624
rect 5868 3612 5874 3664
rect 6549 3655 6607 3661
rect 6549 3621 6561 3655
rect 6595 3652 6607 3655
rect 8588 3652 8616 3692
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 12066 3720 12072 3732
rect 11747 3692 12072 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 13170 3720 13176 3732
rect 12492 3692 13176 3720
rect 12492 3680 12498 3692
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 17310 3720 17316 3732
rect 16899 3692 17316 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 17957 3723 18015 3729
rect 17957 3689 17969 3723
rect 18003 3720 18015 3723
rect 18046 3720 18052 3732
rect 18003 3692 18052 3720
rect 18003 3689 18015 3692
rect 17957 3683 18015 3689
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 21085 3723 21143 3729
rect 21085 3720 21097 3723
rect 20220 3692 21097 3720
rect 20220 3680 20226 3692
rect 21085 3689 21097 3692
rect 21131 3689 21143 3723
rect 21085 3683 21143 3689
rect 28718 3680 28724 3732
rect 28776 3720 28782 3732
rect 30193 3723 30251 3729
rect 30193 3720 30205 3723
rect 28776 3692 30205 3720
rect 28776 3680 28782 3692
rect 30193 3689 30205 3692
rect 30239 3689 30251 3723
rect 30193 3683 30251 3689
rect 30926 3680 30932 3732
rect 30984 3720 30990 3732
rect 31386 3720 31392 3732
rect 30984 3692 31392 3720
rect 30984 3680 30990 3692
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 39485 3723 39543 3729
rect 39485 3689 39497 3723
rect 39531 3720 39543 3723
rect 40034 3720 40040 3732
rect 39531 3692 40040 3720
rect 39531 3689 39543 3692
rect 39485 3683 39543 3689
rect 40034 3680 40040 3692
rect 40092 3680 40098 3732
rect 42429 3723 42487 3729
rect 42429 3689 42441 3723
rect 42475 3720 42487 3723
rect 43346 3720 43352 3732
rect 42475 3692 43352 3720
rect 42475 3689 42487 3692
rect 42429 3683 42487 3689
rect 43346 3680 43352 3692
rect 43404 3680 43410 3732
rect 10410 3652 10416 3664
rect 6595 3624 8616 3652
rect 10244 3624 10416 3652
rect 6595 3621 6607 3624
rect 6549 3615 6607 3621
rect 5166 3584 5172 3596
rect 4632 3556 5172 3584
rect 2498 3476 2504 3528
rect 2556 3476 2562 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3694 3516 3700 3528
rect 3467 3488 3700 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 4632 3525 4660 3556
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 10244 3593 10272 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 12158 3612 12164 3664
rect 12216 3652 12222 3664
rect 13354 3652 13360 3664
rect 12216 3624 13360 3652
rect 12216 3612 12222 3624
rect 13354 3612 13360 3624
rect 13412 3652 13418 3664
rect 16114 3652 16120 3664
rect 13412 3624 16120 3652
rect 13412 3612 13418 3624
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 20806 3652 20812 3664
rect 16224 3624 20812 3652
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 6512 3556 7757 3584
rect 6512 3544 6518 3556
rect 7745 3553 7757 3556
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3553 10287 3587
rect 11514 3584 11520 3596
rect 10229 3547 10287 3553
rect 10428 3556 11520 3584
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 4982 3476 4988 3528
rect 5040 3516 5046 3528
rect 5445 3519 5503 3525
rect 5445 3516 5457 3519
rect 5040 3488 5457 3516
rect 5040 3476 5046 3488
rect 5445 3485 5457 3488
rect 5491 3485 5503 3519
rect 5445 3479 5503 3485
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 5736 3488 7113 3516
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 1673 3451 1731 3457
rect 1673 3448 1685 3451
rect 1084 3420 1685 3448
rect 1084 3408 1090 3420
rect 1673 3417 1685 3420
rect 1719 3417 1731 3451
rect 2516 3448 2544 3476
rect 3602 3448 3608 3460
rect 2516 3420 3608 3448
rect 1673 3411 1731 3417
rect 3602 3408 3608 3420
rect 3660 3408 3666 3460
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 5736 3448 5764 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 9122 3476 9128 3528
rect 9180 3516 9186 3528
rect 10428 3525 10456 3556
rect 11514 3544 11520 3556
rect 11572 3584 11578 3596
rect 11790 3584 11796 3596
rect 11572 3556 11796 3584
rect 11572 3544 11578 3556
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 16224 3584 16252 3624
rect 11940 3556 16252 3584
rect 11940 3544 11946 3556
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9180 3488 10425 3516
rect 9180 3476 9186 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 10413 3479 10471 3485
rect 10520 3488 12265 3516
rect 4120 3420 5764 3448
rect 4120 3408 4126 3420
rect 5994 3408 6000 3460
rect 6052 3448 6058 3460
rect 6365 3451 6423 3457
rect 6365 3448 6377 3451
rect 6052 3420 6377 3448
rect 6052 3408 6058 3420
rect 6365 3417 6377 3420
rect 6411 3417 6423 3451
rect 6365 3411 6423 3417
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 10520 3448 10548 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 12802 3516 12808 3528
rect 12667 3488 12808 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 9456 3420 10548 3448
rect 10597 3451 10655 3457
rect 9456 3408 9462 3420
rect 10597 3417 10609 3451
rect 10643 3448 10655 3451
rect 10643 3420 11468 3448
rect 10643 3417 10655 3420
rect 10597 3411 10655 3417
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 5810 3340 5816 3392
rect 5868 3340 5874 3392
rect 11440 3380 11468 3420
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 11609 3451 11667 3457
rect 11609 3448 11621 3451
rect 11572 3420 11621 3448
rect 11572 3408 11578 3420
rect 11609 3417 11621 3420
rect 11655 3417 11667 3451
rect 11609 3411 11667 3417
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 12452 3448 12480 3479
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 13096 3525 13124 3556
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13228 3488 13273 3516
rect 13228 3476 13234 3488
rect 13354 3476 13360 3528
rect 13412 3476 13418 3528
rect 13538 3476 13544 3528
rect 13596 3525 13602 3528
rect 16224 3525 16252 3556
rect 13596 3519 13645 3525
rect 13596 3485 13599 3519
rect 13633 3516 13645 3519
rect 16209 3519 16267 3525
rect 13633 3488 14688 3516
rect 13633 3485 13645 3488
rect 13596 3479 13645 3485
rect 13596 3476 13602 3479
rect 11848 3420 12480 3448
rect 13449 3451 13507 3457
rect 11848 3408 11854 3420
rect 13449 3417 13461 3451
rect 13495 3448 13507 3451
rect 13495 3420 14044 3448
rect 13495 3417 13507 3420
rect 13449 3411 13507 3417
rect 13630 3380 13636 3392
rect 11440 3352 13636 3380
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13722 3340 13728 3392
rect 13780 3340 13786 3392
rect 14016 3380 14044 3420
rect 14274 3408 14280 3460
rect 14332 3448 14338 3460
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 14332 3420 14473 3448
rect 14332 3408 14338 3420
rect 14461 3417 14473 3420
rect 14507 3417 14519 3451
rect 14461 3411 14519 3417
rect 14553 3383 14611 3389
rect 14553 3380 14565 3383
rect 14016 3352 14565 3380
rect 14553 3349 14565 3352
rect 14599 3349 14611 3383
rect 14660 3380 14688 3488
rect 16209 3485 16221 3519
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 16574 3516 16580 3528
rect 16632 3525 16638 3528
rect 16758 3525 16764 3528
rect 16356 3488 16401 3516
rect 16543 3488 16580 3516
rect 16356 3476 16362 3488
rect 16574 3476 16580 3488
rect 16632 3479 16643 3525
rect 16715 3519 16764 3525
rect 16715 3485 16727 3519
rect 16761 3485 16764 3519
rect 16715 3479 16764 3485
rect 16632 3476 16638 3479
rect 16758 3476 16764 3479
rect 16816 3476 16822 3528
rect 17328 3525 17356 3624
rect 19705 3587 19763 3593
rect 19705 3584 19717 3587
rect 18616 3556 19717 3584
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17862 3525 17868 3528
rect 17819 3519 17868 3525
rect 17460 3488 17505 3516
rect 17460 3476 17466 3488
rect 17819 3485 17831 3519
rect 17865 3485 17868 3519
rect 17819 3479 17868 3485
rect 17862 3476 17868 3479
rect 17920 3476 17926 3528
rect 16114 3408 16120 3460
rect 16172 3448 16178 3460
rect 16485 3451 16543 3457
rect 16485 3448 16497 3451
rect 16172 3420 16497 3448
rect 16172 3408 16178 3420
rect 16485 3417 16497 3420
rect 16531 3448 16543 3451
rect 17589 3451 17647 3457
rect 17589 3448 17601 3451
rect 16531 3420 17601 3448
rect 16531 3417 16543 3420
rect 16485 3411 16543 3417
rect 17589 3417 17601 3420
rect 17635 3417 17647 3451
rect 17589 3411 17647 3417
rect 17681 3451 17739 3457
rect 17681 3417 17693 3451
rect 17727 3448 17739 3451
rect 18616 3448 18644 3556
rect 19705 3553 19717 3556
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19426 3516 19432 3528
rect 19024 3488 19432 3516
rect 19024 3476 19030 3488
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 20456 3525 20484 3624
rect 20806 3612 20812 3624
rect 20864 3612 20870 3664
rect 27154 3612 27160 3664
rect 27212 3652 27218 3664
rect 28902 3652 28908 3664
rect 27212 3624 28908 3652
rect 27212 3612 27218 3624
rect 28902 3612 28908 3624
rect 28960 3612 28966 3664
rect 29181 3655 29239 3661
rect 29181 3621 29193 3655
rect 29227 3621 29239 3655
rect 29181 3615 29239 3621
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 22186 3584 22192 3596
rect 20680 3556 22192 3584
rect 20680 3544 20686 3556
rect 20441 3519 20499 3525
rect 20441 3485 20453 3519
rect 20487 3485 20499 3519
rect 20441 3479 20499 3485
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20906 3519 20964 3525
rect 20588 3488 20633 3516
rect 20588 3476 20594 3488
rect 20906 3485 20918 3519
rect 20952 3516 20964 3519
rect 21008 3516 21036 3556
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 27614 3544 27620 3596
rect 27672 3544 27678 3596
rect 29196 3584 29224 3615
rect 30098 3612 30104 3664
rect 30156 3652 30162 3664
rect 31478 3652 31484 3664
rect 30156 3624 31484 3652
rect 30156 3612 30162 3624
rect 27816 3556 29224 3584
rect 20952 3488 21036 3516
rect 20952 3485 20964 3488
rect 20906 3479 20964 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 21140 3488 22661 3516
rect 21140 3476 21146 3488
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 23658 3476 23664 3528
rect 23716 3516 23722 3528
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 23716 3488 23765 3516
rect 23716 3476 23722 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 23753 3479 23811 3485
rect 24026 3476 24032 3528
rect 24084 3476 24090 3528
rect 25777 3519 25835 3525
rect 25777 3485 25789 3519
rect 25823 3516 25835 3519
rect 25866 3516 25872 3528
rect 25823 3488 25872 3516
rect 25823 3485 25835 3488
rect 25777 3479 25835 3485
rect 25866 3476 25872 3488
rect 25924 3476 25930 3528
rect 27816 3525 27844 3556
rect 29454 3544 29460 3596
rect 29512 3584 29518 3596
rect 29512 3556 30972 3584
rect 29512 3544 29518 3556
rect 30944 3528 30972 3556
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3485 27859 3519
rect 27801 3479 27859 3485
rect 28534 3476 28540 3528
rect 28592 3476 28598 3528
rect 28630 3519 28688 3525
rect 28630 3485 28642 3519
rect 28676 3485 28688 3519
rect 28630 3479 28688 3485
rect 17727 3420 18644 3448
rect 17727 3417 17739 3420
rect 17681 3411 17739 3417
rect 16758 3380 16764 3392
rect 14660 3352 16764 3380
rect 14553 3343 14611 3349
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 17604 3380 17632 3411
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 19521 3451 19579 3457
rect 19521 3448 19533 3451
rect 19392 3420 19533 3448
rect 19392 3408 19398 3420
rect 19521 3417 19533 3420
rect 19567 3417 19579 3451
rect 19521 3411 19579 3417
rect 20717 3451 20775 3457
rect 20717 3417 20729 3451
rect 20763 3417 20775 3451
rect 20717 3411 20775 3417
rect 20809 3451 20867 3457
rect 20809 3417 20821 3451
rect 20855 3448 20867 3451
rect 20855 3420 21404 3448
rect 20855 3417 20867 3420
rect 20809 3411 20867 3417
rect 20732 3380 20760 3411
rect 20990 3380 20996 3392
rect 17604 3352 20996 3380
rect 20990 3340 20996 3352
rect 21048 3380 21054 3392
rect 21266 3380 21272 3392
rect 21048 3352 21272 3380
rect 21048 3340 21054 3352
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 21376 3380 21404 3420
rect 21634 3408 21640 3460
rect 21692 3448 21698 3460
rect 21821 3451 21879 3457
rect 21821 3448 21833 3451
rect 21692 3420 21833 3448
rect 21692 3408 21698 3420
rect 21821 3417 21833 3420
rect 21867 3417 21879 3451
rect 21821 3411 21879 3417
rect 22554 3408 22560 3460
rect 22612 3448 22618 3460
rect 22925 3451 22983 3457
rect 22925 3448 22937 3451
rect 22612 3420 22937 3448
rect 22612 3408 22618 3420
rect 22925 3417 22937 3420
rect 22971 3417 22983 3451
rect 22925 3411 22983 3417
rect 23842 3408 23848 3460
rect 23900 3448 23906 3460
rect 26044 3451 26102 3457
rect 23900 3420 26004 3448
rect 23900 3408 23906 3420
rect 21913 3383 21971 3389
rect 21913 3380 21925 3383
rect 21376 3352 21925 3380
rect 21913 3349 21925 3352
rect 21959 3349 21971 3383
rect 21913 3343 21971 3349
rect 23566 3340 23572 3392
rect 23624 3340 23630 3392
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 25406 3380 25412 3392
rect 23983 3352 25412 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 25406 3340 25412 3352
rect 25464 3340 25470 3392
rect 25976 3380 26004 3420
rect 26044 3417 26056 3451
rect 26090 3448 26102 3451
rect 27985 3451 28043 3457
rect 27985 3448 27997 3451
rect 26090 3420 27997 3448
rect 26090 3417 26102 3420
rect 26044 3411 26102 3417
rect 27985 3417 27997 3420
rect 28031 3417 28043 3451
rect 27985 3411 28043 3417
rect 28644 3380 28672 3479
rect 28902 3476 28908 3528
rect 28960 3476 28966 3528
rect 29043 3519 29101 3525
rect 29043 3485 29055 3519
rect 29089 3516 29101 3519
rect 29089 3488 30420 3516
rect 29089 3485 29101 3488
rect 29043 3479 29101 3485
rect 28813 3451 28871 3457
rect 28813 3417 28825 3451
rect 28859 3448 28871 3451
rect 29914 3448 29920 3460
rect 28859 3420 29920 3448
rect 28859 3417 28871 3420
rect 28813 3411 28871 3417
rect 29914 3408 29920 3420
rect 29972 3408 29978 3460
rect 30101 3451 30159 3457
rect 30101 3417 30113 3451
rect 30147 3448 30159 3451
rect 30282 3448 30288 3460
rect 30147 3420 30288 3448
rect 30147 3417 30159 3420
rect 30101 3411 30159 3417
rect 30282 3408 30288 3420
rect 30340 3408 30346 3460
rect 30006 3380 30012 3392
rect 25976 3352 30012 3380
rect 30006 3340 30012 3352
rect 30064 3340 30070 3392
rect 30392 3380 30420 3488
rect 30558 3476 30564 3528
rect 30616 3516 30622 3528
rect 30742 3516 30748 3528
rect 30616 3488 30748 3516
rect 30616 3476 30622 3488
rect 30742 3476 30748 3488
rect 30800 3476 30806 3528
rect 30926 3476 30932 3528
rect 30984 3476 30990 3528
rect 31021 3519 31079 3525
rect 31021 3485 31033 3519
rect 31067 3485 31079 3519
rect 31021 3479 31079 3485
rect 31113 3519 31171 3525
rect 31113 3485 31125 3519
rect 31159 3516 31171 3519
rect 31220 3516 31248 3624
rect 31478 3612 31484 3624
rect 31536 3612 31542 3664
rect 40405 3655 40463 3661
rect 40405 3621 40417 3655
rect 40451 3652 40463 3655
rect 40494 3652 40500 3664
rect 40451 3624 40500 3652
rect 40451 3621 40463 3624
rect 40405 3615 40463 3621
rect 40494 3612 40500 3624
rect 40552 3612 40558 3664
rect 31938 3544 31944 3596
rect 31996 3544 32002 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 35894 3584 35900 3596
rect 33928 3556 35900 3584
rect 33928 3544 33934 3556
rect 35894 3544 35900 3556
rect 35952 3544 35958 3596
rect 31159 3488 31248 3516
rect 31297 3519 31355 3525
rect 31159 3485 31171 3488
rect 31113 3479 31171 3485
rect 31297 3485 31309 3519
rect 31343 3516 31355 3519
rect 31386 3516 31392 3528
rect 31343 3488 31392 3516
rect 31343 3485 31355 3488
rect 31297 3479 31355 3485
rect 30466 3408 30472 3460
rect 30524 3448 30530 3460
rect 31036 3448 31064 3479
rect 31386 3476 31392 3488
rect 31444 3516 31450 3528
rect 35161 3519 35219 3525
rect 31444 3488 32332 3516
rect 31444 3476 31450 3488
rect 31202 3448 31208 3460
rect 30524 3420 31208 3448
rect 30524 3408 30530 3420
rect 31202 3408 31208 3420
rect 31260 3408 31266 3460
rect 31481 3451 31539 3457
rect 31481 3417 31493 3451
rect 31527 3448 31539 3451
rect 32186 3451 32244 3457
rect 32186 3448 32198 3451
rect 31527 3420 32198 3448
rect 31527 3417 31539 3420
rect 31481 3411 31539 3417
rect 32186 3417 32198 3420
rect 32232 3417 32244 3451
rect 32186 3411 32244 3417
rect 31754 3380 31760 3392
rect 30392 3352 31760 3380
rect 31754 3340 31760 3352
rect 31812 3380 31818 3392
rect 32030 3380 32036 3392
rect 31812 3352 32036 3380
rect 31812 3340 31818 3352
rect 32030 3340 32036 3352
rect 32088 3340 32094 3392
rect 32304 3380 32332 3488
rect 35161 3485 35173 3519
rect 35207 3485 35219 3519
rect 35161 3479 35219 3485
rect 35253 3519 35311 3525
rect 35253 3485 35265 3519
rect 35299 3516 35311 3519
rect 35526 3516 35532 3528
rect 35299 3488 35532 3516
rect 35299 3485 35311 3488
rect 35253 3479 35311 3485
rect 35176 3448 35204 3479
rect 35526 3476 35532 3488
rect 35584 3476 35590 3528
rect 35912 3516 35940 3544
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 35912 3488 38117 3516
rect 38105 3485 38117 3488
rect 38151 3516 38163 3519
rect 38194 3516 38200 3528
rect 38151 3488 38200 3516
rect 38151 3485 38163 3488
rect 38105 3479 38163 3485
rect 38194 3476 38200 3488
rect 38252 3476 38258 3528
rect 38372 3519 38430 3525
rect 38372 3485 38384 3519
rect 38418 3516 38430 3519
rect 38746 3516 38752 3528
rect 38418 3488 38752 3516
rect 38418 3485 38430 3488
rect 38372 3479 38430 3485
rect 38746 3476 38752 3488
rect 38804 3476 38810 3528
rect 41046 3476 41052 3528
rect 41104 3476 41110 3528
rect 41316 3519 41374 3525
rect 41316 3485 41328 3519
rect 41362 3516 41374 3519
rect 42610 3516 42616 3528
rect 41362 3488 42616 3516
rect 41362 3485 41374 3488
rect 41316 3479 41374 3485
rect 42610 3476 42616 3488
rect 42668 3476 42674 3528
rect 44358 3476 44364 3528
rect 44416 3516 44422 3528
rect 57149 3519 57207 3525
rect 57149 3516 57161 3519
rect 44416 3488 57161 3516
rect 44416 3476 44422 3488
rect 57149 3485 57161 3488
rect 57195 3485 57207 3519
rect 57149 3479 57207 3485
rect 35342 3448 35348 3460
rect 35176 3420 35348 3448
rect 35342 3408 35348 3420
rect 35400 3408 35406 3460
rect 35437 3451 35495 3457
rect 35437 3417 35449 3451
rect 35483 3448 35495 3451
rect 36142 3451 36200 3457
rect 36142 3448 36154 3451
rect 35483 3420 36154 3448
rect 35483 3417 35495 3420
rect 35437 3411 35495 3417
rect 36142 3417 36154 3420
rect 36188 3417 36200 3451
rect 36142 3411 36200 3417
rect 40034 3408 40040 3460
rect 40092 3448 40098 3460
rect 40221 3451 40279 3457
rect 40221 3448 40233 3451
rect 40092 3420 40233 3448
rect 40092 3408 40098 3420
rect 40221 3417 40233 3420
rect 40267 3417 40279 3451
rect 40221 3411 40279 3417
rect 57054 3408 57060 3460
rect 57112 3448 57118 3460
rect 57425 3451 57483 3457
rect 57425 3448 57437 3451
rect 57112 3420 57437 3448
rect 57112 3408 57118 3420
rect 57425 3417 57437 3420
rect 57471 3417 57483 3451
rect 57425 3411 57483 3417
rect 33321 3383 33379 3389
rect 33321 3380 33333 3383
rect 32304 3352 33333 3380
rect 33321 3349 33333 3352
rect 33367 3380 33379 3383
rect 34698 3380 34704 3392
rect 33367 3352 34704 3380
rect 33367 3349 33379 3352
rect 33321 3343 33379 3349
rect 34698 3340 34704 3352
rect 34756 3340 34762 3392
rect 37274 3340 37280 3392
rect 37332 3340 37338 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 4890 3176 4896 3188
rect 1596 3148 4896 3176
rect 1596 3049 1624 3148
rect 4890 3136 4896 3148
rect 4948 3176 4954 3188
rect 4985 3179 5043 3185
rect 4985 3176 4997 3179
rect 4948 3148 4997 3176
rect 4948 3136 4954 3148
rect 4985 3145 4997 3148
rect 5031 3145 5043 3179
rect 4985 3139 5043 3145
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 9766 3176 9772 3188
rect 5868 3148 9772 3176
rect 5868 3136 5874 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 21453 3179 21511 3185
rect 10008 3148 13032 3176
rect 10008 3136 10014 3148
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 6362 3108 6368 3120
rect 1912 3080 6368 3108
rect 1912 3068 1918 3080
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 8386 3108 8392 3120
rect 7024 3080 8392 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2222 3000 2228 3052
rect 2280 3040 2286 3052
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2280 3012 2697 3040
rect 2280 3000 2286 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 3872 3043 3930 3049
rect 3872 3009 3884 3043
rect 3918 3040 3930 3043
rect 4430 3040 4436 3052
rect 3918 3012 4436 3040
rect 3918 3009 3930 3012
rect 3872 3003 3930 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5316 3012 5457 3040
rect 5316 3000 5322 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 7024 3049 7052 3080
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 8481 3111 8539 3117
rect 8481 3077 8493 3111
rect 8527 3108 8539 3111
rect 8662 3108 8668 3120
rect 8527 3080 8668 3108
rect 8527 3077 8539 3080
rect 8481 3071 8539 3077
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 10042 3068 10048 3120
rect 10100 3068 10106 3120
rect 10778 3068 10784 3120
rect 10836 3068 10842 3120
rect 7009 3043 7067 3049
rect 5684 3012 6868 3040
rect 5684 3000 5690 3012
rect 934 2932 940 2984
rect 992 2972 998 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 992 2944 1777 2972
rect 992 2932 998 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3234 2972 3240 2984
rect 3007 2944 3240 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 5810 2864 5816 2916
rect 5868 2864 5874 2916
rect 6840 2904 6868 3012
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8754 3040 8760 3052
rect 8343 3012 8760 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 9769 3046 9827 3049
rect 9769 3043 9996 3046
rect 9769 3009 9781 3043
rect 9815 3040 9996 3043
rect 10796 3040 10824 3068
rect 9815 3018 10824 3040
rect 9815 3009 9827 3018
rect 9968 3012 10824 3018
rect 9769 3003 9827 3009
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 13004 3049 13032 3148
rect 18064 3148 20116 3176
rect 13630 3068 13636 3120
rect 13688 3108 13694 3120
rect 14176 3111 14234 3117
rect 13688 3080 14044 3108
rect 13688 3068 13694 3080
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 11020 3012 12357 3040
rect 11020 3000 11026 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13504 3012 13921 3040
rect 13504 3000 13510 3012
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 14016 3040 14044 3080
rect 14176 3077 14188 3111
rect 14222 3108 14234 3111
rect 14642 3108 14648 3120
rect 14222 3080 14648 3108
rect 14222 3077 14234 3080
rect 14176 3071 14234 3077
rect 14642 3068 14648 3080
rect 14700 3068 14706 3120
rect 18064 3049 18092 3148
rect 19236 3111 19294 3117
rect 19236 3077 19248 3111
rect 19282 3108 19294 3111
rect 19978 3108 19984 3120
rect 19282 3080 19984 3108
rect 19282 3077 19294 3080
rect 19236 3071 19294 3077
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 20088 3108 20116 3148
rect 21453 3145 21465 3179
rect 21499 3176 21511 3179
rect 21542 3176 21548 3188
rect 21499 3148 21548 3176
rect 21499 3145 21511 3148
rect 21453 3139 21511 3145
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 23842 3176 23848 3188
rect 22066 3148 23848 3176
rect 22066 3108 22094 3148
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 23934 3136 23940 3188
rect 23992 3136 23998 3188
rect 26142 3136 26148 3188
rect 26200 3176 26206 3188
rect 27433 3179 27491 3185
rect 27433 3176 27445 3179
rect 26200 3148 27445 3176
rect 26200 3136 26206 3148
rect 27433 3145 27445 3148
rect 27479 3145 27491 3179
rect 27433 3139 27491 3145
rect 27798 3136 27804 3188
rect 27856 3176 27862 3188
rect 28169 3179 28227 3185
rect 28169 3176 28181 3179
rect 27856 3148 28181 3176
rect 27856 3136 27862 3148
rect 28169 3145 28181 3148
rect 28215 3145 28227 3179
rect 28169 3139 28227 3145
rect 28994 3136 29000 3188
rect 29052 3136 29058 3188
rect 30006 3136 30012 3188
rect 30064 3176 30070 3188
rect 30101 3179 30159 3185
rect 30101 3176 30113 3179
rect 30064 3148 30113 3176
rect 30064 3136 30070 3148
rect 30101 3145 30113 3148
rect 30147 3145 30159 3179
rect 30101 3139 30159 3145
rect 30466 3136 30472 3188
rect 30524 3176 30530 3188
rect 35253 3179 35311 3185
rect 35253 3176 35265 3179
rect 30524 3148 35265 3176
rect 30524 3136 30530 3148
rect 35253 3145 35265 3148
rect 35299 3145 35311 3179
rect 35253 3139 35311 3145
rect 35710 3136 35716 3188
rect 35768 3176 35774 3188
rect 37645 3179 37703 3185
rect 37645 3176 37657 3179
rect 35768 3148 37657 3176
rect 35768 3136 35774 3148
rect 37645 3145 37657 3148
rect 37691 3145 37703 3179
rect 37645 3139 37703 3145
rect 39114 3136 39120 3188
rect 39172 3176 39178 3188
rect 39577 3179 39635 3185
rect 39577 3176 39589 3179
rect 39172 3148 39589 3176
rect 39172 3136 39178 3148
rect 39577 3145 39589 3148
rect 39623 3145 39635 3179
rect 39577 3139 39635 3145
rect 41230 3136 41236 3188
rect 41288 3176 41294 3188
rect 42797 3179 42855 3185
rect 42797 3176 42809 3179
rect 41288 3148 42809 3176
rect 41288 3136 41294 3148
rect 42797 3145 42809 3148
rect 42843 3145 42855 3179
rect 42797 3139 42855 3145
rect 43162 3136 43168 3188
rect 43220 3176 43226 3188
rect 43533 3179 43591 3185
rect 43533 3176 43545 3179
rect 43220 3148 43545 3176
rect 43220 3136 43226 3148
rect 43533 3145 43545 3148
rect 43579 3145 43591 3179
rect 43533 3139 43591 3145
rect 44450 3136 44456 3188
rect 44508 3136 44514 3188
rect 44910 3136 44916 3188
rect 44968 3176 44974 3188
rect 45833 3179 45891 3185
rect 45833 3176 45845 3179
rect 44968 3148 45845 3176
rect 44968 3136 44974 3148
rect 45833 3145 45845 3148
rect 45879 3145 45891 3179
rect 45833 3139 45891 3145
rect 47946 3136 47952 3188
rect 48004 3136 48010 3188
rect 54110 3136 54116 3188
rect 54168 3136 54174 3188
rect 55950 3136 55956 3188
rect 56008 3136 56014 3188
rect 25866 3108 25872 3120
rect 20088 3080 22094 3108
rect 22572 3080 25872 3108
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 14016 3012 15853 3040
rect 13909 3003 13967 3009
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 6972 2944 7205 2972
rect 6972 2932 6978 2944
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8536 2944 8953 2972
rect 8536 2932 8542 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 9140 2904 9168 3000
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 6840 2876 9168 2904
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 10796 2904 10824 2935
rect 11238 2932 11244 2984
rect 11296 2972 11302 2984
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 11296 2944 12173 2972
rect 11296 2932 11302 2944
rect 12161 2941 12173 2944
rect 12207 2941 12219 2975
rect 12161 2935 12219 2941
rect 12894 2932 12900 2984
rect 12952 2972 12958 2984
rect 13173 2975 13231 2981
rect 13173 2972 13185 2975
rect 12952 2944 13185 2972
rect 12952 2932 12958 2944
rect 13173 2941 13185 2944
rect 13219 2941 13231 2975
rect 13173 2935 13231 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15712 2944 16037 2972
rect 15712 2932 15718 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16025 2935 16083 2941
rect 9272 2876 10824 2904
rect 11149 2907 11207 2913
rect 9272 2864 9278 2876
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 13906 2904 13912 2916
rect 11195 2876 13912 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 17144 2904 17172 3003
rect 18966 3000 18972 3052
rect 19024 3000 19030 3052
rect 19076 3012 20760 3040
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 17494 2972 17500 2984
rect 17451 2944 17500 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 18414 2972 18420 2984
rect 18371 2944 18420 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 19076 2972 19104 3012
rect 18984 2944 19104 2972
rect 20732 2972 20760 3012
rect 20806 3000 20812 3052
rect 20864 3000 20870 3052
rect 20898 3000 20904 3052
rect 20956 3000 20962 3052
rect 20990 3000 20996 3052
rect 21048 3040 21054 3052
rect 21085 3043 21143 3049
rect 21085 3040 21097 3043
rect 21048 3012 21097 3040
rect 21048 3000 21054 3012
rect 21085 3009 21097 3012
rect 21131 3009 21143 3043
rect 21085 3003 21143 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3009 21235 3043
rect 21177 3003 21235 3009
rect 21315 3043 21373 3049
rect 21315 3009 21327 3043
rect 21361 3040 21373 3043
rect 22186 3040 22192 3052
rect 21361 3012 22192 3040
rect 21361 3009 21373 3012
rect 21315 3003 21373 3009
rect 20916 2972 20944 3000
rect 20732 2944 20944 2972
rect 18984 2904 19012 2944
rect 17144 2876 19012 2904
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 9766 2836 9772 2848
rect 9355 2808 9772 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 12529 2839 12587 2845
rect 12529 2805 12541 2839
rect 12575 2836 12587 2839
rect 15194 2836 15200 2848
rect 12575 2808 15200 2836
rect 12575 2805 12587 2808
rect 12529 2799 12587 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15286 2796 15292 2848
rect 15344 2796 15350 2848
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 20349 2839 20407 2845
rect 20349 2836 20361 2839
rect 18012 2808 20361 2836
rect 18012 2796 18018 2808
rect 20349 2805 20361 2808
rect 20395 2836 20407 2839
rect 20530 2836 20536 2848
rect 20395 2808 20536 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 21192 2836 21220 3003
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22572 3049 22600 3080
rect 25866 3068 25872 3080
rect 25924 3068 25930 3120
rect 28077 3111 28135 3117
rect 28077 3077 28089 3111
rect 28123 3108 28135 3111
rect 29012 3108 29040 3136
rect 31297 3111 31355 3117
rect 31297 3108 31309 3111
rect 28123 3080 29040 3108
rect 30116 3080 31309 3108
rect 28123 3077 28135 3080
rect 28077 3071 28135 3077
rect 22557 3043 22615 3049
rect 22557 3009 22569 3043
rect 22603 3009 22615 3043
rect 22557 3003 22615 3009
rect 22824 3043 22882 3049
rect 22824 3009 22836 3043
rect 22870 3040 22882 3043
rect 23566 3040 23572 3052
rect 22870 3012 23572 3040
rect 22870 3009 22882 3012
rect 22824 3003 22882 3009
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 24946 3000 24952 3052
rect 25004 3000 25010 3052
rect 27341 3043 27399 3049
rect 27341 3009 27353 3043
rect 27387 3040 27399 3043
rect 27522 3040 27528 3052
rect 27387 3012 27528 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 27522 3000 27528 3012
rect 27580 3000 27586 3052
rect 28988 3043 29046 3049
rect 28988 3009 29000 3043
rect 29034 3040 29046 3043
rect 30116 3040 30144 3080
rect 31297 3077 31309 3080
rect 31343 3077 31355 3111
rect 31297 3071 31355 3077
rect 32582 3068 32588 3120
rect 32640 3068 32646 3120
rect 33413 3111 33471 3117
rect 33413 3077 33425 3111
rect 33459 3108 33471 3111
rect 33502 3108 33508 3120
rect 33459 3080 33508 3108
rect 33459 3077 33471 3080
rect 33413 3071 33471 3077
rect 33502 3068 33508 3080
rect 33560 3068 33566 3120
rect 35894 3068 35900 3120
rect 35952 3108 35958 3120
rect 37553 3111 37611 3117
rect 37553 3108 37565 3111
rect 35952 3080 37565 3108
rect 35952 3068 35958 3080
rect 37553 3077 37565 3080
rect 37599 3077 37611 3111
rect 41046 3108 41052 3120
rect 37553 3071 37611 3077
rect 38212 3080 41052 3108
rect 38212 3052 38240 3080
rect 29034 3012 30144 3040
rect 29034 3009 29046 3012
rect 28988 3003 29046 3009
rect 30558 3000 30564 3052
rect 30616 3000 30622 3052
rect 30742 2998 30748 3050
rect 30800 2998 30806 3050
rect 30929 3043 30987 3049
rect 30929 3009 30941 3043
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 31113 3043 31171 3049
rect 31113 3009 31125 3043
rect 31159 3040 31171 3043
rect 31202 3040 31208 3052
rect 31159 3012 31208 3040
rect 31159 3009 31171 3012
rect 31113 3003 31171 3009
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 25133 2975 25191 2981
rect 25133 2972 25145 2975
rect 24912 2944 25145 2972
rect 24912 2932 24918 2944
rect 25133 2941 25145 2944
rect 25179 2941 25191 2975
rect 25133 2935 25191 2941
rect 25866 2932 25872 2984
rect 25924 2972 25930 2984
rect 28721 2975 28779 2981
rect 28721 2972 28733 2975
rect 25924 2944 28733 2972
rect 25924 2932 25930 2944
rect 28721 2941 28733 2944
rect 28767 2941 28779 2975
rect 28721 2935 28779 2941
rect 30831 2975 30889 2981
rect 30831 2941 30843 2975
rect 30877 2941 30889 2975
rect 30944 2972 30972 3003
rect 31202 3000 31208 3012
rect 31260 3000 31266 3052
rect 31754 3000 31760 3052
rect 31812 3040 31818 3052
rect 32401 3043 32459 3049
rect 32401 3040 32413 3043
rect 31812 3012 32413 3040
rect 31812 3000 31818 3012
rect 32401 3009 32413 3012
rect 32447 3009 32459 3043
rect 32401 3003 32459 3009
rect 33134 3000 33140 3052
rect 33192 3040 33198 3052
rect 33229 3043 33287 3049
rect 33229 3040 33241 3043
rect 33192 3012 33241 3040
rect 33192 3000 33198 3012
rect 33229 3009 33241 3012
rect 33275 3009 33287 3043
rect 33229 3003 33287 3009
rect 33870 3000 33876 3052
rect 33928 3000 33934 3052
rect 33962 3000 33968 3052
rect 34020 3040 34026 3052
rect 34129 3043 34187 3049
rect 34129 3040 34141 3043
rect 34020 3012 34141 3040
rect 34020 3000 34026 3012
rect 34129 3009 34141 3012
rect 34175 3009 34187 3043
rect 34129 3003 34187 3009
rect 36446 3000 36452 3052
rect 36504 3000 36510 3052
rect 38194 3000 38200 3052
rect 38252 3000 38258 3052
rect 38286 3000 38292 3052
rect 38344 3040 38350 3052
rect 40604 3049 40632 3080
rect 41046 3068 41052 3080
rect 41104 3068 41110 3120
rect 41506 3068 41512 3120
rect 41564 3108 41570 3120
rect 42705 3111 42763 3117
rect 42705 3108 42717 3111
rect 41564 3080 42717 3108
rect 41564 3068 41570 3080
rect 42705 3077 42717 3080
rect 42751 3077 42763 3111
rect 42705 3071 42763 3077
rect 45278 3068 45284 3120
rect 45336 3108 45342 3120
rect 45336 3080 48912 3108
rect 45336 3068 45342 3080
rect 38453 3043 38511 3049
rect 38453 3040 38465 3043
rect 38344 3012 38465 3040
rect 38344 3000 38350 3012
rect 38453 3009 38465 3012
rect 38499 3009 38511 3043
rect 38453 3003 38511 3009
rect 40589 3043 40647 3049
rect 40589 3009 40601 3043
rect 40635 3009 40647 3043
rect 40589 3003 40647 3009
rect 40856 3043 40914 3049
rect 40856 3009 40868 3043
rect 40902 3040 40914 3043
rect 41414 3040 41420 3052
rect 40902 3012 41420 3040
rect 40902 3009 40914 3012
rect 40856 3003 40914 3009
rect 41414 3000 41420 3012
rect 41472 3000 41478 3052
rect 42794 3000 42800 3052
rect 42852 3040 42858 3052
rect 43441 3043 43499 3049
rect 43441 3040 43453 3043
rect 42852 3012 43453 3040
rect 42852 3000 42858 3012
rect 43441 3009 43453 3012
rect 43487 3009 43499 3043
rect 43441 3003 43499 3009
rect 44174 3000 44180 3052
rect 44232 3040 44238 3052
rect 44361 3043 44419 3049
rect 44361 3040 44373 3043
rect 44232 3012 44373 3040
rect 44232 3000 44238 3012
rect 44361 3009 44373 3012
rect 44407 3009 44419 3043
rect 44361 3003 44419 3009
rect 45554 3000 45560 3052
rect 45612 3040 45618 3052
rect 45741 3043 45799 3049
rect 45741 3040 45753 3043
rect 45612 3012 45753 3040
rect 45612 3000 45618 3012
rect 45741 3009 45753 3012
rect 45787 3009 45799 3043
rect 45741 3003 45799 3009
rect 46934 3000 46940 3052
rect 46992 3040 46998 3052
rect 48884 3049 48912 3080
rect 56962 3068 56968 3120
rect 57020 3068 57026 3120
rect 47857 3043 47915 3049
rect 47857 3040 47869 3043
rect 46992 3012 47869 3040
rect 46992 3000 46998 3012
rect 47857 3009 47869 3012
rect 47903 3009 47915 3043
rect 47857 3003 47915 3009
rect 48869 3043 48927 3049
rect 48869 3009 48881 3043
rect 48915 3009 48927 3043
rect 48869 3003 48927 3009
rect 49694 3000 49700 3052
rect 49752 3040 49758 3052
rect 50249 3043 50307 3049
rect 50249 3040 50261 3043
rect 49752 3012 50261 3040
rect 49752 3000 49758 3012
rect 50249 3009 50261 3012
rect 50295 3009 50307 3043
rect 50249 3003 50307 3009
rect 51626 3000 51632 3052
rect 51684 3000 51690 3052
rect 53834 3000 53840 3052
rect 53892 3040 53898 3052
rect 54021 3043 54079 3049
rect 54021 3040 54033 3043
rect 53892 3012 54033 3040
rect 53892 3000 53898 3012
rect 54021 3009 54033 3012
rect 54067 3009 54079 3043
rect 54021 3003 54079 3009
rect 54846 3000 54852 3052
rect 54904 3000 54910 3052
rect 55861 3043 55919 3049
rect 55861 3009 55873 3043
rect 55907 3009 55919 3043
rect 55861 3003 55919 3009
rect 31478 2972 31484 2984
rect 30944 2944 31484 2972
rect 30831 2935 30889 2941
rect 23492 2876 24992 2904
rect 23492 2836 23520 2876
rect 24964 2848 24992 2876
rect 30742 2864 30748 2916
rect 30800 2904 30806 2916
rect 30852 2904 30880 2935
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 36354 2932 36360 2984
rect 36412 2972 36418 2984
rect 36633 2975 36691 2981
rect 36633 2972 36645 2975
rect 36412 2944 36645 2972
rect 36412 2932 36418 2944
rect 36633 2941 36645 2944
rect 36679 2941 36691 2975
rect 36633 2935 36691 2941
rect 48774 2932 48780 2984
rect 48832 2972 48838 2984
rect 49053 2975 49111 2981
rect 49053 2972 49065 2975
rect 48832 2944 49065 2972
rect 48832 2932 48838 2944
rect 49053 2941 49065 2944
rect 49099 2941 49111 2975
rect 49053 2935 49111 2941
rect 50154 2932 50160 2984
rect 50212 2972 50218 2984
rect 50433 2975 50491 2981
rect 50433 2972 50445 2975
rect 50212 2944 50445 2972
rect 50212 2932 50218 2944
rect 50433 2941 50445 2944
rect 50479 2941 50491 2975
rect 50433 2935 50491 2941
rect 51534 2932 51540 2984
rect 51592 2972 51598 2984
rect 51813 2975 51871 2981
rect 51813 2972 51825 2975
rect 51592 2944 51825 2972
rect 51592 2932 51598 2944
rect 51813 2941 51825 2944
rect 51859 2941 51871 2975
rect 51813 2935 51871 2941
rect 54294 2932 54300 2984
rect 54352 2972 54358 2984
rect 55033 2975 55091 2981
rect 55033 2972 55045 2975
rect 54352 2944 55045 2972
rect 54352 2932 54358 2944
rect 55033 2941 55045 2944
rect 55079 2941 55091 2975
rect 55876 2972 55904 3003
rect 56594 3000 56600 3052
rect 56652 3040 56658 3052
rect 56689 3043 56747 3049
rect 56689 3040 56701 3043
rect 56652 3012 56701 3040
rect 56652 3000 56658 3012
rect 56689 3009 56701 3012
rect 56735 3009 56747 3043
rect 56689 3003 56747 3009
rect 57974 2972 57980 2984
rect 55876 2944 57980 2972
rect 55033 2935 55091 2941
rect 57974 2932 57980 2944
rect 58032 2932 58038 2984
rect 30800 2876 30880 2904
rect 41969 2907 42027 2913
rect 30800 2864 30806 2876
rect 41969 2873 41981 2907
rect 42015 2904 42027 2907
rect 44358 2904 44364 2916
rect 42015 2876 44364 2904
rect 42015 2873 42027 2876
rect 41969 2867 42027 2873
rect 21192 2808 23520 2836
rect 24946 2796 24952 2848
rect 25004 2796 25010 2848
rect 40218 2796 40224 2848
rect 40276 2836 40282 2848
rect 41984 2836 42012 2867
rect 44358 2864 44364 2876
rect 44416 2864 44422 2916
rect 40276 2808 42012 2836
rect 40276 2796 40282 2808
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 32306 2632 32312 2644
rect 7944 2604 21956 2632
rect 5442 2496 5448 2508
rect 4264 2468 5448 2496
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 4264 2437 4292 2468
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 5166 2388 5172 2440
rect 5224 2388 5230 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7098 2428 7104 2440
rect 7055 2400 7104 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7944 2437 7972 2604
rect 15286 2564 15292 2576
rect 12360 2536 15292 2564
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 12360 2437 12388 2536
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 21818 2564 21824 2576
rect 18432 2536 21824 2564
rect 13648 2468 18368 2496
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 12345 2431 12403 2437
rect 10735 2400 12296 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 2317 2363 2375 2369
rect 2317 2329 2329 2363
rect 2363 2360 2375 2363
rect 2774 2360 2780 2372
rect 2363 2332 2780 2360
rect 2363 2329 2375 2332
rect 2317 2323 2375 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 4062 2360 4068 2372
rect 3283 2332 4068 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 4614 2360 4620 2372
rect 4571 2332 4620 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 5445 2363 5503 2369
rect 5445 2360 5457 2363
rect 5132 2332 5457 2360
rect 5132 2320 5138 2332
rect 5445 2329 5457 2332
rect 5491 2329 5503 2363
rect 5445 2323 5503 2329
rect 7285 2363 7343 2369
rect 7285 2329 7297 2363
rect 7331 2360 7343 2363
rect 7374 2360 7380 2372
rect 7331 2332 7380 2360
rect 7331 2329 7343 2332
rect 7285 2323 7343 2329
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 7834 2320 7840 2372
rect 7892 2360 7898 2372
rect 8205 2363 8263 2369
rect 8205 2360 8217 2363
rect 7892 2332 8217 2360
rect 7892 2320 7898 2332
rect 8205 2329 8217 2332
rect 8251 2329 8263 2363
rect 8205 2323 8263 2329
rect 10045 2363 10103 2369
rect 10045 2329 10057 2363
rect 10091 2360 10103 2363
rect 10134 2360 10140 2372
rect 10091 2332 10140 2360
rect 10091 2329 10103 2332
rect 10045 2323 10103 2329
rect 10134 2320 10140 2332
rect 10192 2320 10198 2372
rect 10594 2320 10600 2372
rect 10652 2360 10658 2372
rect 10965 2363 11023 2369
rect 10965 2360 10977 2363
rect 10652 2332 10977 2360
rect 10652 2320 10658 2332
rect 10965 2329 10977 2332
rect 11011 2329 11023 2363
rect 10965 2323 11023 2329
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 8570 2292 8576 2304
rect 3476 2264 8576 2292
rect 3476 2252 3482 2264
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 9214 2292 9220 2304
rect 9171 2264 9220 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 11974 2292 11980 2304
rect 11747 2264 11980 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 12268 2292 12296 2400
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 12492 2332 12633 2360
rect 12492 2320 12498 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 13354 2320 13360 2372
rect 13412 2360 13418 2372
rect 13541 2363 13599 2369
rect 13541 2360 13553 2363
rect 13412 2332 13553 2360
rect 13412 2320 13418 2332
rect 13541 2329 13553 2332
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 13648 2292 13676 2468
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15838 2388 15844 2440
rect 15896 2388 15902 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 15194 2320 15200 2372
rect 15252 2320 15258 2372
rect 16114 2320 16120 2372
rect 16172 2320 16178 2372
rect 17773 2363 17831 2369
rect 17773 2329 17785 2363
rect 17819 2360 17831 2363
rect 17862 2360 17868 2372
rect 17819 2332 17868 2360
rect 17819 2329 17831 2332
rect 17773 2323 17831 2329
rect 17862 2320 17868 2332
rect 17920 2320 17926 2372
rect 18340 2360 18368 2468
rect 18432 2437 18460 2536
rect 21818 2524 21824 2536
rect 21876 2524 21882 2576
rect 21928 2564 21956 2604
rect 25424 2604 32312 2632
rect 24762 2564 24768 2576
rect 21928 2536 24768 2564
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 24857 2567 24915 2573
rect 24857 2533 24869 2567
rect 24903 2564 24915 2567
rect 24946 2564 24952 2576
rect 24903 2536 24952 2564
rect 24903 2533 24915 2536
rect 24857 2527 24915 2533
rect 24946 2524 24952 2536
rect 25004 2524 25010 2576
rect 22462 2496 22468 2508
rect 18524 2468 22468 2496
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 18524 2360 18552 2468
rect 22462 2456 22468 2468
rect 22520 2456 22526 2508
rect 25130 2496 25136 2508
rect 22664 2468 25136 2496
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2428 21051 2431
rect 22094 2428 22100 2440
rect 21039 2400 22100 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 18340 2332 18552 2360
rect 18690 2320 18696 2372
rect 18748 2320 18754 2372
rect 12268 2264 13676 2292
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 14734 2292 14740 2304
rect 14323 2264 14740 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 20088 2292 20116 2391
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 22664 2437 22692 2468
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 20349 2363 20407 2369
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 20622 2360 20628 2372
rect 20395 2332 20628 2360
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 22002 2360 22008 2372
rect 21315 2332 22008 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 22002 2320 22008 2332
rect 22060 2320 22066 2372
rect 22925 2363 22983 2369
rect 22925 2329 22937 2363
rect 22971 2360 22983 2363
rect 23014 2360 23020 2372
rect 22971 2332 23020 2360
rect 22971 2329 22983 2332
rect 22925 2323 22983 2329
rect 23014 2320 23020 2332
rect 23072 2320 23078 2372
rect 23474 2292 23480 2304
rect 20088 2264 23480 2292
rect 23474 2252 23480 2264
rect 23532 2252 23538 2304
rect 23584 2292 23612 2391
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 25424 2437 25452 2604
rect 32306 2592 32312 2604
rect 32364 2592 32370 2644
rect 33502 2592 33508 2644
rect 33560 2632 33566 2644
rect 34238 2632 34244 2644
rect 33560 2604 34244 2632
rect 33560 2592 33566 2604
rect 34238 2592 34244 2604
rect 34296 2592 34302 2644
rect 35526 2592 35532 2644
rect 35584 2592 35590 2644
rect 36906 2592 36912 2644
rect 36964 2632 36970 2644
rect 38933 2635 38991 2641
rect 38933 2632 38945 2635
rect 36964 2604 38945 2632
rect 36964 2592 36970 2604
rect 38933 2601 38945 2604
rect 38979 2601 38991 2635
rect 38933 2595 38991 2601
rect 40310 2592 40316 2644
rect 40368 2632 40374 2644
rect 40368 2604 49740 2632
rect 40368 2592 40374 2604
rect 26605 2567 26663 2573
rect 26605 2533 26617 2567
rect 26651 2564 26663 2567
rect 27430 2564 27436 2576
rect 26651 2536 27436 2564
rect 26651 2533 26663 2536
rect 26605 2527 26663 2533
rect 27430 2524 27436 2536
rect 27488 2524 27494 2576
rect 30190 2524 30196 2576
rect 30248 2564 30254 2576
rect 49712 2564 49740 2604
rect 53098 2592 53104 2644
rect 53156 2592 53162 2644
rect 30248 2536 46980 2564
rect 49712 2536 53880 2564
rect 30248 2524 30254 2536
rect 33502 2496 33508 2508
rect 31956 2468 33508 2496
rect 24673 2431 24731 2437
rect 24673 2428 24685 2431
rect 23992 2400 24685 2428
rect 23992 2388 23998 2400
rect 24673 2397 24685 2400
rect 24719 2397 24731 2431
rect 24673 2391 24731 2397
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 27157 2431 27215 2437
rect 27157 2397 27169 2431
rect 27203 2428 27215 2431
rect 28169 2431 28227 2437
rect 27203 2400 28028 2428
rect 27203 2397 27215 2400
rect 27157 2391 27215 2397
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24394 2360 24400 2372
rect 23891 2332 24400 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24394 2320 24400 2332
rect 24452 2320 24458 2372
rect 25314 2320 25320 2372
rect 25372 2360 25378 2372
rect 25685 2363 25743 2369
rect 25685 2360 25697 2363
rect 25372 2332 25697 2360
rect 25372 2320 25378 2332
rect 25685 2329 25697 2332
rect 25731 2329 25743 2363
rect 25685 2323 25743 2329
rect 26234 2320 26240 2372
rect 26292 2360 26298 2372
rect 26421 2363 26479 2369
rect 26421 2360 26433 2363
rect 26292 2332 26433 2360
rect 26292 2320 26298 2332
rect 26421 2329 26433 2332
rect 26467 2329 26479 2363
rect 26421 2323 26479 2329
rect 26694 2320 26700 2372
rect 26752 2360 26758 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 26752 2332 27445 2360
rect 26752 2320 26758 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 26326 2292 26332 2304
rect 23584 2264 26332 2292
rect 26326 2252 26332 2264
rect 26384 2252 26390 2304
rect 28000 2292 28028 2400
rect 28169 2397 28181 2431
rect 28215 2428 28227 2431
rect 28258 2428 28264 2440
rect 28215 2400 28264 2428
rect 28215 2397 28227 2400
rect 28169 2391 28227 2397
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30926 2388 30932 2440
rect 30984 2388 30990 2440
rect 28074 2320 28080 2372
rect 28132 2360 28138 2372
rect 28445 2363 28503 2369
rect 28445 2360 28457 2363
rect 28132 2332 28457 2360
rect 28132 2320 28138 2332
rect 28445 2329 28457 2332
rect 28491 2329 28503 2363
rect 28445 2323 28503 2329
rect 29454 2320 29460 2372
rect 29512 2360 29518 2372
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 29512 2332 30021 2360
rect 29512 2320 29518 2332
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 30009 2323 30067 2329
rect 30834 2320 30840 2372
rect 30892 2360 30898 2372
rect 31205 2363 31263 2369
rect 31205 2360 31217 2363
rect 30892 2332 31217 2360
rect 30892 2320 30898 2332
rect 31205 2329 31217 2332
rect 31251 2329 31263 2363
rect 31205 2323 31263 2329
rect 31956 2292 31984 2468
rect 33502 2456 33508 2468
rect 33560 2456 33566 2508
rect 33594 2456 33600 2508
rect 33652 2456 33658 2508
rect 37274 2496 37280 2508
rect 35268 2468 37280 2496
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2428 32367 2431
rect 33612 2428 33640 2456
rect 35268 2440 35296 2468
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 42426 2456 42432 2508
rect 42484 2496 42490 2508
rect 42484 2468 43668 2496
rect 42484 2456 42490 2468
rect 32355 2400 33640 2428
rect 32355 2397 32367 2400
rect 32309 2391 32367 2397
rect 33686 2388 33692 2440
rect 33744 2388 33750 2440
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34664 2400 34897 2428
rect 34664 2388 34670 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35032 2400 35077 2428
rect 35032 2388 35038 2400
rect 35250 2388 35256 2440
rect 35308 2388 35314 2440
rect 35350 2431 35408 2437
rect 35350 2397 35362 2431
rect 35396 2397 35408 2431
rect 35350 2391 35408 2397
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 32585 2363 32643 2369
rect 32585 2360 32597 2363
rect 32272 2332 32597 2360
rect 32272 2320 32278 2332
rect 32585 2329 32597 2332
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 33594 2320 33600 2372
rect 33652 2360 33658 2372
rect 33965 2363 34023 2369
rect 33965 2360 33977 2363
rect 33652 2332 33977 2360
rect 33652 2320 33658 2332
rect 33965 2329 33977 2332
rect 34011 2329 34023 2363
rect 33965 2323 34023 2329
rect 34054 2320 34060 2372
rect 34112 2360 34118 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 34112 2332 35173 2360
rect 34112 2320 34118 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 28000 2264 31984 2292
rect 32030 2252 32036 2304
rect 32088 2292 32094 2304
rect 35360 2292 35388 2391
rect 35618 2388 35624 2440
rect 35676 2428 35682 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35676 2400 36001 2428
rect 35676 2388 35682 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 37826 2388 37832 2440
rect 37884 2388 37890 2440
rect 39206 2388 39212 2440
rect 39264 2428 39270 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39264 2400 40049 2428
rect 39264 2388 39270 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 40954 2388 40960 2440
rect 41012 2388 41018 2440
rect 42518 2388 42524 2440
rect 42576 2428 42582 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 42576 2400 42625 2428
rect 42576 2388 42582 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 43438 2388 43444 2440
rect 43496 2428 43502 2440
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 43496 2400 43545 2428
rect 43496 2388 43502 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43640 2428 43668 2468
rect 43806 2456 43812 2508
rect 43864 2496 43870 2508
rect 46952 2496 46980 2536
rect 50709 2499 50767 2505
rect 50709 2496 50721 2499
rect 43864 2468 45554 2496
rect 46952 2468 50721 2496
rect 43864 2456 43870 2468
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 43640 2400 45201 2428
rect 43533 2391 43591 2397
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 45526 2428 45554 2468
rect 50709 2465 50721 2468
rect 50755 2465 50767 2499
rect 50709 2459 50767 2465
rect 53852 2437 53880 2536
rect 46109 2431 46167 2437
rect 46109 2428 46121 2431
rect 45526 2400 46121 2428
rect 45189 2391 45247 2397
rect 46109 2397 46121 2400
rect 46155 2397 46167 2431
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46109 2391 46167 2397
rect 46676 2400 47777 2428
rect 36262 2320 36268 2372
rect 36320 2320 36326 2372
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 38105 2363 38163 2369
rect 38105 2360 38117 2363
rect 37792 2332 38117 2360
rect 37792 2320 37798 2332
rect 38105 2329 38117 2332
rect 38151 2329 38163 2363
rect 38105 2323 38163 2329
rect 38838 2320 38844 2372
rect 38896 2320 38902 2372
rect 40310 2320 40316 2372
rect 40368 2320 40374 2372
rect 40494 2320 40500 2372
rect 40552 2360 40558 2372
rect 41233 2363 41291 2369
rect 41233 2360 41245 2363
rect 40552 2332 41245 2360
rect 40552 2320 40558 2332
rect 41233 2329 41245 2332
rect 41279 2329 41291 2363
rect 41233 2323 41291 2329
rect 42886 2320 42892 2372
rect 42944 2320 42950 2372
rect 43254 2320 43260 2372
rect 43312 2360 43318 2372
rect 43809 2363 43867 2369
rect 43809 2360 43821 2363
rect 43312 2332 43821 2360
rect 43312 2320 43318 2332
rect 43809 2329 43821 2332
rect 43855 2329 43867 2363
rect 43809 2323 43867 2329
rect 44634 2320 44640 2372
rect 44692 2360 44698 2372
rect 45465 2363 45523 2369
rect 45465 2360 45477 2363
rect 44692 2332 45477 2360
rect 44692 2320 44698 2332
rect 45465 2329 45477 2332
rect 45511 2329 45523 2363
rect 45465 2323 45523 2329
rect 46014 2320 46020 2372
rect 46072 2360 46078 2372
rect 46385 2363 46443 2369
rect 46385 2360 46397 2363
rect 46072 2332 46397 2360
rect 46072 2320 46078 2332
rect 46385 2329 46397 2332
rect 46431 2329 46443 2363
rect 46385 2323 46443 2329
rect 32088 2264 35388 2292
rect 32088 2252 32094 2264
rect 44266 2252 44272 2304
rect 44324 2292 44330 2304
rect 46676 2292 46704 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 53837 2431 53895 2437
rect 53837 2397 53849 2431
rect 53883 2397 53895 2431
rect 53837 2391 53895 2397
rect 55214 2388 55220 2440
rect 55272 2428 55278 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55272 2400 55505 2428
rect 55272 2388 55278 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 56410 2388 56416 2440
rect 56468 2388 56474 2440
rect 47394 2320 47400 2372
rect 47452 2360 47458 2372
rect 48041 2363 48099 2369
rect 48041 2360 48053 2363
rect 47452 2332 48053 2360
rect 47452 2320 47458 2332
rect 48041 2329 48053 2332
rect 48087 2329 48099 2363
rect 48041 2323 48099 2329
rect 48314 2320 48320 2372
rect 48372 2360 48378 2372
rect 48777 2363 48835 2369
rect 48777 2360 48789 2363
rect 48372 2332 48789 2360
rect 48372 2320 48378 2332
rect 48777 2329 48789 2332
rect 48823 2329 48835 2363
rect 48777 2323 48835 2329
rect 49694 2320 49700 2372
rect 49752 2360 49758 2372
rect 50433 2363 50491 2369
rect 50433 2360 50445 2363
rect 49752 2332 50445 2360
rect 49752 2320 49758 2332
rect 50433 2329 50445 2332
rect 50479 2329 50491 2363
rect 50433 2323 50491 2329
rect 51074 2320 51080 2372
rect 51132 2360 51138 2372
rect 51353 2363 51411 2369
rect 51353 2360 51365 2363
rect 51132 2332 51365 2360
rect 51132 2320 51138 2332
rect 51353 2329 51365 2332
rect 51399 2329 51411 2363
rect 51353 2323 51411 2329
rect 52454 2320 52460 2372
rect 52512 2360 52518 2372
rect 53009 2363 53067 2369
rect 53009 2360 53021 2363
rect 52512 2332 53021 2360
rect 52512 2320 52518 2332
rect 53009 2329 53021 2332
rect 53055 2329 53067 2363
rect 53009 2323 53067 2329
rect 54110 2320 54116 2372
rect 54168 2320 54174 2372
rect 55766 2320 55772 2372
rect 55824 2320 55830 2372
rect 56686 2320 56692 2372
rect 56744 2320 56750 2372
rect 44324 2264 46704 2292
rect 44324 2252 44330 2264
rect 48866 2252 48872 2304
rect 48924 2252 48930 2304
rect 51442 2252 51448 2304
rect 51500 2252 51506 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 22462 2048 22468 2100
rect 22520 2088 22526 2100
rect 30466 2088 30472 2100
rect 22520 2060 30472 2088
rect 22520 2048 22526 2060
rect 30466 2048 30472 2060
rect 30524 2048 30530 2100
rect 2866 1980 2872 2032
rect 2924 2020 2930 2032
rect 4798 2020 4804 2032
rect 2924 1992 4804 2020
rect 2924 1980 2930 1992
rect 4798 1980 4804 1992
rect 4856 1980 4862 2032
rect 5166 1980 5172 2032
rect 5224 2020 5230 2032
rect 11330 2020 11336 2032
rect 5224 1992 11336 2020
rect 5224 1980 5230 1992
rect 11330 1980 11336 1992
rect 11388 1980 11394 2032
rect 12986 1980 12992 2032
rect 13044 2020 13050 2032
rect 48866 2020 48872 2032
rect 13044 1992 48872 2020
rect 13044 1980 13050 1992
rect 48866 1980 48872 1992
rect 48924 1980 48930 2032
rect 2958 1912 2964 1964
rect 3016 1952 3022 1964
rect 11146 1952 11152 1964
rect 3016 1924 11152 1952
rect 3016 1912 3022 1924
rect 11146 1912 11152 1924
rect 11204 1912 11210 1964
rect 15838 1912 15844 1964
rect 15896 1952 15902 1964
rect 15896 1924 22094 1952
rect 15896 1912 15902 1924
rect 2038 1844 2044 1896
rect 2096 1884 2102 1896
rect 11698 1884 11704 1896
rect 2096 1856 11704 1884
rect 2096 1844 2102 1856
rect 11698 1844 11704 1856
rect 11756 1844 11762 1896
rect 22066 1884 22094 1924
rect 23474 1912 23480 1964
rect 23532 1952 23538 1964
rect 27154 1952 27160 1964
rect 23532 1924 27160 1952
rect 23532 1912 23538 1924
rect 27154 1912 27160 1924
rect 27212 1912 27218 1964
rect 46842 1912 46848 1964
rect 46900 1952 46906 1964
rect 56410 1952 56416 1964
rect 46900 1924 56416 1952
rect 46900 1912 46906 1924
rect 56410 1912 56416 1924
rect 56468 1912 56474 1964
rect 30742 1884 30748 1896
rect 22066 1856 30748 1884
rect 30742 1844 30748 1856
rect 30800 1884 30806 1896
rect 35250 1884 35256 1896
rect 30800 1856 35256 1884
rect 30800 1844 30806 1856
rect 35250 1844 35256 1856
rect 35308 1844 35314 1896
rect 6086 1776 6092 1828
rect 6144 1816 6150 1828
rect 51442 1816 51448 1828
rect 6144 1788 51448 1816
rect 6144 1776 6150 1788
rect 51442 1776 51448 1788
rect 51500 1776 51506 1828
rect 13262 1708 13268 1760
rect 13320 1748 13326 1760
rect 31386 1748 31392 1760
rect 13320 1720 31392 1748
rect 13320 1708 13326 1720
rect 31386 1708 31392 1720
rect 31444 1708 31450 1760
rect 8846 1640 8852 1692
rect 8904 1680 8910 1692
rect 55766 1680 55772 1692
rect 8904 1652 55772 1680
rect 8904 1640 8910 1652
rect 55766 1640 55772 1652
rect 55824 1640 55830 1692
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 21910 1340 21916 1352
rect 3384 1312 21916 1340
rect 3384 1300 3390 1312
rect 21910 1300 21916 1312
rect 21968 1300 21974 1352
rect 18690 892 18696 944
rect 18748 932 18754 944
rect 19794 932 19800 944
rect 18748 904 19800 932
rect 18748 892 18754 904
rect 19794 892 19800 904
rect 19852 892 19858 944
rect 34974 892 34980 944
rect 35032 932 35038 944
rect 36262 932 36268 944
rect 35032 904 36268 932
rect 35032 892 35038 904
rect 36262 892 36268 904
rect 36320 892 36326 944
rect 37274 892 37280 944
rect 37332 932 37338 944
rect 38838 932 38844 944
rect 37332 904 38844 932
rect 37332 892 37338 904
rect 38838 892 38844 904
rect 38896 892 38902 944
rect 39114 892 39120 944
rect 39172 932 39178 944
rect 40310 932 40316 944
rect 39172 904 40316 932
rect 39172 892 39178 904
rect 40310 892 40316 904
rect 40368 892 40374 944
rect 41874 892 41880 944
rect 41932 932 41938 944
rect 42886 932 42892 944
rect 41932 904 42892 932
rect 41932 892 41938 904
rect 42886 892 42892 904
rect 42944 892 42950 944
rect 52914 892 52920 944
rect 52972 932 52978 944
rect 54110 932 54116 944
rect 52972 904 54116 932
rect 52972 892 52978 904
rect 54110 892 54116 904
rect 54168 892 54174 944
rect 55674 892 55680 944
rect 55732 932 55738 944
rect 56686 932 56692 944
rect 55732 904 56692 932
rect 55732 892 55738 904
rect 56686 892 56692 904
rect 56744 892 56750 944
<< via1 >>
rect 3884 41080 3936 41132
rect 4620 41080 4672 41132
rect 18788 41080 18840 41132
rect 19432 41080 19484 41132
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 41420 39627 41472 39636
rect 41420 39593 41429 39627
rect 41429 39593 41463 39627
rect 41463 39593 41472 39627
rect 41420 39584 41472 39593
rect 48596 39584 48648 39636
rect 940 39448 992 39500
rect 3424 39448 3476 39500
rect 4620 39448 4672 39500
rect 19432 39491 19484 39500
rect 19432 39457 19441 39491
rect 19441 39457 19475 39491
rect 19475 39457 19484 39491
rect 19432 39448 19484 39457
rect 26240 39448 26292 39500
rect 56048 39448 56100 39500
rect 2504 39423 2556 39432
rect 2504 39389 2513 39423
rect 2513 39389 2547 39423
rect 2547 39389 2556 39423
rect 2504 39380 2556 39389
rect 1032 39312 1084 39364
rect 27160 39423 27212 39432
rect 27160 39389 27169 39423
rect 27169 39389 27203 39423
rect 27203 39389 27212 39423
rect 27160 39380 27212 39389
rect 33692 39380 33744 39432
rect 42156 39380 42208 39432
rect 28264 39312 28316 39364
rect 33324 39244 33376 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 7656 38972 7708 39024
rect 6184 38904 6236 38956
rect 940 38836 992 38888
rect 1124 38768 1176 38820
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 10324 38292 10376 38344
rect 940 38224 992 38276
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 6184 37884 6236 37936
rect 14280 37884 14332 37936
rect 2504 37612 2556 37664
rect 6000 37612 6052 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 3424 37408 3476 37460
rect 5356 37408 5408 37460
rect 4068 37204 4120 37256
rect 940 37136 992 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 11980 36728 12032 36780
rect 940 36660 992 36712
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 11704 35640 11756 35692
rect 940 35572 992 35624
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5540 35028 5592 35080
rect 940 34960 992 35012
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4620 34620 4672 34672
rect 1032 34552 1084 34604
rect 940 34484 992 34536
rect 2688 34484 2740 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1124 33872 1176 33924
rect 2136 33872 2188 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 23756 33464 23808 33516
rect 940 33396 992 33448
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 940 32784 992 32836
rect 2504 32784 2556 32836
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 5540 32444 5592 32496
rect 22836 32444 22888 32496
rect 12440 32376 12492 32428
rect 940 32308 992 32360
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1032 31832 1084 31884
rect 4068 31900 4120 31952
rect 6184 31900 6236 31952
rect 940 31764 992 31816
rect 6644 31832 6696 31884
rect 2596 31807 2648 31816
rect 2596 31773 2605 31807
rect 2605 31773 2639 31807
rect 2639 31773 2648 31807
rect 2596 31764 2648 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 26056 31288 26108 31340
rect 940 31220 992 31272
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 940 30608 992 30660
rect 1860 30540 1912 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 10416 30268 10468 30320
rect 940 30132 992 30184
rect 1032 30064 1084 30116
rect 10784 30064 10836 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12440 29588 12492 29640
rect 25596 29588 25648 29640
rect 940 29520 992 29572
rect 2412 29520 2464 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 13544 29180 13596 29232
rect 1032 29044 1084 29096
rect 940 28976 992 29028
rect 6460 28976 6512 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 940 28432 992 28484
rect 4620 28432 4672 28484
rect 10692 28432 10744 28484
rect 31944 28364 31996 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4068 28092 4120 28144
rect 940 27956 992 28008
rect 1032 27888 1084 27940
rect 4620 27888 4672 27940
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 10324 27548 10376 27600
rect 11244 27548 11296 27600
rect 940 27344 992 27396
rect 20628 27412 20680 27464
rect 1952 27319 2004 27328
rect 1952 27285 1961 27319
rect 1961 27285 1995 27319
rect 1995 27285 2004 27319
rect 1952 27276 2004 27285
rect 19064 27276 19116 27328
rect 19984 27276 20036 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1952 27072 2004 27124
rect 19340 27072 19392 27124
rect 19984 27072 20036 27124
rect 20628 27115 20680 27124
rect 20628 27081 20637 27115
rect 20637 27081 20671 27115
rect 20671 27081 20680 27115
rect 20628 27072 20680 27081
rect 1032 27004 1084 27056
rect 5264 27004 5316 27056
rect 33784 27004 33836 27056
rect 3976 26936 4028 26988
rect 14648 26979 14700 26988
rect 14648 26945 14657 26979
rect 14657 26945 14691 26979
rect 14691 26945 14700 26979
rect 14648 26936 14700 26945
rect 1124 26868 1176 26920
rect 4068 26868 4120 26920
rect 14096 26868 14148 26920
rect 2780 26843 2832 26852
rect 2780 26809 2789 26843
rect 2789 26809 2823 26843
rect 2823 26809 2832 26843
rect 2780 26800 2832 26809
rect 15936 26936 15988 26988
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 14924 26911 14976 26920
rect 14924 26877 14933 26911
rect 14933 26877 14967 26911
rect 14967 26877 14976 26911
rect 14924 26868 14976 26877
rect 20352 26936 20404 26988
rect 24952 26936 25004 26988
rect 34612 26979 34664 26988
rect 34612 26945 34621 26979
rect 34621 26945 34655 26979
rect 34655 26945 34664 26979
rect 34612 26936 34664 26945
rect 19800 26911 19852 26920
rect 19800 26877 19809 26911
rect 19809 26877 19843 26911
rect 19843 26877 19852 26911
rect 19800 26868 19852 26877
rect 19524 26800 19576 26852
rect 20444 26800 20496 26852
rect 34152 26868 34204 26920
rect 36360 26868 36412 26920
rect 14740 26775 14792 26784
rect 14740 26741 14749 26775
rect 14749 26741 14783 26775
rect 14783 26741 14792 26775
rect 14740 26732 14792 26741
rect 15384 26775 15436 26784
rect 15384 26741 15393 26775
rect 15393 26741 15427 26775
rect 15427 26741 15436 26775
rect 15384 26732 15436 26741
rect 19800 26732 19852 26784
rect 20536 26732 20588 26784
rect 20628 26732 20680 26784
rect 22008 26732 22060 26784
rect 24400 26775 24452 26784
rect 24400 26741 24409 26775
rect 24409 26741 24443 26775
rect 24443 26741 24452 26775
rect 24400 26732 24452 26741
rect 24584 26732 24636 26784
rect 34428 26775 34480 26784
rect 34428 26741 34437 26775
rect 34437 26741 34471 26775
rect 34471 26741 34480 26775
rect 34428 26732 34480 26741
rect 34796 26775 34848 26784
rect 34796 26741 34805 26775
rect 34805 26741 34839 26775
rect 34839 26741 34848 26775
rect 34796 26732 34848 26741
rect 35808 26732 35860 26784
rect 38016 26732 38068 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5264 26528 5316 26580
rect 14832 26528 14884 26580
rect 15936 26571 15988 26580
rect 15936 26537 15945 26571
rect 15945 26537 15979 26571
rect 15979 26537 15988 26571
rect 15936 26528 15988 26537
rect 20076 26528 20128 26580
rect 37832 26528 37884 26580
rect 14740 26460 14792 26512
rect 20628 26460 20680 26512
rect 2504 26392 2556 26444
rect 4344 26392 4396 26444
rect 6460 26435 6512 26444
rect 6460 26401 6469 26435
rect 6469 26401 6503 26435
rect 6503 26401 6512 26435
rect 6460 26392 6512 26401
rect 8024 26435 8076 26444
rect 8024 26401 8033 26435
rect 8033 26401 8067 26435
rect 8067 26401 8076 26435
rect 8024 26392 8076 26401
rect 6644 26324 6696 26376
rect 940 26256 992 26308
rect 7656 26256 7708 26308
rect 2320 26188 2372 26240
rect 3424 26188 3476 26240
rect 6000 26231 6052 26240
rect 6000 26197 6009 26231
rect 6009 26197 6043 26231
rect 6043 26197 6052 26231
rect 6000 26188 6052 26197
rect 6368 26231 6420 26240
rect 6368 26197 6377 26231
rect 6377 26197 6411 26231
rect 6411 26197 6420 26231
rect 6368 26188 6420 26197
rect 7472 26231 7524 26240
rect 7472 26197 7481 26231
rect 7481 26197 7515 26231
rect 7515 26197 7524 26231
rect 7472 26188 7524 26197
rect 14740 26367 14792 26376
rect 14740 26333 14749 26367
rect 14749 26333 14783 26367
rect 14783 26333 14792 26367
rect 14740 26324 14792 26333
rect 15016 26324 15068 26376
rect 20352 26367 20404 26376
rect 20352 26333 20361 26367
rect 20361 26333 20395 26367
rect 20395 26333 20404 26367
rect 20352 26324 20404 26333
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 13636 26299 13688 26308
rect 13636 26265 13645 26299
rect 13645 26265 13679 26299
rect 13679 26265 13688 26299
rect 13636 26256 13688 26265
rect 14648 26256 14700 26308
rect 15108 26188 15160 26240
rect 15660 26256 15712 26308
rect 19248 26256 19300 26308
rect 20628 26367 20680 26376
rect 20628 26333 20637 26367
rect 20637 26333 20671 26367
rect 20671 26333 20680 26367
rect 20628 26324 20680 26333
rect 20720 26324 20772 26376
rect 15844 26188 15896 26240
rect 24860 26460 24912 26512
rect 33508 26503 33560 26512
rect 33508 26469 33517 26503
rect 33517 26469 33551 26503
rect 33551 26469 33560 26503
rect 33508 26460 33560 26469
rect 24400 26392 24452 26444
rect 22008 26367 22060 26376
rect 22008 26333 22017 26367
rect 22017 26333 22051 26367
rect 22051 26333 22060 26367
rect 22008 26324 22060 26333
rect 22284 26367 22336 26376
rect 22284 26333 22293 26367
rect 22293 26333 22327 26367
rect 22327 26333 22336 26367
rect 22284 26324 22336 26333
rect 24584 26367 24636 26376
rect 24584 26333 24593 26367
rect 24593 26333 24627 26367
rect 24627 26333 24636 26367
rect 24584 26324 24636 26333
rect 28264 26392 28316 26444
rect 28724 26392 28776 26444
rect 32128 26324 32180 26376
rect 21548 26231 21600 26240
rect 21548 26197 21557 26231
rect 21557 26197 21591 26231
rect 21591 26197 21600 26231
rect 21548 26188 21600 26197
rect 24952 26256 25004 26308
rect 25964 26256 26016 26308
rect 32496 26392 32548 26444
rect 32312 26367 32364 26376
rect 32312 26333 32321 26367
rect 32321 26333 32355 26367
rect 32355 26333 32364 26367
rect 32312 26324 32364 26333
rect 34152 26367 34204 26376
rect 34152 26333 34161 26367
rect 34161 26333 34195 26367
rect 34195 26333 34204 26367
rect 34152 26324 34204 26333
rect 34428 26324 34480 26376
rect 35256 26367 35308 26376
rect 35256 26333 35265 26367
rect 35265 26333 35299 26367
rect 35299 26333 35308 26367
rect 35256 26324 35308 26333
rect 37648 26324 37700 26376
rect 37832 26324 37884 26376
rect 38016 26367 38068 26376
rect 38016 26333 38025 26367
rect 38025 26333 38059 26367
rect 38059 26333 38068 26367
rect 38016 26324 38068 26333
rect 38844 26392 38896 26444
rect 39212 26392 39264 26444
rect 40316 26460 40368 26512
rect 39396 26392 39448 26444
rect 32680 26299 32732 26308
rect 32680 26265 32689 26299
rect 32689 26265 32723 26299
rect 32723 26265 32732 26299
rect 32680 26256 32732 26265
rect 33692 26256 33744 26308
rect 34796 26256 34848 26308
rect 34980 26256 35032 26308
rect 36360 26299 36412 26308
rect 36360 26265 36394 26299
rect 36394 26265 36412 26299
rect 40040 26367 40092 26376
rect 40040 26333 40049 26367
rect 40049 26333 40083 26367
rect 40083 26333 40092 26367
rect 40040 26324 40092 26333
rect 40224 26367 40276 26376
rect 40224 26333 40233 26367
rect 40233 26333 40267 26367
rect 40267 26333 40276 26367
rect 40224 26324 40276 26333
rect 36360 26256 36412 26265
rect 36544 26231 36596 26240
rect 36544 26197 36553 26231
rect 36553 26197 36587 26231
rect 36587 26197 36596 26231
rect 36544 26188 36596 26197
rect 40132 26256 40184 26308
rect 38752 26188 38804 26240
rect 40040 26188 40092 26240
rect 40408 26367 40460 26376
rect 40408 26333 40417 26367
rect 40417 26333 40451 26367
rect 40451 26333 40460 26367
rect 40408 26324 40460 26333
rect 40868 26256 40920 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4620 25984 4672 26036
rect 8024 26027 8076 26036
rect 8024 25993 8033 26027
rect 8033 25993 8067 26027
rect 8067 25993 8076 26027
rect 8024 25984 8076 25993
rect 10692 26027 10744 26036
rect 10692 25993 10701 26027
rect 10701 25993 10735 26027
rect 10735 25993 10744 26027
rect 10692 25984 10744 25993
rect 15108 26027 15160 26036
rect 15108 25993 15117 26027
rect 15117 25993 15151 26027
rect 15151 25993 15160 26027
rect 15108 25984 15160 25993
rect 20444 25984 20496 26036
rect 34888 25984 34940 26036
rect 36544 25984 36596 26036
rect 1124 25916 1176 25968
rect 19248 25916 19300 25968
rect 1032 25780 1084 25832
rect 4988 25848 5040 25900
rect 7380 25848 7432 25900
rect 10692 25848 10744 25900
rect 14740 25848 14792 25900
rect 15844 25848 15896 25900
rect 30288 25916 30340 25968
rect 4344 25823 4396 25832
rect 4344 25789 4353 25823
rect 4353 25789 4387 25823
rect 4387 25789 4396 25823
rect 4344 25780 4396 25789
rect 8024 25780 8076 25832
rect 10876 25780 10928 25832
rect 14924 25780 14976 25832
rect 15936 25780 15988 25832
rect 17776 25780 17828 25832
rect 29000 25780 29052 25832
rect 30104 25891 30156 25900
rect 30104 25857 30113 25891
rect 30113 25857 30147 25891
rect 30147 25857 30156 25891
rect 30104 25848 30156 25857
rect 30196 25891 30248 25900
rect 30196 25857 30205 25891
rect 30205 25857 30239 25891
rect 30239 25857 30248 25891
rect 30196 25848 30248 25857
rect 3884 25644 3936 25696
rect 4620 25712 4672 25764
rect 19340 25712 19392 25764
rect 30840 25712 30892 25764
rect 32128 25848 32180 25900
rect 32496 25891 32548 25900
rect 32496 25857 32505 25891
rect 32505 25857 32539 25891
rect 32539 25857 32548 25891
rect 32496 25848 32548 25857
rect 33508 25848 33560 25900
rect 33692 25891 33744 25900
rect 33692 25857 33701 25891
rect 33701 25857 33735 25891
rect 33735 25857 33744 25891
rect 33692 25848 33744 25857
rect 37372 25916 37424 25968
rect 38844 25959 38896 25968
rect 38844 25925 38853 25959
rect 38853 25925 38887 25959
rect 38887 25925 38896 25959
rect 38844 25916 38896 25925
rect 40132 25984 40184 26036
rect 40224 25916 40276 25968
rect 35256 25848 35308 25900
rect 35900 25780 35952 25832
rect 6736 25644 6788 25696
rect 10232 25687 10284 25696
rect 10232 25653 10241 25687
rect 10241 25653 10275 25687
rect 10275 25653 10284 25687
rect 10232 25644 10284 25653
rect 15016 25644 15068 25696
rect 19616 25644 19668 25696
rect 29920 25644 29972 25696
rect 35256 25712 35308 25764
rect 36176 25891 36228 25900
rect 36176 25857 36185 25891
rect 36185 25857 36219 25891
rect 36219 25857 36228 25891
rect 36176 25848 36228 25857
rect 38752 25891 38804 25900
rect 38752 25857 38761 25891
rect 38761 25857 38795 25891
rect 38795 25857 38804 25891
rect 38752 25848 38804 25857
rect 37648 25780 37700 25832
rect 39212 25891 39264 25900
rect 39212 25857 39221 25891
rect 39221 25857 39255 25891
rect 39255 25857 39264 25891
rect 39212 25848 39264 25857
rect 40040 25891 40092 25900
rect 40040 25857 40049 25891
rect 40049 25857 40083 25891
rect 40083 25857 40092 25891
rect 40040 25848 40092 25857
rect 40316 25848 40368 25900
rect 40408 25780 40460 25832
rect 41052 25823 41104 25832
rect 41052 25789 41061 25823
rect 41061 25789 41095 25823
rect 41095 25789 41104 25823
rect 41052 25780 41104 25789
rect 42616 25891 42668 25900
rect 42616 25857 42625 25891
rect 42625 25857 42659 25891
rect 42659 25857 42668 25891
rect 42616 25848 42668 25857
rect 36084 25687 36136 25696
rect 36084 25653 36093 25687
rect 36093 25653 36127 25687
rect 36127 25653 36136 25687
rect 36084 25644 36136 25653
rect 40132 25687 40184 25696
rect 40132 25653 40141 25687
rect 40141 25653 40175 25687
rect 40175 25653 40184 25687
rect 40132 25644 40184 25653
rect 41236 25687 41288 25696
rect 41236 25653 41245 25687
rect 41245 25653 41279 25687
rect 41279 25653 41288 25687
rect 41236 25644 41288 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 6368 25440 6420 25492
rect 7196 25440 7248 25492
rect 15844 25440 15896 25492
rect 22284 25483 22336 25492
rect 22284 25449 22293 25483
rect 22293 25449 22327 25483
rect 22327 25449 22336 25483
rect 22284 25440 22336 25449
rect 25964 25483 26016 25492
rect 25964 25449 25973 25483
rect 25973 25449 26007 25483
rect 26007 25449 26016 25483
rect 25964 25440 26016 25449
rect 34612 25440 34664 25492
rect 39948 25440 40000 25492
rect 41052 25440 41104 25492
rect 36544 25415 36596 25424
rect 36544 25381 36553 25415
rect 36553 25381 36587 25415
rect 36587 25381 36596 25415
rect 36544 25372 36596 25381
rect 10784 25347 10836 25356
rect 10784 25313 10793 25347
rect 10793 25313 10827 25347
rect 10827 25313 10836 25347
rect 10784 25304 10836 25313
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 28908 25304 28960 25356
rect 32956 25304 33008 25356
rect 36084 25304 36136 25356
rect 36820 25304 36872 25356
rect 2044 25279 2096 25288
rect 2044 25245 2053 25279
rect 2053 25245 2087 25279
rect 2087 25245 2096 25279
rect 2044 25236 2096 25245
rect 2320 25279 2372 25288
rect 2320 25245 2354 25279
rect 2354 25245 2372 25279
rect 2320 25236 2372 25245
rect 3608 25236 3660 25288
rect 6552 25236 6604 25288
rect 7472 25279 7524 25288
rect 7472 25245 7506 25279
rect 7506 25245 7524 25279
rect 7472 25236 7524 25245
rect 15016 25236 15068 25288
rect 19432 25279 19484 25288
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 19616 25279 19668 25288
rect 19616 25245 19625 25279
rect 19625 25245 19659 25279
rect 19659 25245 19668 25279
rect 19616 25236 19668 25245
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 21548 25236 21600 25288
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 24860 25279 24912 25288
rect 24860 25245 24894 25279
rect 24894 25245 24912 25279
rect 24860 25236 24912 25245
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 37648 25236 37700 25288
rect 38752 25236 38804 25288
rect 6000 25168 6052 25220
rect 15384 25168 15436 25220
rect 3424 25143 3476 25152
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 7656 25100 7708 25152
rect 10324 25143 10376 25152
rect 10324 25109 10333 25143
rect 10333 25109 10367 25143
rect 10367 25109 10376 25143
rect 10324 25100 10376 25109
rect 10784 25100 10836 25152
rect 19340 25100 19392 25152
rect 30380 25100 30432 25152
rect 37280 25100 37332 25152
rect 37924 25143 37976 25152
rect 37924 25109 37933 25143
rect 37933 25109 37967 25143
rect 37967 25109 37976 25143
rect 37924 25100 37976 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4988 24939 5040 24948
rect 4988 24905 4997 24939
rect 4997 24905 5031 24939
rect 5031 24905 5040 24939
rect 4988 24896 5040 24905
rect 20444 24896 20496 24948
rect 30012 24896 30064 24948
rect 37648 24896 37700 24948
rect 38384 24896 38436 24948
rect 10232 24828 10284 24880
rect 940 24760 992 24812
rect 1032 24692 1084 24744
rect 3884 24803 3936 24812
rect 3884 24769 3918 24803
rect 3918 24769 3936 24803
rect 3884 24760 3936 24769
rect 15016 24828 15068 24880
rect 13636 24803 13688 24812
rect 13636 24769 13670 24803
rect 13670 24769 13688 24803
rect 13636 24760 13688 24769
rect 16120 24760 16172 24812
rect 19064 24803 19116 24812
rect 19064 24769 19098 24803
rect 19098 24769 19116 24803
rect 19064 24760 19116 24769
rect 19616 24760 19668 24812
rect 20628 24760 20680 24812
rect 24584 24828 24636 24880
rect 30104 24828 30156 24880
rect 33508 24828 33560 24880
rect 34612 24871 34664 24880
rect 34612 24837 34621 24871
rect 34621 24837 34655 24871
rect 34655 24837 34664 24871
rect 34612 24828 34664 24837
rect 39212 24896 39264 24948
rect 24768 24760 24820 24812
rect 27712 24760 27764 24812
rect 28908 24760 28960 24812
rect 29920 24803 29972 24812
rect 29920 24769 29929 24803
rect 29929 24769 29963 24803
rect 29963 24769 29972 24803
rect 29920 24760 29972 24769
rect 30288 24760 30340 24812
rect 30380 24803 30432 24812
rect 30380 24769 30389 24803
rect 30389 24769 30423 24803
rect 30423 24769 30432 24803
rect 30380 24760 30432 24769
rect 32496 24803 32548 24812
rect 32496 24769 32505 24803
rect 32505 24769 32539 24803
rect 32539 24769 32548 24803
rect 32496 24760 32548 24769
rect 32588 24803 32640 24812
rect 32588 24769 32597 24803
rect 32597 24769 32631 24803
rect 32631 24769 32640 24803
rect 32588 24760 32640 24769
rect 33048 24760 33100 24812
rect 34428 24803 34480 24812
rect 34428 24769 34437 24803
rect 34437 24769 34471 24803
rect 34471 24769 34480 24803
rect 34428 24760 34480 24769
rect 36360 24760 36412 24812
rect 37924 24760 37976 24812
rect 38752 24803 38804 24812
rect 38752 24769 38761 24803
rect 38761 24769 38795 24803
rect 38795 24769 38804 24803
rect 38752 24760 38804 24769
rect 40316 24760 40368 24812
rect 40868 24803 40920 24812
rect 40868 24769 40902 24803
rect 40902 24769 40920 24803
rect 40868 24760 40920 24769
rect 2044 24692 2096 24744
rect 3608 24735 3660 24744
rect 3608 24701 3617 24735
rect 3617 24701 3651 24735
rect 3651 24701 3660 24735
rect 3608 24692 3660 24701
rect 9680 24692 9732 24744
rect 3516 24624 3568 24676
rect 2228 24556 2280 24608
rect 2596 24556 2648 24608
rect 4896 24556 4948 24608
rect 10692 24556 10744 24608
rect 14740 24599 14792 24608
rect 14740 24565 14749 24599
rect 14749 24565 14783 24599
rect 14783 24565 14792 24599
rect 14740 24556 14792 24565
rect 15016 24556 15068 24608
rect 17868 24556 17920 24608
rect 18788 24556 18840 24608
rect 20904 24624 20956 24676
rect 28816 24692 28868 24744
rect 20352 24556 20404 24608
rect 25596 24599 25648 24608
rect 25596 24565 25605 24599
rect 25605 24565 25639 24599
rect 25639 24565 25648 24599
rect 25596 24556 25648 24565
rect 29736 24624 29788 24676
rect 33784 24624 33836 24676
rect 35716 24624 35768 24676
rect 40592 24735 40644 24744
rect 40592 24701 40601 24735
rect 40601 24701 40635 24735
rect 40635 24701 40644 24735
rect 40592 24692 40644 24701
rect 28816 24556 28868 24608
rect 29368 24556 29420 24608
rect 32220 24556 32272 24608
rect 33140 24556 33192 24608
rect 39120 24556 39172 24608
rect 40040 24556 40092 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1952 24352 2004 24404
rect 15936 24395 15988 24404
rect 15936 24361 15945 24395
rect 15945 24361 15979 24395
rect 15979 24361 15988 24395
rect 15936 24352 15988 24361
rect 16120 24395 16172 24404
rect 16120 24361 16129 24395
rect 16129 24361 16163 24395
rect 16163 24361 16172 24395
rect 16120 24352 16172 24361
rect 19432 24284 19484 24336
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 29000 24352 29052 24404
rect 36360 24352 36412 24404
rect 38384 24395 38436 24404
rect 38384 24361 38393 24395
rect 38393 24361 38427 24395
rect 38427 24361 38436 24395
rect 38384 24352 38436 24361
rect 42616 24352 42668 24404
rect 29460 24284 29512 24336
rect 32404 24284 32456 24336
rect 14740 24216 14792 24268
rect 19708 24216 19760 24268
rect 20904 24216 20956 24268
rect 24584 24216 24636 24268
rect 1676 24148 1728 24200
rect 2044 24191 2096 24200
rect 2044 24157 2053 24191
rect 2053 24157 2087 24191
rect 2087 24157 2096 24191
rect 2044 24148 2096 24157
rect 4620 24148 4672 24200
rect 2504 24080 2556 24132
rect 9680 24148 9732 24200
rect 10324 24148 10376 24200
rect 15568 24191 15620 24200
rect 15568 24157 15577 24191
rect 15577 24157 15611 24191
rect 15611 24157 15620 24191
rect 15568 24148 15620 24157
rect 17868 24148 17920 24200
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 31760 24216 31812 24268
rect 32588 24216 32640 24268
rect 27712 24148 27764 24200
rect 32956 24148 33008 24200
rect 33140 24191 33192 24200
rect 33140 24157 33174 24191
rect 33174 24157 33192 24191
rect 33140 24148 33192 24157
rect 36544 24148 36596 24200
rect 37280 24191 37332 24200
rect 37280 24157 37314 24191
rect 37314 24157 37332 24191
rect 37280 24148 37332 24157
rect 39120 24191 39172 24200
rect 39120 24157 39129 24191
rect 39129 24157 39163 24191
rect 39163 24157 39172 24191
rect 39120 24148 39172 24157
rect 40132 24148 40184 24200
rect 40224 24148 40276 24200
rect 40592 24148 40644 24200
rect 41236 24191 41288 24200
rect 41236 24157 41270 24191
rect 41270 24157 41288 24191
rect 41236 24148 41288 24157
rect 11336 24080 11388 24132
rect 16580 24080 16632 24132
rect 4804 24012 4856 24064
rect 10784 24012 10836 24064
rect 19616 24055 19668 24064
rect 19616 24021 19625 24055
rect 19625 24021 19659 24055
rect 19659 24021 19668 24055
rect 19616 24012 19668 24021
rect 19708 24055 19760 24064
rect 19708 24021 19717 24055
rect 19717 24021 19751 24055
rect 19751 24021 19760 24055
rect 19708 24012 19760 24021
rect 20536 24080 20588 24132
rect 25596 24080 25648 24132
rect 26148 24080 26200 24132
rect 34796 24080 34848 24132
rect 36176 24080 36228 24132
rect 20996 24012 21048 24064
rect 30564 24012 30616 24064
rect 34612 24012 34664 24064
rect 38936 24012 38988 24064
rect 39396 24055 39448 24064
rect 39396 24021 39405 24055
rect 39405 24021 39439 24055
rect 39439 24021 39448 24055
rect 39396 24012 39448 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 1952 23851 2004 23860
rect 1952 23817 1961 23851
rect 1961 23817 1995 23851
rect 1995 23817 2004 23851
rect 1952 23808 2004 23817
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 2780 23808 2832 23860
rect 3516 23808 3568 23860
rect 4988 23740 5040 23792
rect 940 23672 992 23724
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 6644 23672 6696 23724
rect 17040 23740 17092 23792
rect 20076 23783 20128 23792
rect 20076 23749 20085 23783
rect 20085 23749 20119 23783
rect 20119 23749 20128 23783
rect 20076 23740 20128 23749
rect 20536 23783 20588 23792
rect 20536 23749 20545 23783
rect 20545 23749 20579 23783
rect 20579 23749 20588 23783
rect 20536 23740 20588 23749
rect 26148 23851 26200 23860
rect 26148 23817 26157 23851
rect 26157 23817 26191 23851
rect 26191 23817 26200 23851
rect 26148 23808 26200 23817
rect 17868 23672 17920 23724
rect 2964 23604 3016 23656
rect 4804 23604 4856 23656
rect 17132 23604 17184 23656
rect 20444 23647 20496 23656
rect 20444 23613 20453 23647
rect 20453 23613 20487 23647
rect 20487 23613 20496 23647
rect 20444 23604 20496 23613
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 26332 23715 26384 23724
rect 26332 23681 26341 23715
rect 26341 23681 26375 23715
rect 26375 23681 26384 23715
rect 26332 23672 26384 23681
rect 29368 23783 29420 23792
rect 29368 23749 29377 23783
rect 29377 23749 29411 23783
rect 29411 23749 29420 23783
rect 29368 23740 29420 23749
rect 31760 23851 31812 23860
rect 31760 23817 31769 23851
rect 31769 23817 31803 23851
rect 31803 23817 31812 23851
rect 31760 23808 31812 23817
rect 32496 23851 32548 23860
rect 32496 23817 32505 23851
rect 32505 23817 32539 23851
rect 32539 23817 32548 23851
rect 32496 23808 32548 23817
rect 40316 23808 40368 23860
rect 36728 23740 36780 23792
rect 39396 23740 39448 23792
rect 7748 23536 7800 23588
rect 9864 23536 9916 23588
rect 15568 23536 15620 23588
rect 28264 23536 28316 23588
rect 30196 23715 30248 23724
rect 30196 23681 30205 23715
rect 30205 23681 30239 23715
rect 30239 23681 30248 23715
rect 30196 23672 30248 23681
rect 30472 23672 30524 23724
rect 32312 23715 32364 23724
rect 32312 23681 32321 23715
rect 32321 23681 32355 23715
rect 32355 23681 32364 23715
rect 32312 23672 32364 23681
rect 31760 23604 31812 23656
rect 34612 23672 34664 23724
rect 33324 23647 33376 23656
rect 33324 23613 33333 23647
rect 33333 23613 33367 23647
rect 33367 23613 33376 23647
rect 33324 23604 33376 23613
rect 40224 23604 40276 23656
rect 31208 23536 31260 23588
rect 33048 23536 33100 23588
rect 5080 23468 5132 23520
rect 6552 23468 6604 23520
rect 11704 23468 11756 23520
rect 13452 23468 13504 23520
rect 16856 23468 16908 23520
rect 17776 23468 17828 23520
rect 18880 23468 18932 23520
rect 26516 23511 26568 23520
rect 26516 23477 26525 23511
rect 26525 23477 26559 23511
rect 26559 23477 26568 23511
rect 26516 23468 26568 23477
rect 29000 23468 29052 23520
rect 32312 23468 32364 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6644 23264 6696 23316
rect 7196 23264 7248 23316
rect 13544 23307 13596 23316
rect 13544 23273 13553 23307
rect 13553 23273 13587 23307
rect 13587 23273 13596 23307
rect 13544 23264 13596 23273
rect 16580 23307 16632 23316
rect 16580 23273 16589 23307
rect 16589 23273 16623 23307
rect 16623 23273 16632 23307
rect 16580 23264 16632 23273
rect 3424 23196 3476 23248
rect 1032 23128 1084 23180
rect 2964 23128 3016 23180
rect 7288 23128 7340 23180
rect 16948 23196 17000 23248
rect 17040 23196 17092 23248
rect 26516 23264 26568 23316
rect 29736 23307 29788 23316
rect 29736 23273 29745 23307
rect 29745 23273 29779 23307
rect 29779 23273 29788 23307
rect 29736 23264 29788 23273
rect 33048 23264 33100 23316
rect 42156 23307 42208 23316
rect 42156 23273 42165 23307
rect 42165 23273 42199 23307
rect 42199 23273 42208 23307
rect 42156 23264 42208 23273
rect 28724 23196 28776 23248
rect 30564 23196 30616 23248
rect 7656 23171 7708 23180
rect 7656 23137 7665 23171
rect 7665 23137 7699 23171
rect 7699 23137 7708 23171
rect 7656 23128 7708 23137
rect 940 22924 992 22976
rect 5172 22992 5224 23044
rect 6736 23035 6788 23044
rect 6736 23001 6745 23035
rect 6745 23001 6779 23035
rect 6779 23001 6788 23035
rect 6736 22992 6788 23001
rect 7748 23103 7800 23112
rect 7748 23069 7757 23103
rect 7757 23069 7791 23103
rect 7791 23069 7800 23103
rect 7748 23060 7800 23069
rect 12900 23060 12952 23112
rect 16764 23103 16816 23112
rect 16764 23069 16773 23103
rect 16773 23069 16807 23103
rect 16807 23069 16816 23103
rect 16764 23060 16816 23069
rect 16856 23103 16908 23112
rect 16856 23069 16865 23103
rect 16865 23069 16899 23103
rect 16899 23069 16908 23103
rect 16856 23060 16908 23069
rect 2412 22924 2464 22976
rect 4436 22967 4488 22976
rect 4436 22933 4445 22967
rect 4445 22933 4479 22967
rect 4479 22933 4488 22967
rect 4436 22924 4488 22933
rect 4896 22967 4948 22976
rect 4896 22933 4905 22967
rect 4905 22933 4939 22967
rect 4939 22933 4948 22967
rect 4896 22924 4948 22933
rect 6644 22967 6696 22976
rect 6644 22933 6653 22967
rect 6653 22933 6687 22967
rect 6687 22933 6696 22967
rect 6644 22924 6696 22933
rect 8208 22924 8260 22976
rect 12808 22992 12860 23044
rect 14648 22992 14700 23044
rect 16856 22924 16908 22976
rect 17132 23060 17184 23112
rect 17776 23060 17828 23112
rect 28264 23128 28316 23180
rect 20812 23060 20864 23112
rect 22192 23060 22244 23112
rect 20260 22992 20312 23044
rect 20444 22992 20496 23044
rect 21364 22992 21416 23044
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 28448 23103 28500 23112
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 22100 22924 22152 22976
rect 28724 23103 28776 23112
rect 28724 23069 28733 23103
rect 28733 23069 28767 23103
rect 28767 23069 28776 23103
rect 28724 23060 28776 23069
rect 35900 23128 35952 23180
rect 36268 23128 36320 23180
rect 30012 23103 30064 23112
rect 30012 23069 30021 23103
rect 30021 23069 30055 23103
rect 30055 23069 30064 23103
rect 30012 23060 30064 23069
rect 30656 23060 30708 23112
rect 29184 22992 29236 23044
rect 31392 22992 31444 23044
rect 32128 23060 32180 23112
rect 33324 23060 33376 23112
rect 35440 23060 35492 23112
rect 36176 23060 36228 23112
rect 37372 23128 37424 23180
rect 34520 22992 34572 23044
rect 36820 23103 36872 23112
rect 36820 23069 36829 23103
rect 36829 23069 36863 23103
rect 36863 23069 36872 23103
rect 36820 23060 36872 23069
rect 40224 23060 40276 23112
rect 38844 22992 38896 23044
rect 28356 22924 28408 22976
rect 29092 22924 29144 22976
rect 36820 22924 36872 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2412 22763 2464 22772
rect 2412 22729 2421 22763
rect 2421 22729 2455 22763
rect 2455 22729 2464 22763
rect 2412 22720 2464 22729
rect 5172 22720 5224 22772
rect 12808 22763 12860 22772
rect 12808 22729 12817 22763
rect 12817 22729 12851 22763
rect 12851 22729 12860 22763
rect 12808 22720 12860 22729
rect 13544 22720 13596 22772
rect 18420 22720 18472 22772
rect 18880 22720 18932 22772
rect 23756 22763 23808 22772
rect 23756 22729 23765 22763
rect 23765 22729 23799 22763
rect 23799 22729 23808 22763
rect 23756 22720 23808 22729
rect 26056 22720 26108 22772
rect 28448 22720 28500 22772
rect 4436 22652 4488 22704
rect 3056 22584 3108 22636
rect 3240 22627 3292 22636
rect 3240 22593 3249 22627
rect 3249 22593 3283 22627
rect 3283 22593 3292 22627
rect 3240 22584 3292 22593
rect 3608 22584 3660 22636
rect 10784 22652 10836 22704
rect 14372 22652 14424 22704
rect 22192 22652 22244 22704
rect 8208 22627 8260 22636
rect 8208 22593 8217 22627
rect 8217 22593 8251 22627
rect 8251 22593 8260 22627
rect 8208 22584 8260 22593
rect 9036 22584 9088 22636
rect 9680 22627 9732 22636
rect 9680 22593 9714 22627
rect 9714 22593 9732 22627
rect 9680 22584 9732 22593
rect 13084 22584 13136 22636
rect 13268 22627 13320 22636
rect 13268 22593 13277 22627
rect 13277 22593 13311 22627
rect 13311 22593 13320 22627
rect 13268 22584 13320 22593
rect 2596 22559 2648 22568
rect 2596 22525 2605 22559
rect 2605 22525 2639 22559
rect 2639 22525 2648 22559
rect 2596 22516 2648 22525
rect 2964 22516 3016 22568
rect 9404 22559 9456 22568
rect 9404 22525 9413 22559
rect 9413 22525 9447 22559
rect 9447 22525 9456 22559
rect 9404 22516 9456 22525
rect 12900 22516 12952 22568
rect 15016 22584 15068 22636
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17776 22584 17828 22636
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 22284 22584 22336 22636
rect 29184 22695 29236 22704
rect 29184 22661 29193 22695
rect 29193 22661 29227 22695
rect 29227 22661 29236 22695
rect 29184 22652 29236 22661
rect 23388 22584 23440 22636
rect 24584 22584 24636 22636
rect 25044 22627 25096 22636
rect 25044 22593 25078 22627
rect 25078 22593 25096 22627
rect 25044 22584 25096 22593
rect 1952 22423 2004 22432
rect 1952 22389 1961 22423
rect 1961 22389 1995 22423
rect 1995 22389 2004 22423
rect 1952 22380 2004 22389
rect 3332 22423 3384 22432
rect 3332 22389 3341 22423
rect 3341 22389 3375 22423
rect 3375 22389 3384 22423
rect 3332 22380 3384 22389
rect 6736 22380 6788 22432
rect 10416 22448 10468 22500
rect 19340 22516 19392 22568
rect 16856 22448 16908 22500
rect 20352 22448 20404 22500
rect 30012 22720 30064 22772
rect 31760 22720 31812 22772
rect 35808 22652 35860 22704
rect 10692 22380 10744 22432
rect 16948 22380 17000 22432
rect 19708 22380 19760 22432
rect 30196 22380 30248 22432
rect 30564 22380 30616 22432
rect 32312 22380 32364 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3056 22219 3108 22228
rect 3056 22185 3065 22219
rect 3065 22185 3099 22219
rect 3099 22185 3108 22219
rect 3056 22176 3108 22185
rect 5172 22219 5224 22228
rect 5172 22185 5181 22219
rect 5181 22185 5215 22219
rect 5215 22185 5224 22219
rect 5172 22176 5224 22185
rect 9680 22176 9732 22228
rect 19340 22176 19392 22228
rect 23388 22219 23440 22228
rect 23388 22185 23397 22219
rect 23397 22185 23431 22219
rect 23431 22185 23440 22219
rect 23388 22176 23440 22185
rect 25044 22176 25096 22228
rect 27528 22176 27580 22228
rect 29184 22176 29236 22228
rect 30288 22176 30340 22228
rect 30840 22219 30892 22228
rect 30840 22185 30849 22219
rect 30849 22185 30883 22219
rect 30883 22185 30892 22219
rect 30840 22176 30892 22185
rect 31484 22176 31536 22228
rect 37464 22176 37516 22228
rect 4804 22040 4856 22092
rect 16764 22108 16816 22160
rect 19708 22108 19760 22160
rect 20076 22108 20128 22160
rect 30656 22108 30708 22160
rect 1676 22015 1728 22024
rect 1676 21981 1685 22015
rect 1685 21981 1719 22015
rect 1719 21981 1728 22015
rect 1676 21972 1728 21981
rect 1952 22015 2004 22024
rect 1952 21981 1986 22015
rect 1986 21981 2004 22015
rect 1952 21972 2004 21981
rect 940 21904 992 21956
rect 4988 21904 5040 21956
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 5264 21972 5316 22024
rect 13176 22040 13228 22092
rect 13268 22040 13320 22092
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 11888 21904 11940 21956
rect 14096 21904 14148 21956
rect 17684 21972 17736 22024
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 22284 21972 22336 22024
rect 23480 21972 23532 22024
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 2228 21836 2280 21888
rect 5264 21836 5316 21888
rect 6460 21836 6512 21888
rect 10416 21836 10468 21888
rect 14280 21879 14332 21888
rect 14280 21845 14289 21879
rect 14289 21845 14323 21879
rect 14323 21845 14332 21879
rect 14280 21836 14332 21845
rect 18052 21836 18104 21888
rect 22192 21904 22244 21956
rect 25228 21972 25280 22024
rect 25320 22015 25372 22024
rect 25320 21981 25329 22015
rect 25329 21981 25363 22015
rect 25363 21981 25372 22015
rect 25320 21972 25372 21981
rect 26332 22040 26384 22092
rect 27528 22040 27580 22092
rect 30196 22015 30248 22024
rect 30196 21981 30205 22015
rect 30205 21981 30239 22015
rect 30239 21981 30248 22015
rect 30196 21972 30248 21981
rect 26056 21904 26108 21956
rect 30748 21904 30800 21956
rect 20720 21836 20772 21888
rect 22284 21836 22336 21888
rect 22560 21836 22612 21888
rect 22836 21879 22888 21888
rect 22836 21845 22845 21879
rect 22845 21845 22879 21879
rect 22879 21845 22888 21879
rect 22836 21836 22888 21845
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 30104 21879 30156 21888
rect 30104 21845 30113 21879
rect 30113 21845 30147 21879
rect 30147 21845 30156 21879
rect 30104 21836 30156 21845
rect 30472 21836 30524 21888
rect 35808 22040 35860 22092
rect 36544 22083 36596 22092
rect 36544 22049 36553 22083
rect 36553 22049 36587 22083
rect 36587 22049 36596 22083
rect 36544 22040 36596 22049
rect 36820 22083 36872 22092
rect 36820 22049 36829 22083
rect 36829 22049 36863 22083
rect 36863 22049 36872 22083
rect 36820 22040 36872 22049
rect 32956 22015 33008 22024
rect 32956 21981 32965 22015
rect 32965 21981 32999 22015
rect 32999 21981 33008 22015
rect 32956 21972 33008 21981
rect 40224 22015 40276 22024
rect 40224 21981 40233 22015
rect 40233 21981 40267 22015
rect 40267 21981 40276 22015
rect 40224 21972 40276 21981
rect 33324 21904 33376 21956
rect 33600 21836 33652 21888
rect 34336 21879 34388 21888
rect 34336 21845 34345 21879
rect 34345 21845 34379 21879
rect 34379 21845 34388 21879
rect 34336 21836 34388 21845
rect 34796 21836 34848 21888
rect 40592 21904 40644 21956
rect 40960 21836 41012 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 940 21632 992 21684
rect 3240 21632 3292 21684
rect 3976 21632 4028 21684
rect 9680 21632 9732 21684
rect 8484 21564 8536 21616
rect 4068 21496 4120 21548
rect 5080 21539 5132 21548
rect 5080 21505 5089 21539
rect 5089 21505 5123 21539
rect 5123 21505 5132 21539
rect 5080 21496 5132 21505
rect 5540 21496 5592 21548
rect 1032 21428 1084 21480
rect 940 21360 992 21412
rect 3424 21428 3476 21480
rect 9496 21496 9548 21548
rect 9588 21539 9640 21548
rect 9588 21505 9597 21539
rect 9597 21505 9631 21539
rect 9631 21505 9640 21539
rect 9588 21496 9640 21505
rect 7196 21428 7248 21480
rect 32864 21632 32916 21684
rect 33324 21675 33376 21684
rect 33324 21641 33333 21675
rect 33333 21641 33367 21675
rect 33367 21641 33376 21675
rect 33324 21632 33376 21641
rect 34336 21632 34388 21684
rect 34704 21632 34756 21684
rect 11888 21607 11940 21616
rect 11888 21573 11897 21607
rect 11897 21573 11931 21607
rect 11931 21573 11940 21607
rect 11888 21564 11940 21573
rect 14280 21564 14332 21616
rect 15936 21564 15988 21616
rect 11520 21496 11572 21548
rect 12992 21496 13044 21548
rect 17960 21564 18012 21616
rect 20168 21564 20220 21616
rect 22100 21607 22152 21616
rect 22100 21573 22109 21607
rect 22109 21573 22143 21607
rect 22143 21573 22152 21607
rect 22100 21564 22152 21573
rect 20352 21496 20404 21548
rect 26332 21564 26384 21616
rect 29736 21564 29788 21616
rect 30840 21564 30892 21616
rect 34520 21564 34572 21616
rect 19984 21428 20036 21480
rect 20444 21428 20496 21480
rect 1860 21292 1912 21344
rect 5172 21335 5224 21344
rect 5172 21301 5181 21335
rect 5181 21301 5215 21335
rect 5215 21301 5224 21335
rect 5172 21292 5224 21301
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 6644 21335 6696 21344
rect 6644 21301 6653 21335
rect 6653 21301 6687 21335
rect 6687 21301 6696 21335
rect 6644 21292 6696 21301
rect 7196 21335 7248 21344
rect 7196 21301 7205 21335
rect 7205 21301 7239 21335
rect 7239 21301 7248 21335
rect 7196 21292 7248 21301
rect 8576 21292 8628 21344
rect 11060 21292 11112 21344
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 14096 21360 14148 21412
rect 18512 21360 18564 21412
rect 17776 21335 17828 21344
rect 17776 21301 17785 21335
rect 17785 21301 17819 21335
rect 17819 21301 17828 21335
rect 17776 21292 17828 21301
rect 20996 21292 21048 21344
rect 21640 21292 21692 21344
rect 27160 21496 27212 21548
rect 30656 21539 30708 21548
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 33508 21539 33560 21548
rect 33508 21505 33517 21539
rect 33517 21505 33551 21539
rect 33551 21505 33560 21539
rect 33508 21496 33560 21505
rect 33784 21539 33836 21548
rect 25872 21428 25924 21480
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 26240 21471 26292 21480
rect 26240 21437 26249 21471
rect 26249 21437 26283 21471
rect 26283 21437 26292 21471
rect 26240 21428 26292 21437
rect 27344 21471 27396 21480
rect 27344 21437 27353 21471
rect 27353 21437 27387 21471
rect 27387 21437 27396 21471
rect 27344 21428 27396 21437
rect 27068 21360 27120 21412
rect 27528 21471 27580 21480
rect 27528 21437 27537 21471
rect 27537 21437 27571 21471
rect 27571 21437 27580 21471
rect 27528 21428 27580 21437
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 28632 21471 28684 21480
rect 28632 21437 28641 21471
rect 28641 21437 28675 21471
rect 28675 21437 28684 21471
rect 28632 21428 28684 21437
rect 30840 21471 30892 21480
rect 30840 21437 30849 21471
rect 30849 21437 30883 21471
rect 30883 21437 30892 21471
rect 30840 21428 30892 21437
rect 31208 21428 31260 21480
rect 33784 21505 33793 21539
rect 33793 21505 33827 21539
rect 33827 21505 33836 21539
rect 33784 21496 33836 21505
rect 33876 21496 33928 21548
rect 34428 21539 34480 21548
rect 34428 21505 34437 21539
rect 34437 21505 34471 21539
rect 34471 21505 34480 21539
rect 34428 21496 34480 21505
rect 37372 21496 37424 21548
rect 34336 21471 34388 21480
rect 34336 21437 34345 21471
rect 34345 21437 34379 21471
rect 34379 21437 34388 21471
rect 34336 21428 34388 21437
rect 37556 21564 37608 21616
rect 40592 21675 40644 21684
rect 40592 21641 40601 21675
rect 40601 21641 40635 21675
rect 40635 21641 40644 21675
rect 40592 21632 40644 21641
rect 40960 21675 41012 21684
rect 40960 21641 40969 21675
rect 40969 21641 41003 21675
rect 41003 21641 41012 21675
rect 40960 21632 41012 21641
rect 40408 21428 40460 21480
rect 45192 21496 45244 21548
rect 45836 21428 45888 21480
rect 25780 21335 25832 21344
rect 25780 21301 25789 21335
rect 25789 21301 25823 21335
rect 25823 21301 25832 21335
rect 25780 21292 25832 21301
rect 25964 21292 26016 21344
rect 28540 21292 28592 21344
rect 30104 21292 30156 21344
rect 32864 21292 32916 21344
rect 41236 21292 41288 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 7748 21131 7800 21140
rect 7748 21097 7757 21131
rect 7757 21097 7791 21131
rect 7791 21097 7800 21131
rect 7748 21088 7800 21097
rect 10048 21088 10100 21140
rect 11980 21131 12032 21140
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 17960 21131 18012 21140
rect 17960 21097 17969 21131
rect 17969 21097 18003 21131
rect 18003 21097 18012 21131
rect 17960 21088 18012 21097
rect 18512 21131 18564 21140
rect 18512 21097 18521 21131
rect 18521 21097 18555 21131
rect 18555 21097 18564 21131
rect 18512 21088 18564 21097
rect 22192 21131 22244 21140
rect 22192 21097 22201 21131
rect 22201 21097 22235 21131
rect 22235 21097 22244 21131
rect 22192 21088 22244 21097
rect 23480 21131 23532 21140
rect 23480 21097 23489 21131
rect 23489 21097 23523 21131
rect 23523 21097 23532 21131
rect 23480 21088 23532 21097
rect 27528 21088 27580 21140
rect 25780 21020 25832 21072
rect 27252 21020 27304 21072
rect 30564 21063 30616 21072
rect 30564 21029 30573 21063
rect 30573 21029 30607 21063
rect 30607 21029 30616 21063
rect 30564 21020 30616 21029
rect 31208 21063 31260 21072
rect 31208 21029 31217 21063
rect 31217 21029 31251 21063
rect 31251 21029 31260 21063
rect 31208 21020 31260 21029
rect 34796 21088 34848 21140
rect 40960 21088 41012 21140
rect 43444 21020 43496 21072
rect 2596 20995 2648 21004
rect 2596 20961 2605 20995
rect 2605 20961 2639 20995
rect 2639 20961 2648 20995
rect 2596 20952 2648 20961
rect 1676 20884 1728 20936
rect 9404 20884 9456 20936
rect 12992 20884 13044 20936
rect 13176 20884 13228 20936
rect 18420 20927 18472 20936
rect 18420 20893 18429 20927
rect 18429 20893 18463 20927
rect 18463 20893 18472 20927
rect 18420 20884 18472 20893
rect 3332 20816 3384 20868
rect 6644 20859 6696 20868
rect 6644 20825 6678 20859
rect 6678 20825 6696 20859
rect 6644 20816 6696 20825
rect 9128 20859 9180 20868
rect 9128 20825 9137 20859
rect 9137 20825 9171 20859
rect 9171 20825 9180 20859
rect 9128 20816 9180 20825
rect 12348 20816 12400 20868
rect 15108 20816 15160 20868
rect 15292 20816 15344 20868
rect 17684 20816 17736 20868
rect 19248 20884 19300 20936
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 21364 20884 21416 20936
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 2228 20748 2280 20800
rect 3424 20748 3476 20800
rect 9588 20748 9640 20800
rect 12440 20748 12492 20800
rect 13268 20748 13320 20800
rect 18604 20748 18656 20800
rect 23204 20952 23256 21004
rect 25964 20995 26016 21004
rect 25964 20961 25973 20995
rect 25973 20961 26007 20995
rect 26007 20961 26016 20995
rect 25964 20952 26016 20961
rect 28540 20952 28592 21004
rect 28632 20952 28684 21004
rect 30932 20952 30984 21004
rect 32956 20995 33008 21004
rect 32956 20961 32965 20995
rect 32965 20961 32999 20995
rect 32999 20961 33008 20995
rect 32956 20952 33008 20961
rect 40224 20952 40276 21004
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 23756 20927 23808 20936
rect 23756 20893 23765 20927
rect 23765 20893 23799 20927
rect 23799 20893 23808 20927
rect 23756 20884 23808 20893
rect 23572 20816 23624 20868
rect 26056 20927 26108 20936
rect 26056 20893 26065 20927
rect 26065 20893 26099 20927
rect 26099 20893 26108 20927
rect 26056 20884 26108 20893
rect 26148 20927 26200 20936
rect 26148 20893 26157 20927
rect 26157 20893 26191 20927
rect 26191 20893 26200 20927
rect 26148 20884 26200 20893
rect 26240 20927 26292 20936
rect 26240 20893 26249 20927
rect 26249 20893 26283 20927
rect 26283 20893 26292 20927
rect 26240 20884 26292 20893
rect 26976 20927 27028 20936
rect 26976 20893 26985 20927
rect 26985 20893 27019 20927
rect 27019 20893 27028 20927
rect 26976 20884 27028 20893
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 27620 20884 27672 20936
rect 30472 20884 30524 20936
rect 31024 20884 31076 20936
rect 28724 20816 28776 20868
rect 30564 20816 30616 20868
rect 31392 20927 31444 20936
rect 31392 20893 31401 20927
rect 31401 20893 31435 20927
rect 31435 20893 31444 20927
rect 31392 20884 31444 20893
rect 34336 20884 34388 20936
rect 34796 20884 34848 20936
rect 36636 20927 36688 20936
rect 36636 20893 36645 20927
rect 36645 20893 36679 20927
rect 36679 20893 36688 20927
rect 36636 20884 36688 20893
rect 41236 20927 41288 20936
rect 41236 20893 41270 20927
rect 41270 20893 41288 20927
rect 41236 20884 41288 20893
rect 45192 21131 45244 21140
rect 45192 21097 45201 21131
rect 45201 21097 45235 21131
rect 45235 21097 45244 21131
rect 45192 21088 45244 21097
rect 33600 20816 33652 20868
rect 25320 20748 25372 20800
rect 26792 20791 26844 20800
rect 26792 20757 26801 20791
rect 26801 20757 26835 20791
rect 26835 20757 26844 20791
rect 26792 20748 26844 20757
rect 34980 20791 35032 20800
rect 34980 20757 34989 20791
rect 34989 20757 35023 20791
rect 35023 20757 35032 20791
rect 34980 20748 35032 20757
rect 38016 20791 38068 20800
rect 38016 20757 38025 20791
rect 38025 20757 38059 20791
rect 38059 20757 38068 20791
rect 38016 20748 38068 20757
rect 38660 20816 38712 20868
rect 45836 20927 45888 20936
rect 45836 20893 45845 20927
rect 45845 20893 45879 20927
rect 45879 20893 45888 20927
rect 45836 20884 45888 20893
rect 45928 20816 45980 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 2136 20544 2188 20596
rect 2964 20544 3016 20596
rect 3424 20544 3476 20596
rect 6644 20587 6696 20596
rect 6644 20553 6653 20587
rect 6653 20553 6687 20587
rect 6687 20553 6696 20587
rect 6644 20544 6696 20553
rect 7748 20544 7800 20596
rect 2228 20519 2280 20528
rect 2228 20485 2262 20519
rect 2262 20485 2280 20519
rect 2228 20476 2280 20485
rect 2504 20476 2556 20528
rect 8576 20519 8628 20528
rect 8576 20485 8610 20519
rect 8610 20485 8628 20519
rect 8576 20476 8628 20485
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 11980 20544 12032 20596
rect 12348 20587 12400 20596
rect 12348 20553 12357 20587
rect 12357 20553 12391 20587
rect 12391 20553 12400 20587
rect 12348 20544 12400 20553
rect 13452 20544 13504 20596
rect 11428 20476 11480 20528
rect 1676 20408 1728 20460
rect 940 20340 992 20392
rect 2964 20340 3016 20392
rect 6828 20408 6880 20460
rect 4712 20340 4764 20392
rect 7288 20383 7340 20392
rect 7288 20349 7297 20383
rect 7297 20349 7331 20383
rect 7331 20349 7340 20383
rect 7288 20340 7340 20349
rect 8208 20340 8260 20392
rect 10416 20408 10468 20460
rect 11612 20408 11664 20460
rect 11796 20451 11848 20460
rect 11796 20417 11806 20451
rect 11806 20417 11840 20451
rect 11840 20417 11848 20451
rect 11796 20408 11848 20417
rect 12256 20408 12308 20460
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 14832 20476 14884 20528
rect 12992 20408 13044 20417
rect 13728 20408 13780 20460
rect 26700 20544 26752 20596
rect 27160 20587 27212 20596
rect 27160 20553 27169 20587
rect 27169 20553 27203 20587
rect 27203 20553 27212 20587
rect 27160 20544 27212 20553
rect 28908 20544 28960 20596
rect 33876 20544 33928 20596
rect 37648 20544 37700 20596
rect 38016 20544 38068 20596
rect 44456 20544 44508 20596
rect 17776 20476 17828 20528
rect 20168 20476 20220 20528
rect 12348 20340 12400 20392
rect 2320 20204 2372 20256
rect 3976 20247 4028 20256
rect 3976 20213 3985 20247
rect 3985 20213 4019 20247
rect 4019 20213 4028 20247
rect 3976 20204 4028 20213
rect 6184 20204 6236 20256
rect 6644 20204 6696 20256
rect 6828 20204 6880 20256
rect 8668 20204 8720 20256
rect 10508 20204 10560 20256
rect 11704 20204 11756 20256
rect 12900 20204 12952 20256
rect 18788 20408 18840 20460
rect 19340 20451 19392 20460
rect 19340 20417 19374 20451
rect 19374 20417 19392 20451
rect 19340 20408 19392 20417
rect 18512 20340 18564 20392
rect 20720 20340 20772 20392
rect 26792 20408 26844 20460
rect 27068 20408 27120 20460
rect 28816 20408 28868 20460
rect 26148 20383 26200 20392
rect 26148 20349 26157 20383
rect 26157 20349 26191 20383
rect 26191 20349 26200 20383
rect 26148 20340 26200 20349
rect 26240 20383 26292 20392
rect 26240 20349 26249 20383
rect 26249 20349 26283 20383
rect 26283 20349 26292 20383
rect 26240 20340 26292 20349
rect 26884 20340 26936 20392
rect 27160 20340 27212 20392
rect 27344 20383 27396 20392
rect 27344 20349 27353 20383
rect 27353 20349 27387 20383
rect 27387 20349 27396 20383
rect 27344 20340 27396 20349
rect 27436 20383 27488 20392
rect 27436 20349 27445 20383
rect 27445 20349 27479 20383
rect 27479 20349 27488 20383
rect 27436 20340 27488 20349
rect 27528 20383 27580 20392
rect 27528 20349 27537 20383
rect 27537 20349 27571 20383
rect 27571 20349 27580 20383
rect 27528 20340 27580 20349
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 17684 20272 17736 20324
rect 20168 20272 20220 20324
rect 26332 20272 26384 20324
rect 15292 20204 15344 20256
rect 19432 20204 19484 20256
rect 34520 20476 34572 20528
rect 30012 20408 30064 20460
rect 34704 20408 34756 20460
rect 34796 20408 34848 20460
rect 34980 20408 35032 20460
rect 36544 20408 36596 20460
rect 37096 20408 37148 20460
rect 40224 20476 40276 20528
rect 37740 20451 37792 20460
rect 37740 20417 37774 20451
rect 37774 20417 37792 20451
rect 37740 20408 37792 20417
rect 41420 20408 41472 20460
rect 29920 20340 29972 20392
rect 30196 20340 30248 20392
rect 32036 20340 32088 20392
rect 33784 20340 33836 20392
rect 29828 20204 29880 20256
rect 30012 20204 30064 20256
rect 34428 20204 34480 20256
rect 34704 20204 34756 20256
rect 38108 20204 38160 20256
rect 38844 20247 38896 20256
rect 38844 20213 38853 20247
rect 38853 20213 38887 20247
rect 38887 20213 38896 20247
rect 38844 20204 38896 20213
rect 42064 20247 42116 20256
rect 42064 20213 42073 20247
rect 42073 20213 42107 20247
rect 42107 20213 42116 20247
rect 42064 20204 42116 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6552 20000 6604 20052
rect 10416 20000 10468 20052
rect 10508 20043 10560 20052
rect 10508 20009 10517 20043
rect 10517 20009 10551 20043
rect 10551 20009 10560 20043
rect 10508 20000 10560 20009
rect 7472 19932 7524 19984
rect 940 19864 992 19916
rect 1032 19796 1084 19848
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 940 19728 992 19780
rect 4620 19728 4672 19780
rect 5540 19907 5592 19916
rect 5540 19873 5549 19907
rect 5549 19873 5583 19907
rect 5583 19873 5592 19907
rect 5540 19864 5592 19873
rect 6460 19907 6512 19916
rect 6460 19873 6469 19907
rect 6469 19873 6503 19907
rect 6503 19873 6512 19907
rect 6460 19864 6512 19873
rect 8668 19864 8720 19916
rect 5448 19796 5500 19848
rect 6000 19796 6052 19848
rect 6736 19796 6788 19848
rect 8208 19796 8260 19848
rect 11796 20000 11848 20052
rect 12808 20000 12860 20052
rect 12900 20000 12952 20052
rect 13636 20000 13688 20052
rect 13728 20043 13780 20052
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 16120 20000 16172 20052
rect 19340 20000 19392 20052
rect 23664 20000 23716 20052
rect 24952 20000 25004 20052
rect 28816 20000 28868 20052
rect 37740 20043 37792 20052
rect 37740 20009 37749 20043
rect 37749 20009 37783 20043
rect 37783 20009 37792 20043
rect 37740 20000 37792 20009
rect 41420 20043 41472 20052
rect 41420 20009 41429 20043
rect 41429 20009 41463 20043
rect 41463 20009 41472 20043
rect 41420 20000 41472 20009
rect 11428 19864 11480 19916
rect 11888 19864 11940 19916
rect 13268 19864 13320 19916
rect 11612 19796 11664 19848
rect 13176 19839 13228 19848
rect 13176 19805 13186 19839
rect 13186 19805 13220 19839
rect 13220 19805 13228 19839
rect 13176 19796 13228 19805
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 13636 19864 13688 19916
rect 14832 19796 14884 19848
rect 18052 19864 18104 19916
rect 19248 19796 19300 19848
rect 7840 19728 7892 19780
rect 9128 19771 9180 19780
rect 9128 19737 9137 19771
rect 9137 19737 9171 19771
rect 9171 19737 9180 19771
rect 9128 19728 9180 19737
rect 11152 19728 11204 19780
rect 13360 19771 13412 19780
rect 13360 19737 13369 19771
rect 13369 19737 13403 19771
rect 13403 19737 13412 19771
rect 13360 19728 13412 19737
rect 15108 19771 15160 19780
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 5448 19660 5500 19712
rect 6276 19660 6328 19712
rect 7196 19660 7248 19712
rect 15108 19737 15117 19771
rect 15117 19737 15151 19771
rect 15151 19737 15160 19771
rect 15108 19728 15160 19737
rect 16120 19728 16172 19780
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 20260 19796 20312 19848
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 25136 19932 25188 19984
rect 27528 19932 27580 19984
rect 23572 19864 23624 19916
rect 26700 19864 26752 19916
rect 29368 19864 29420 19916
rect 30932 19907 30984 19916
rect 30932 19873 30941 19907
rect 30941 19873 30975 19907
rect 30975 19873 30984 19907
rect 30932 19864 30984 19873
rect 33508 19864 33560 19916
rect 22284 19728 22336 19780
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 24860 19839 24912 19848
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 24400 19728 24452 19780
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 26056 19796 26108 19848
rect 26240 19839 26292 19848
rect 26240 19805 26249 19839
rect 26249 19805 26283 19839
rect 26283 19805 26292 19839
rect 26240 19796 26292 19805
rect 26332 19839 26384 19848
rect 26332 19805 26341 19839
rect 26341 19805 26375 19839
rect 26375 19805 26384 19839
rect 26332 19796 26384 19805
rect 28724 19796 28776 19848
rect 29920 19796 29972 19848
rect 34520 19796 34572 19848
rect 37464 19932 37516 19984
rect 37096 19907 37148 19916
rect 37096 19873 37105 19907
rect 37105 19873 37139 19907
rect 37139 19873 37148 19907
rect 37096 19864 37148 19873
rect 38844 19932 38896 19984
rect 38660 19864 38712 19916
rect 16488 19703 16540 19712
rect 16488 19669 16497 19703
rect 16497 19669 16531 19703
rect 16531 19669 16540 19703
rect 16488 19660 16540 19669
rect 19432 19660 19484 19712
rect 20904 19703 20956 19712
rect 20904 19669 20913 19703
rect 20913 19669 20947 19703
rect 20947 19669 20956 19703
rect 20904 19660 20956 19669
rect 23480 19703 23532 19712
rect 23480 19669 23489 19703
rect 23489 19669 23523 19703
rect 23523 19669 23532 19703
rect 23480 19660 23532 19669
rect 24308 19660 24360 19712
rect 30012 19728 30064 19780
rect 30104 19728 30156 19780
rect 34796 19728 34848 19780
rect 36360 19771 36412 19780
rect 36360 19737 36369 19771
rect 36369 19737 36403 19771
rect 36403 19737 36412 19771
rect 36360 19728 36412 19737
rect 37464 19796 37516 19848
rect 38016 19839 38068 19848
rect 38016 19805 38025 19839
rect 38025 19805 38059 19839
rect 38059 19805 38068 19839
rect 38016 19796 38068 19805
rect 28908 19660 28960 19712
rect 29184 19660 29236 19712
rect 30288 19660 30340 19712
rect 34336 19703 34388 19712
rect 34336 19669 34345 19703
rect 34345 19669 34379 19703
rect 34379 19669 34388 19703
rect 34336 19660 34388 19669
rect 34888 19660 34940 19712
rect 40408 19796 40460 19848
rect 41604 19839 41656 19848
rect 41604 19805 41613 19839
rect 41613 19805 41647 19839
rect 41647 19805 41656 19839
rect 41604 19796 41656 19805
rect 42064 19796 42116 19848
rect 44180 19796 44232 19848
rect 44456 19796 44508 19848
rect 45560 19839 45612 19848
rect 45560 19805 45569 19839
rect 45569 19805 45603 19839
rect 45603 19805 45612 19839
rect 45560 19796 45612 19805
rect 45652 19839 45704 19848
rect 45652 19805 45661 19839
rect 45661 19805 45695 19839
rect 45695 19805 45704 19839
rect 45652 19796 45704 19805
rect 45836 19839 45888 19848
rect 45836 19805 45845 19839
rect 45845 19805 45879 19839
rect 45879 19805 45888 19839
rect 45836 19796 45888 19805
rect 42892 19728 42944 19780
rect 38568 19660 38620 19712
rect 43352 19660 43404 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 3976 19456 4028 19508
rect 6000 19499 6052 19508
rect 6000 19465 6009 19499
rect 6009 19465 6043 19499
rect 6043 19465 6052 19499
rect 6000 19456 6052 19465
rect 6368 19456 6420 19508
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 12808 19456 12860 19508
rect 16120 19456 16172 19508
rect 16764 19456 16816 19508
rect 20904 19456 20956 19508
rect 24308 19456 24360 19508
rect 24400 19499 24452 19508
rect 24400 19465 24409 19499
rect 24409 19465 24443 19499
rect 24443 19465 24452 19499
rect 24400 19456 24452 19465
rect 26056 19499 26108 19508
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 32496 19456 32548 19508
rect 32588 19499 32640 19508
rect 32588 19465 32597 19499
rect 32597 19465 32631 19499
rect 32631 19465 32640 19499
rect 32588 19456 32640 19465
rect 3240 19388 3292 19440
rect 5540 19388 5592 19440
rect 6184 19388 6236 19440
rect 2688 19252 2740 19304
rect 940 19184 992 19236
rect 6276 19320 6328 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 6736 19388 6788 19440
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 9588 19388 9640 19440
rect 16488 19388 16540 19440
rect 20996 19388 21048 19440
rect 8208 19320 8260 19372
rect 10140 19320 10192 19372
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 23480 19388 23532 19440
rect 25964 19388 26016 19440
rect 27436 19388 27488 19440
rect 4712 19252 4764 19304
rect 6920 19252 6972 19304
rect 2136 19116 2188 19168
rect 5264 19116 5316 19168
rect 9496 19116 9548 19168
rect 22928 19184 22980 19236
rect 27160 19320 27212 19372
rect 25596 19252 25648 19304
rect 24860 19184 24912 19236
rect 25964 19184 26016 19236
rect 26516 19295 26568 19304
rect 26516 19261 26525 19295
rect 26525 19261 26559 19295
rect 26559 19261 26568 19295
rect 26516 19252 26568 19261
rect 28908 19320 28960 19372
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 29368 19363 29420 19372
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 29828 19363 29880 19372
rect 29828 19329 29844 19363
rect 29844 19329 29878 19363
rect 29878 19329 29880 19363
rect 30288 19388 30340 19440
rect 30380 19388 30432 19440
rect 29828 19320 29880 19329
rect 31944 19388 31996 19440
rect 27344 19295 27396 19304
rect 27344 19261 27353 19295
rect 27353 19261 27387 19295
rect 27387 19261 27396 19295
rect 27344 19252 27396 19261
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 27528 19295 27580 19304
rect 27528 19261 27537 19295
rect 27537 19261 27571 19295
rect 27571 19261 27580 19295
rect 27528 19252 27580 19261
rect 27620 19295 27672 19304
rect 27620 19261 27629 19295
rect 27629 19261 27663 19295
rect 27663 19261 27672 19295
rect 27620 19252 27672 19261
rect 31392 19252 31444 19304
rect 32496 19320 32548 19372
rect 32772 19320 32824 19372
rect 34336 19388 34388 19440
rect 27160 19227 27212 19236
rect 27160 19193 27169 19227
rect 27169 19193 27203 19227
rect 27203 19193 27212 19227
rect 27160 19184 27212 19193
rect 23940 19116 23992 19168
rect 26516 19116 26568 19168
rect 31576 19184 31628 19236
rect 33508 19184 33560 19236
rect 34520 19320 34572 19372
rect 34704 19320 34756 19372
rect 34336 19252 34388 19304
rect 35440 19320 35492 19372
rect 36268 19363 36320 19372
rect 36268 19329 36277 19363
rect 36277 19329 36311 19363
rect 36311 19329 36320 19363
rect 36268 19320 36320 19329
rect 37372 19388 37424 19440
rect 38476 19388 38528 19440
rect 37280 19320 37332 19372
rect 37648 19363 37700 19372
rect 37648 19329 37655 19363
rect 37655 19329 37700 19363
rect 37648 19320 37700 19329
rect 38016 19320 38068 19372
rect 38108 19320 38160 19372
rect 42432 19388 42484 19440
rect 34612 19184 34664 19236
rect 36176 19184 36228 19236
rect 37280 19184 37332 19236
rect 27528 19116 27580 19168
rect 31208 19159 31260 19168
rect 31208 19125 31217 19159
rect 31217 19125 31251 19159
rect 31251 19125 31260 19159
rect 31208 19116 31260 19125
rect 37096 19116 37148 19168
rect 37464 19116 37516 19168
rect 41604 19320 41656 19372
rect 45652 19456 45704 19508
rect 43352 19363 43404 19372
rect 43352 19329 43361 19363
rect 43361 19329 43395 19363
rect 43395 19329 43404 19363
rect 43352 19320 43404 19329
rect 43904 19363 43956 19372
rect 43904 19329 43913 19363
rect 43913 19329 43947 19363
rect 43947 19329 43956 19363
rect 43904 19320 43956 19329
rect 44180 19320 44232 19372
rect 45560 19388 45612 19440
rect 42892 19295 42944 19304
rect 42892 19261 42901 19295
rect 42901 19261 42935 19295
rect 42935 19261 42944 19295
rect 42892 19252 42944 19261
rect 44456 19252 44508 19304
rect 45928 19184 45980 19236
rect 40960 19159 41012 19168
rect 40960 19125 40969 19159
rect 40969 19125 41003 19159
rect 41003 19125 41012 19159
rect 40960 19116 41012 19125
rect 42800 19116 42852 19168
rect 43904 19116 43956 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3240 18955 3292 18964
rect 3240 18921 3249 18955
rect 3249 18921 3283 18955
rect 3283 18921 3292 18955
rect 3240 18912 3292 18921
rect 4068 18912 4120 18964
rect 6736 18912 6788 18964
rect 9588 18912 9640 18964
rect 9956 18912 10008 18964
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 11704 18912 11756 18964
rect 12440 18912 12492 18964
rect 13360 18955 13412 18964
rect 13360 18921 13369 18955
rect 13369 18921 13403 18955
rect 13403 18921 13412 18955
rect 13360 18912 13412 18921
rect 22376 18912 22428 18964
rect 26148 18912 26200 18964
rect 9772 18844 9824 18896
rect 6828 18776 6880 18828
rect 1768 18708 1820 18760
rect 2136 18751 2188 18760
rect 2136 18717 2170 18751
rect 2170 18717 2188 18751
rect 2136 18708 2188 18717
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 6368 18708 6420 18760
rect 5908 18640 5960 18692
rect 7932 18708 7984 18760
rect 20168 18844 20220 18896
rect 11428 18776 11480 18828
rect 22284 18844 22336 18896
rect 22652 18844 22704 18896
rect 26424 18887 26476 18896
rect 26424 18853 26433 18887
rect 26433 18853 26467 18887
rect 26467 18853 26476 18887
rect 26424 18844 26476 18853
rect 9956 18751 10008 18760
rect 9956 18717 9970 18751
rect 9970 18717 10004 18751
rect 10004 18717 10008 18751
rect 9956 18708 10008 18717
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 11888 18708 11940 18760
rect 16396 18708 16448 18760
rect 9864 18683 9916 18692
rect 9864 18649 9873 18683
rect 9873 18649 9907 18683
rect 9907 18649 9916 18683
rect 9864 18640 9916 18649
rect 11704 18683 11756 18692
rect 11704 18649 11713 18683
rect 11713 18649 11747 18683
rect 11747 18649 11756 18683
rect 11704 18640 11756 18649
rect 12164 18572 12216 18624
rect 12900 18640 12952 18692
rect 19340 18572 19392 18624
rect 23664 18776 23716 18828
rect 24768 18776 24820 18828
rect 25596 18776 25648 18828
rect 26976 18844 27028 18896
rect 27344 18844 27396 18896
rect 31392 18955 31444 18964
rect 31392 18921 31401 18955
rect 31401 18921 31435 18955
rect 31435 18921 31444 18955
rect 31392 18912 31444 18921
rect 32588 18912 32640 18964
rect 27160 18776 27212 18828
rect 30104 18776 30156 18828
rect 42432 18887 42484 18896
rect 42432 18853 42441 18887
rect 42441 18853 42475 18887
rect 42475 18853 42484 18887
rect 42432 18844 42484 18853
rect 42800 18844 42852 18896
rect 20076 18708 20128 18760
rect 20904 18708 20956 18760
rect 20996 18708 21048 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 19984 18640 20036 18692
rect 21732 18708 21784 18760
rect 22836 18751 22888 18760
rect 22836 18717 22845 18751
rect 22845 18717 22879 18751
rect 22879 18717 22888 18751
rect 22836 18708 22888 18717
rect 23296 18708 23348 18760
rect 24860 18708 24912 18760
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 20720 18572 20772 18624
rect 21456 18572 21508 18624
rect 24768 18640 24820 18692
rect 26332 18640 26384 18692
rect 26884 18751 26936 18760
rect 26884 18717 26893 18751
rect 26893 18717 26927 18751
rect 26927 18717 26936 18751
rect 26884 18708 26936 18717
rect 28724 18708 28776 18760
rect 31024 18708 31076 18760
rect 31116 18708 31168 18760
rect 31576 18751 31628 18760
rect 31576 18717 31585 18751
rect 31585 18717 31619 18751
rect 31619 18717 31628 18751
rect 31576 18708 31628 18717
rect 32588 18708 32640 18760
rect 36360 18751 36412 18760
rect 36360 18717 36369 18751
rect 36369 18717 36403 18751
rect 36403 18717 36412 18751
rect 36360 18708 36412 18717
rect 37464 18708 37516 18760
rect 37648 18708 37700 18760
rect 41328 18776 41380 18828
rect 30104 18640 30156 18692
rect 30380 18640 30432 18692
rect 31208 18640 31260 18692
rect 32036 18683 32088 18692
rect 32036 18649 32045 18683
rect 32045 18649 32079 18683
rect 32079 18649 32088 18683
rect 32036 18640 32088 18649
rect 34796 18640 34848 18692
rect 36544 18640 36596 18692
rect 40316 18640 40368 18692
rect 40960 18708 41012 18760
rect 42156 18640 42208 18692
rect 25872 18572 25924 18624
rect 40592 18572 40644 18624
rect 41604 18615 41656 18624
rect 41604 18581 41613 18615
rect 41613 18581 41647 18615
rect 41647 18581 41656 18615
rect 41604 18572 41656 18581
rect 42340 18708 42392 18760
rect 44456 18955 44508 18964
rect 44456 18921 44465 18955
rect 44465 18921 44499 18955
rect 44499 18921 44508 18955
rect 44456 18912 44508 18921
rect 43904 18844 43956 18896
rect 44180 18776 44232 18828
rect 45928 18819 45980 18828
rect 45928 18785 45937 18819
rect 45937 18785 45971 18819
rect 45971 18785 45980 18819
rect 45928 18776 45980 18785
rect 44180 18640 44232 18692
rect 44272 18683 44324 18692
rect 44272 18649 44281 18683
rect 44281 18649 44315 18683
rect 44315 18649 44324 18683
rect 44272 18640 44324 18649
rect 45560 18683 45612 18692
rect 45560 18649 45569 18683
rect 45569 18649 45603 18683
rect 45603 18649 45612 18683
rect 45560 18640 45612 18649
rect 43720 18572 43772 18624
rect 43812 18572 43864 18624
rect 45744 18572 45796 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 1032 18368 1084 18420
rect 940 18300 992 18352
rect 2780 18368 2832 18420
rect 11704 18368 11756 18420
rect 19984 18368 20036 18420
rect 3424 18300 3476 18352
rect 21456 18300 21508 18352
rect 14740 18232 14792 18284
rect 15016 18164 15068 18216
rect 16672 18164 16724 18216
rect 16856 18164 16908 18216
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17132 18232 17184 18284
rect 19432 18232 19484 18284
rect 2780 18139 2832 18148
rect 2780 18105 2789 18139
rect 2789 18105 2823 18139
rect 2823 18105 2832 18139
rect 2780 18096 2832 18105
rect 9772 18096 9824 18148
rect 17224 18096 17276 18148
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 17960 18164 18012 18216
rect 22192 18368 22244 18420
rect 22928 18368 22980 18420
rect 25044 18368 25096 18420
rect 25872 18368 25924 18420
rect 26516 18368 26568 18420
rect 26700 18368 26752 18420
rect 40500 18368 40552 18420
rect 40592 18411 40644 18420
rect 40592 18377 40601 18411
rect 40601 18377 40635 18411
rect 40635 18377 40644 18411
rect 40592 18368 40644 18377
rect 42156 18368 42208 18420
rect 44456 18368 44508 18420
rect 23940 18300 23992 18352
rect 22100 18232 22152 18284
rect 24860 18275 24912 18284
rect 24860 18241 24869 18275
rect 24869 18241 24903 18275
rect 24903 18241 24912 18275
rect 24860 18232 24912 18241
rect 24952 18232 25004 18284
rect 25688 18275 25740 18284
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 30472 18232 30524 18284
rect 30656 18275 30708 18284
rect 30656 18241 30690 18275
rect 30690 18241 30708 18275
rect 30656 18232 30708 18241
rect 31024 18232 31076 18284
rect 31576 18232 31628 18284
rect 24768 18207 24820 18216
rect 24768 18173 24777 18207
rect 24777 18173 24811 18207
rect 24811 18173 24820 18207
rect 24768 18164 24820 18173
rect 25596 18207 25648 18216
rect 25596 18173 25605 18207
rect 25605 18173 25639 18207
rect 25639 18173 25648 18207
rect 25596 18164 25648 18173
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 30380 18207 30432 18216
rect 30380 18173 30389 18207
rect 30389 18173 30423 18207
rect 30423 18173 30432 18207
rect 30380 18164 30432 18173
rect 32680 18300 32732 18352
rect 37280 18300 37332 18352
rect 32772 18232 32824 18284
rect 37464 18275 37516 18284
rect 37464 18241 37473 18275
rect 37473 18241 37507 18275
rect 37507 18241 37516 18275
rect 37464 18232 37516 18241
rect 37648 18275 37700 18284
rect 37648 18241 37657 18275
rect 37657 18241 37691 18275
rect 37691 18241 37700 18275
rect 37648 18232 37700 18241
rect 41236 18300 41288 18352
rect 43076 18300 43128 18352
rect 34152 18164 34204 18216
rect 36452 18164 36504 18216
rect 26884 18096 26936 18148
rect 31392 18096 31444 18148
rect 20720 18028 20772 18080
rect 22008 18028 22060 18080
rect 23664 18028 23716 18080
rect 24768 18028 24820 18080
rect 31300 18028 31352 18080
rect 31852 18028 31904 18080
rect 38108 18096 38160 18148
rect 40224 18275 40276 18284
rect 40224 18241 40233 18275
rect 40233 18241 40267 18275
rect 40267 18241 40276 18275
rect 40224 18232 40276 18241
rect 40592 18232 40644 18284
rect 41328 18232 41380 18284
rect 41512 18232 41564 18284
rect 42064 18164 42116 18216
rect 43260 18275 43312 18284
rect 43260 18241 43269 18275
rect 43269 18241 43303 18275
rect 43303 18241 43312 18275
rect 43260 18232 43312 18241
rect 43444 18275 43496 18284
rect 43444 18241 43451 18275
rect 43451 18241 43496 18275
rect 43444 18232 43496 18241
rect 43536 18275 43588 18284
rect 43536 18241 43545 18275
rect 43545 18241 43579 18275
rect 43579 18241 43588 18275
rect 43536 18232 43588 18241
rect 43720 18275 43772 18284
rect 43720 18241 43734 18275
rect 43734 18241 43768 18275
rect 43768 18241 43772 18275
rect 43720 18232 43772 18241
rect 45560 18300 45612 18352
rect 40040 18096 40092 18148
rect 43260 18096 43312 18148
rect 37280 18028 37332 18080
rect 38660 18028 38712 18080
rect 41512 18028 41564 18080
rect 41604 18028 41656 18080
rect 44272 18164 44324 18216
rect 44180 18096 44232 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1768 17688 1820 17740
rect 5172 17824 5224 17876
rect 5356 17867 5408 17876
rect 5356 17833 5365 17867
rect 5365 17833 5399 17867
rect 5399 17833 5408 17867
rect 5356 17824 5408 17833
rect 17132 17824 17184 17876
rect 19432 17867 19484 17876
rect 19432 17833 19441 17867
rect 19441 17833 19475 17867
rect 19475 17833 19484 17867
rect 19432 17824 19484 17833
rect 22100 17824 22152 17876
rect 22836 17824 22888 17876
rect 27620 17824 27672 17876
rect 30656 17867 30708 17876
rect 30656 17833 30665 17867
rect 30665 17833 30699 17867
rect 30699 17833 30708 17867
rect 30656 17824 30708 17833
rect 940 17620 992 17672
rect 1124 17552 1176 17604
rect 8484 17756 8536 17808
rect 19524 17756 19576 17808
rect 28080 17756 28132 17808
rect 15292 17688 15344 17740
rect 5172 17620 5224 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 8208 17620 8260 17672
rect 12992 17620 13044 17672
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 14648 17663 14700 17672
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 17960 17620 18012 17672
rect 4988 17552 5040 17604
rect 8944 17552 8996 17604
rect 11704 17552 11756 17604
rect 16856 17552 16908 17604
rect 17224 17552 17276 17604
rect 19340 17620 19392 17672
rect 23388 17688 23440 17740
rect 30472 17688 30524 17740
rect 31300 17688 31352 17740
rect 20076 17620 20128 17672
rect 21824 17663 21876 17672
rect 21824 17629 21833 17663
rect 21833 17629 21867 17663
rect 21867 17629 21876 17663
rect 21824 17620 21876 17629
rect 22008 17663 22060 17672
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 22192 17620 22244 17672
rect 27528 17620 27580 17672
rect 37924 17824 37976 17876
rect 40500 17824 40552 17876
rect 38016 17756 38068 17808
rect 40592 17756 40644 17808
rect 36544 17731 36596 17740
rect 36544 17697 36553 17731
rect 36553 17697 36587 17731
rect 36587 17697 36596 17731
rect 36544 17688 36596 17697
rect 19984 17552 20036 17604
rect 26240 17552 26292 17604
rect 30656 17552 30708 17604
rect 35532 17620 35584 17672
rect 35624 17663 35676 17672
rect 35624 17629 35633 17663
rect 35633 17629 35667 17663
rect 35667 17629 35676 17663
rect 35624 17620 35676 17629
rect 35808 17663 35860 17672
rect 35808 17629 35817 17663
rect 35817 17629 35851 17663
rect 35851 17629 35860 17663
rect 35808 17620 35860 17629
rect 37280 17620 37332 17672
rect 40040 17663 40092 17672
rect 40040 17629 40049 17663
rect 40049 17629 40083 17663
rect 40083 17629 40092 17663
rect 40040 17620 40092 17629
rect 41604 17688 41656 17740
rect 40592 17620 40644 17672
rect 31116 17552 31168 17604
rect 32036 17552 32088 17604
rect 33876 17552 33928 17604
rect 36360 17552 36412 17604
rect 37372 17552 37424 17604
rect 2412 17484 2464 17536
rect 11336 17484 11388 17536
rect 11980 17484 12032 17536
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 17408 17484 17460 17536
rect 20260 17484 20312 17536
rect 21916 17484 21968 17536
rect 23572 17484 23624 17536
rect 25228 17484 25280 17536
rect 34428 17484 34480 17536
rect 34612 17484 34664 17536
rect 36084 17484 36136 17536
rect 37188 17484 37240 17536
rect 37280 17484 37332 17536
rect 40224 17484 40276 17536
rect 40500 17484 40552 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 3424 17280 3476 17332
rect 4528 17280 4580 17332
rect 4712 17280 4764 17332
rect 4988 17323 5040 17332
rect 4988 17289 4997 17323
rect 4997 17289 5031 17323
rect 5031 17289 5040 17323
rect 4988 17280 5040 17289
rect 7288 17280 7340 17332
rect 8944 17323 8996 17332
rect 8944 17289 8953 17323
rect 8953 17289 8987 17323
rect 8987 17289 8996 17323
rect 8944 17280 8996 17289
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 940 17212 992 17264
rect 5632 17212 5684 17264
rect 8024 17212 8076 17264
rect 8484 17212 8536 17264
rect 4528 17187 4580 17196
rect 4528 17153 4535 17187
rect 4535 17153 4580 17187
rect 4528 17144 4580 17153
rect 2688 17076 2740 17128
rect 3240 17008 3292 17060
rect 5356 17076 5408 17128
rect 5908 17008 5960 17060
rect 2044 16940 2096 16992
rect 2412 16940 2464 16992
rect 2688 16940 2740 16992
rect 6644 16940 6696 16992
rect 6736 16940 6788 16992
rect 7288 17144 7340 17196
rect 9588 17144 9640 17196
rect 11980 17212 12032 17264
rect 14280 17212 14332 17264
rect 17040 17280 17092 17332
rect 17316 17280 17368 17332
rect 18512 17280 18564 17332
rect 11612 17076 11664 17128
rect 9680 17008 9732 17060
rect 10324 17008 10376 17060
rect 14740 17144 14792 17196
rect 15844 17144 15896 17196
rect 16396 17144 16448 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 17500 17144 17552 17196
rect 17960 17187 18012 17196
rect 17960 17153 17969 17187
rect 17969 17153 18003 17187
rect 18003 17153 18012 17187
rect 17960 17144 18012 17153
rect 18236 17187 18288 17196
rect 18236 17153 18270 17187
rect 18270 17153 18288 17187
rect 18236 17144 18288 17153
rect 23572 17144 23624 17196
rect 33692 17280 33744 17332
rect 33876 17323 33928 17332
rect 33876 17289 33885 17323
rect 33885 17289 33919 17323
rect 33919 17289 33928 17323
rect 33876 17280 33928 17289
rect 34152 17280 34204 17332
rect 37464 17323 37516 17332
rect 37464 17289 37473 17323
rect 37473 17289 37507 17323
rect 37507 17289 37516 17323
rect 37464 17280 37516 17289
rect 43536 17280 43588 17332
rect 45744 17323 45796 17332
rect 45744 17289 45753 17323
rect 45753 17289 45787 17323
rect 45787 17289 45796 17323
rect 45744 17280 45796 17289
rect 45928 17280 45980 17332
rect 46388 17280 46440 17332
rect 23940 17212 23992 17264
rect 24124 17144 24176 17196
rect 30380 17212 30432 17264
rect 34428 17255 34480 17264
rect 34428 17221 34437 17255
rect 34437 17221 34471 17255
rect 34471 17221 34480 17255
rect 34428 17212 34480 17221
rect 34796 17212 34848 17264
rect 27436 17187 27488 17196
rect 27436 17153 27470 17187
rect 27470 17153 27488 17187
rect 27436 17144 27488 17153
rect 29184 17144 29236 17196
rect 29460 17187 29512 17196
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 30288 17144 30340 17196
rect 32312 17187 32364 17196
rect 32312 17153 32321 17187
rect 32321 17153 32355 17187
rect 32355 17153 32364 17187
rect 32312 17144 32364 17153
rect 32680 17144 32732 17196
rect 12992 17119 13044 17128
rect 12992 17085 13001 17119
rect 13001 17085 13035 17119
rect 13035 17085 13044 17119
rect 12992 17076 13044 17085
rect 17132 17119 17184 17128
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 17132 17076 17184 17085
rect 14648 17008 14700 17060
rect 17868 17008 17920 17060
rect 23664 17008 23716 17060
rect 24216 17076 24268 17128
rect 24584 17076 24636 17128
rect 24676 17076 24728 17128
rect 24860 17119 24912 17128
rect 24860 17085 24869 17119
rect 24869 17085 24903 17119
rect 24903 17085 24912 17119
rect 24860 17076 24912 17085
rect 9588 16940 9640 16992
rect 16580 16940 16632 16992
rect 18972 16940 19024 16992
rect 23480 16940 23532 16992
rect 28172 17076 28224 17128
rect 30472 17076 30524 17128
rect 30656 17076 30708 17128
rect 32588 17051 32640 17060
rect 32588 17017 32597 17051
rect 32597 17017 32631 17051
rect 32631 17017 32640 17051
rect 32588 17008 32640 17017
rect 33508 17144 33560 17196
rect 35992 17212 36044 17264
rect 35900 17144 35952 17196
rect 36084 17187 36136 17196
rect 36084 17153 36093 17187
rect 36093 17153 36127 17187
rect 36127 17153 36136 17187
rect 36084 17144 36136 17153
rect 37280 17212 37332 17264
rect 36360 17187 36412 17196
rect 36360 17153 36369 17187
rect 36369 17153 36403 17187
rect 36403 17153 36412 17187
rect 36360 17144 36412 17153
rect 35532 17076 35584 17128
rect 36636 17144 36688 17196
rect 38016 17212 38068 17264
rect 40224 17212 40276 17264
rect 43904 17212 43956 17264
rect 44456 17212 44508 17264
rect 37556 17144 37608 17196
rect 37924 17187 37976 17196
rect 37924 17153 37933 17187
rect 37933 17153 37967 17187
rect 37967 17153 37976 17187
rect 37924 17144 37976 17153
rect 43536 17144 43588 17196
rect 43812 17187 43864 17196
rect 43812 17153 43822 17187
rect 43822 17153 43856 17187
rect 43856 17153 43864 17187
rect 44180 17187 44232 17196
rect 43812 17144 43864 17153
rect 44180 17153 44194 17187
rect 44194 17153 44228 17187
rect 44228 17153 44232 17187
rect 44180 17144 44232 17153
rect 45652 17187 45704 17196
rect 45652 17153 45661 17187
rect 45661 17153 45695 17187
rect 45695 17153 45704 17187
rect 45652 17144 45704 17153
rect 36912 17076 36964 17128
rect 38660 17076 38712 17128
rect 45744 17076 45796 17128
rect 46112 17076 46164 17128
rect 27896 16940 27948 16992
rect 28908 16940 28960 16992
rect 33324 16940 33376 16992
rect 35624 16940 35676 16992
rect 35900 16940 35952 16992
rect 36360 16940 36412 16992
rect 36544 17008 36596 17060
rect 37188 17008 37240 17060
rect 37832 17051 37884 17060
rect 37832 17017 37841 17051
rect 37841 17017 37875 17051
rect 37875 17017 37884 17051
rect 37832 17008 37884 17017
rect 45468 17051 45520 17060
rect 45468 17017 45477 17051
rect 45477 17017 45511 17051
rect 45511 17017 45520 17051
rect 45468 17008 45520 17017
rect 45836 17008 45888 17060
rect 45284 16940 45336 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7012 16736 7064 16788
rect 10508 16736 10560 16788
rect 14464 16736 14516 16788
rect 24032 16736 24084 16788
rect 24768 16736 24820 16788
rect 24952 16736 25004 16788
rect 6184 16668 6236 16720
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 5172 16600 5224 16652
rect 15200 16600 15252 16652
rect 15384 16600 15436 16652
rect 20720 16668 20772 16720
rect 21364 16668 21416 16720
rect 27436 16736 27488 16788
rect 28908 16779 28960 16788
rect 28908 16745 28917 16779
rect 28917 16745 28951 16779
rect 28951 16745 28960 16779
rect 28908 16736 28960 16745
rect 940 16532 992 16584
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 5632 16575 5684 16584
rect 5632 16541 5641 16575
rect 5641 16541 5675 16575
rect 5675 16541 5684 16575
rect 5632 16532 5684 16541
rect 5816 16575 5868 16584
rect 5816 16541 5823 16575
rect 5823 16541 5868 16575
rect 5816 16532 5868 16541
rect 5908 16575 5960 16584
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 6000 16575 6052 16584
rect 6000 16541 6009 16575
rect 6009 16541 6043 16575
rect 6043 16541 6052 16575
rect 6000 16532 6052 16541
rect 6644 16532 6696 16584
rect 7012 16575 7064 16584
rect 7012 16541 7046 16575
rect 7046 16541 7064 16575
rect 7012 16532 7064 16541
rect 9772 16532 9824 16584
rect 11796 16532 11848 16584
rect 14556 16532 14608 16584
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 16580 16575 16632 16584
rect 16580 16541 16590 16575
rect 16590 16541 16624 16575
rect 16624 16541 16632 16575
rect 16580 16532 16632 16541
rect 17040 16600 17092 16652
rect 17316 16600 17368 16652
rect 19432 16600 19484 16652
rect 23480 16643 23532 16652
rect 23480 16609 23489 16643
rect 23489 16609 23523 16643
rect 23523 16609 23532 16643
rect 23480 16600 23532 16609
rect 24952 16600 25004 16652
rect 25320 16643 25372 16652
rect 25320 16609 25329 16643
rect 25329 16609 25363 16643
rect 25363 16609 25372 16643
rect 25320 16600 25372 16609
rect 6828 16464 6880 16516
rect 17684 16532 17736 16584
rect 17040 16464 17092 16516
rect 21180 16532 21232 16584
rect 23664 16575 23716 16584
rect 23664 16541 23673 16575
rect 23673 16541 23707 16575
rect 23707 16541 23716 16575
rect 23664 16532 23716 16541
rect 20812 16464 20864 16516
rect 22192 16464 22244 16516
rect 23296 16464 23348 16516
rect 24216 16532 24268 16584
rect 24676 16532 24728 16584
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 23848 16464 23900 16516
rect 24768 16464 24820 16516
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 28172 16668 28224 16720
rect 27528 16643 27580 16652
rect 27528 16609 27537 16643
rect 27537 16609 27571 16643
rect 27571 16609 27580 16643
rect 27528 16600 27580 16609
rect 29092 16643 29144 16652
rect 29092 16609 29101 16643
rect 29101 16609 29135 16643
rect 29135 16609 29144 16643
rect 29092 16600 29144 16609
rect 30380 16736 30432 16788
rect 31300 16736 31352 16788
rect 32588 16736 32640 16788
rect 35900 16736 35952 16788
rect 37832 16736 37884 16788
rect 43812 16736 43864 16788
rect 34152 16668 34204 16720
rect 36728 16668 36780 16720
rect 43720 16668 43772 16720
rect 27896 16575 27948 16584
rect 27896 16541 27905 16575
rect 27905 16541 27939 16575
rect 27939 16541 27948 16575
rect 27896 16532 27948 16541
rect 11520 16396 11572 16448
rect 11704 16396 11756 16448
rect 16304 16396 16356 16448
rect 17132 16396 17184 16448
rect 17408 16396 17460 16448
rect 20076 16396 20128 16448
rect 21364 16396 21416 16448
rect 23572 16396 23624 16448
rect 27528 16396 27580 16448
rect 29184 16532 29236 16584
rect 33324 16600 33376 16652
rect 37280 16643 37332 16652
rect 34612 16532 34664 16584
rect 37280 16609 37289 16643
rect 37289 16609 37323 16643
rect 37323 16609 37332 16643
rect 37280 16600 37332 16609
rect 38660 16600 38712 16652
rect 40316 16643 40368 16652
rect 40316 16609 40325 16643
rect 40325 16609 40359 16643
rect 40359 16609 40368 16643
rect 40316 16600 40368 16609
rect 45744 16600 45796 16652
rect 34520 16464 34572 16516
rect 30748 16396 30800 16448
rect 34796 16396 34848 16448
rect 43812 16532 43864 16584
rect 45652 16532 45704 16584
rect 46112 16575 46164 16584
rect 46112 16541 46121 16575
rect 46121 16541 46155 16575
rect 46155 16541 46164 16575
rect 46112 16532 46164 16541
rect 46388 16575 46440 16584
rect 46388 16541 46397 16575
rect 46397 16541 46431 16575
rect 46431 16541 46440 16575
rect 46388 16532 46440 16541
rect 36728 16464 36780 16516
rect 37648 16507 37700 16516
rect 37648 16473 37657 16507
rect 37657 16473 37691 16507
rect 37691 16473 37700 16507
rect 37648 16464 37700 16473
rect 40040 16464 40092 16516
rect 45560 16464 45612 16516
rect 37280 16396 37332 16448
rect 37464 16439 37516 16448
rect 37464 16405 37473 16439
rect 37473 16405 37507 16439
rect 37507 16405 37516 16439
rect 37464 16396 37516 16405
rect 38844 16396 38896 16448
rect 43628 16396 43680 16448
rect 45468 16396 45520 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2780 16192 2832 16244
rect 5816 16192 5868 16244
rect 940 16124 992 16176
rect 11520 16124 11572 16176
rect 4068 16056 4120 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7196 16056 7248 16108
rect 7748 16056 7800 16108
rect 2596 15988 2648 16040
rect 6736 16031 6788 16040
rect 6736 15997 6745 16031
rect 6745 15997 6779 16031
rect 6779 15997 6788 16031
rect 6736 15988 6788 15997
rect 2964 15895 3016 15904
rect 2964 15861 2973 15895
rect 2973 15861 3007 15895
rect 3007 15861 3016 15895
rect 2964 15852 3016 15861
rect 8024 15852 8076 15904
rect 9312 15852 9364 15904
rect 14188 16192 14240 16244
rect 14648 16192 14700 16244
rect 16304 16235 16356 16244
rect 16304 16201 16313 16235
rect 16313 16201 16347 16235
rect 16347 16201 16356 16235
rect 16304 16192 16356 16201
rect 18236 16192 18288 16244
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 25136 16192 25188 16244
rect 31024 16192 31076 16244
rect 33692 16192 33744 16244
rect 37280 16192 37332 16244
rect 40040 16235 40092 16244
rect 40040 16201 40049 16235
rect 40049 16201 40083 16235
rect 40083 16201 40092 16235
rect 40040 16192 40092 16201
rect 40408 16235 40460 16244
rect 40408 16201 40417 16235
rect 40417 16201 40451 16235
rect 40451 16201 40460 16235
rect 40408 16192 40460 16201
rect 12992 16124 13044 16176
rect 15200 16167 15252 16176
rect 14832 16056 14884 16108
rect 15200 16133 15234 16167
rect 15234 16133 15252 16167
rect 15200 16124 15252 16133
rect 17592 16124 17644 16176
rect 18880 16124 18932 16176
rect 18972 16124 19024 16176
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 18052 15988 18104 16040
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 20996 16124 21048 16176
rect 25044 16124 25096 16176
rect 25596 16124 25648 16176
rect 29184 16124 29236 16176
rect 30472 16124 30524 16176
rect 33784 16124 33836 16176
rect 18052 15852 18104 15904
rect 18788 15852 18840 15904
rect 19800 16031 19852 16040
rect 19800 15997 19809 16031
rect 19809 15997 19843 16031
rect 19843 15997 19852 16031
rect 19800 15988 19852 15997
rect 20260 15988 20312 16040
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 21272 16056 21324 16108
rect 21732 16056 21784 16108
rect 22100 16056 22152 16108
rect 24492 16099 24544 16108
rect 24492 16065 24501 16099
rect 24501 16065 24535 16099
rect 24535 16065 24544 16099
rect 24492 16056 24544 16065
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 25688 16056 25740 16108
rect 26148 16099 26200 16108
rect 26148 16065 26157 16099
rect 26157 16065 26191 16099
rect 26191 16065 26200 16099
rect 26148 16056 26200 16065
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 29920 16056 29972 16108
rect 20720 15852 20772 15904
rect 21088 15988 21140 16040
rect 30748 16099 30800 16108
rect 30748 16065 30757 16099
rect 30757 16065 30791 16099
rect 30791 16065 30800 16099
rect 30748 16056 30800 16065
rect 33140 16056 33192 16108
rect 33876 16099 33928 16108
rect 33876 16065 33885 16099
rect 33885 16065 33919 16099
rect 33919 16065 33928 16099
rect 33876 16056 33928 16065
rect 37464 16167 37516 16176
rect 37464 16133 37473 16167
rect 37473 16133 37507 16167
rect 37507 16133 37516 16167
rect 37464 16124 37516 16133
rect 37648 16167 37700 16176
rect 34060 16056 34112 16108
rect 34244 16099 34296 16108
rect 34244 16065 34253 16099
rect 34253 16065 34287 16099
rect 34287 16065 34296 16099
rect 34244 16056 34296 16065
rect 34520 16056 34572 16108
rect 36728 16056 36780 16108
rect 37648 16133 37673 16167
rect 37673 16133 37700 16167
rect 37648 16124 37700 16133
rect 40224 16099 40276 16108
rect 40224 16065 40233 16099
rect 40233 16065 40267 16099
rect 40267 16065 40276 16099
rect 40224 16056 40276 16065
rect 43720 16124 43772 16176
rect 43536 16099 43588 16108
rect 43536 16065 43545 16099
rect 43545 16065 43579 16099
rect 43579 16065 43588 16099
rect 43536 16056 43588 16065
rect 43628 16099 43680 16108
rect 43628 16065 43638 16099
rect 43638 16065 43672 16099
rect 43672 16065 43680 16099
rect 43628 16056 43680 16065
rect 43812 16099 43864 16108
rect 43812 16065 43821 16099
rect 43821 16065 43855 16099
rect 43855 16065 43864 16099
rect 43812 16056 43864 16065
rect 44916 16192 44968 16244
rect 45560 16235 45612 16244
rect 45560 16201 45569 16235
rect 45569 16201 45603 16235
rect 45603 16201 45612 16235
rect 45560 16192 45612 16201
rect 43996 16099 44048 16108
rect 43996 16065 44010 16099
rect 44010 16065 44044 16099
rect 44044 16065 44048 16099
rect 43996 16056 44048 16065
rect 38108 15988 38160 16040
rect 45744 16031 45796 16040
rect 45744 15997 45753 16031
rect 45753 15997 45787 16031
rect 45787 15997 45796 16031
rect 45744 15988 45796 15997
rect 45836 16031 45888 16040
rect 45836 15997 45845 16031
rect 45845 15997 45879 16031
rect 45879 15997 45888 16031
rect 45836 15988 45888 15997
rect 36268 15920 36320 15972
rect 36728 15920 36780 15972
rect 22008 15852 22060 15904
rect 24676 15852 24728 15904
rect 30196 15852 30248 15904
rect 33876 15852 33928 15904
rect 36084 15852 36136 15904
rect 36820 15852 36872 15904
rect 44180 15963 44232 15972
rect 44180 15929 44189 15963
rect 44189 15929 44223 15963
rect 44223 15929 44232 15963
rect 44180 15920 44232 15929
rect 42984 15852 43036 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 7748 15648 7800 15700
rect 11704 15648 11756 15700
rect 11888 15648 11940 15700
rect 5632 15580 5684 15632
rect 7932 15580 7984 15632
rect 14832 15648 14884 15700
rect 17500 15648 17552 15700
rect 21088 15648 21140 15700
rect 22100 15691 22152 15700
rect 22100 15657 22109 15691
rect 22109 15657 22143 15691
rect 22143 15657 22152 15691
rect 22100 15648 22152 15657
rect 23388 15648 23440 15700
rect 6184 15512 6236 15564
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 14096 15444 14148 15496
rect 17040 15580 17092 15632
rect 27804 15580 27856 15632
rect 29092 15648 29144 15700
rect 32404 15648 32456 15700
rect 33048 15648 33100 15700
rect 33784 15648 33836 15700
rect 34152 15648 34204 15700
rect 34520 15648 34572 15700
rect 31024 15580 31076 15632
rect 40224 15648 40276 15700
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 14740 15487 14792 15496
rect 14740 15453 14754 15487
rect 14754 15453 14788 15487
rect 14788 15453 14792 15487
rect 17500 15555 17552 15564
rect 17500 15521 17509 15555
rect 17509 15521 17543 15555
rect 17543 15521 17552 15555
rect 17500 15512 17552 15521
rect 19800 15512 19852 15564
rect 21180 15512 21232 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 22008 15512 22060 15564
rect 14740 15444 14792 15453
rect 19064 15444 19116 15496
rect 940 15376 992 15428
rect 1032 15308 1084 15360
rect 5540 15376 5592 15428
rect 12440 15376 12492 15428
rect 12808 15376 12860 15428
rect 19432 15376 19484 15428
rect 22100 15444 22152 15496
rect 22192 15444 22244 15496
rect 21272 15376 21324 15428
rect 22744 15419 22796 15428
rect 22744 15385 22753 15419
rect 22753 15385 22787 15419
rect 22787 15385 22796 15419
rect 22744 15376 22796 15385
rect 26332 15444 26384 15496
rect 24676 15376 24728 15428
rect 24952 15376 25004 15428
rect 27528 15512 27580 15564
rect 26700 15444 26752 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 30748 15512 30800 15564
rect 36728 15580 36780 15632
rect 36820 15623 36872 15632
rect 36820 15589 36829 15623
rect 36829 15589 36863 15623
rect 36863 15589 36872 15623
rect 36820 15580 36872 15589
rect 37280 15580 37332 15632
rect 30196 15487 30248 15496
rect 30196 15453 30205 15487
rect 30205 15453 30239 15487
rect 30239 15453 30248 15487
rect 30196 15444 30248 15453
rect 27528 15376 27580 15428
rect 28080 15376 28132 15428
rect 33140 15444 33192 15496
rect 40316 15512 40368 15564
rect 33692 15487 33744 15496
rect 33692 15453 33706 15487
rect 33706 15453 33740 15487
rect 33740 15453 33744 15487
rect 33692 15444 33744 15453
rect 34152 15444 34204 15496
rect 36728 15487 36780 15496
rect 36728 15453 36737 15487
rect 36737 15453 36771 15487
rect 36771 15453 36780 15487
rect 36728 15444 36780 15453
rect 33416 15376 33468 15428
rect 9312 15308 9364 15360
rect 11520 15308 11572 15360
rect 19984 15308 20036 15360
rect 27712 15308 27764 15360
rect 34704 15376 34756 15428
rect 35992 15376 36044 15428
rect 36636 15376 36688 15428
rect 42616 15376 42668 15428
rect 34060 15308 34112 15360
rect 35900 15308 35952 15360
rect 36728 15308 36780 15360
rect 37556 15308 37608 15360
rect 43812 15308 43864 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 11244 15104 11296 15156
rect 19432 15104 19484 15156
rect 1124 15036 1176 15088
rect 2964 15079 3016 15088
rect 2964 15045 2998 15079
rect 2998 15045 3016 15079
rect 2964 15036 3016 15045
rect 7104 15011 7156 15020
rect 7104 14977 7138 15011
rect 7138 14977 7156 15011
rect 7104 14968 7156 14977
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 3976 14764 4028 14816
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 4896 14764 4948 14816
rect 8300 14764 8352 14816
rect 9220 14764 9272 14816
rect 11704 15036 11756 15088
rect 12348 15036 12400 15088
rect 11796 14968 11848 15020
rect 18604 14968 18656 15020
rect 19892 15079 19944 15088
rect 19892 15045 19901 15079
rect 19901 15045 19935 15079
rect 19935 15045 19944 15079
rect 19892 15036 19944 15045
rect 20720 15104 20772 15156
rect 22100 15036 22152 15088
rect 24124 15036 24176 15088
rect 28080 15079 28132 15088
rect 28080 15045 28089 15079
rect 28089 15045 28123 15079
rect 28123 15045 28132 15079
rect 28080 15036 28132 15045
rect 15016 14900 15068 14952
rect 17500 14900 17552 14952
rect 21272 14968 21324 15020
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 24768 14968 24820 15020
rect 25504 14968 25556 15020
rect 23020 14943 23072 14952
rect 23020 14909 23029 14943
rect 23029 14909 23063 14943
rect 23063 14909 23072 14943
rect 23020 14900 23072 14909
rect 11336 14832 11388 14884
rect 22928 14832 22980 14884
rect 23296 14943 23348 14952
rect 23296 14909 23305 14943
rect 23305 14909 23339 14943
rect 23339 14909 23348 14943
rect 23296 14900 23348 14909
rect 12256 14764 12308 14816
rect 13452 14764 13504 14816
rect 23848 14764 23900 14816
rect 25320 14875 25372 14884
rect 25320 14841 25329 14875
rect 25329 14841 25363 14875
rect 25363 14841 25372 14875
rect 25320 14832 25372 14841
rect 26424 15011 26476 15020
rect 26424 14977 26438 15011
rect 26438 14977 26472 15011
rect 26472 14977 26476 15011
rect 26424 14968 26476 14977
rect 27804 15011 27856 15020
rect 27804 14977 27813 15011
rect 27813 14977 27847 15011
rect 27847 14977 27856 15011
rect 27804 14968 27856 14977
rect 29000 14968 29052 15020
rect 29920 14968 29972 15020
rect 27344 14900 27396 14952
rect 27620 14900 27672 14952
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 31300 14968 31352 15020
rect 33048 15036 33100 15088
rect 28632 14832 28684 14884
rect 27620 14764 27672 14816
rect 30196 14764 30248 14816
rect 33324 14764 33376 14816
rect 35808 15011 35860 15020
rect 35808 14977 35817 15011
rect 35817 14977 35851 15011
rect 35851 14977 35860 15011
rect 35808 14968 35860 14977
rect 34520 14900 34572 14952
rect 38844 15147 38896 15156
rect 38844 15113 38853 15147
rect 38853 15113 38887 15147
rect 38887 15113 38896 15147
rect 38844 15104 38896 15113
rect 42616 15147 42668 15156
rect 42616 15113 42625 15147
rect 42625 15113 42659 15147
rect 42659 15113 42668 15147
rect 42616 15104 42668 15113
rect 42984 15147 43036 15156
rect 42984 15113 42993 15147
rect 42993 15113 43027 15147
rect 43027 15113 43036 15147
rect 42984 15104 43036 15113
rect 43812 15104 43864 15156
rect 37188 14968 37240 15020
rect 36452 14900 36504 14952
rect 43904 15036 43956 15088
rect 43720 15011 43772 15020
rect 43720 14977 43729 15011
rect 43729 14977 43763 15011
rect 43763 14977 43772 15011
rect 43720 14968 43772 14977
rect 43812 15011 43864 15020
rect 43812 14977 43822 15011
rect 43822 14977 43856 15011
rect 43856 14977 43864 15011
rect 43812 14968 43864 14977
rect 44088 15011 44140 15020
rect 44088 14977 44097 15011
rect 44097 14977 44131 15011
rect 44131 14977 44140 15011
rect 44088 14968 44140 14977
rect 44180 15011 44232 15020
rect 44180 14977 44194 15011
rect 44194 14977 44228 15011
rect 44228 14977 44232 15011
rect 44180 14968 44232 14977
rect 45284 14900 45336 14952
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 7104 14560 7156 14612
rect 11796 14603 11848 14612
rect 11796 14569 11805 14603
rect 11805 14569 11839 14603
rect 11839 14569 11848 14603
rect 11796 14560 11848 14569
rect 11980 14560 12032 14612
rect 33784 14560 33836 14612
rect 36636 14603 36688 14612
rect 36636 14569 36645 14603
rect 36645 14569 36679 14603
rect 36679 14569 36688 14603
rect 36636 14560 36688 14569
rect 37004 14560 37056 14612
rect 40316 14560 40368 14612
rect 11244 14492 11296 14544
rect 16212 14492 16264 14544
rect 17500 14492 17552 14544
rect 18604 14492 18656 14544
rect 24676 14535 24728 14544
rect 24676 14501 24685 14535
rect 24685 14501 24719 14535
rect 24719 14501 24728 14535
rect 24676 14492 24728 14501
rect 24768 14535 24820 14544
rect 24768 14501 24777 14535
rect 24777 14501 24811 14535
rect 24811 14501 24820 14535
rect 24768 14492 24820 14501
rect 26240 14492 26292 14544
rect 26700 14535 26752 14544
rect 26700 14501 26709 14535
rect 26709 14501 26743 14535
rect 26743 14501 26752 14535
rect 26700 14492 26752 14501
rect 940 14424 992 14476
rect 2504 14356 2556 14408
rect 3976 14467 4028 14476
rect 3976 14433 3985 14467
rect 3985 14433 4019 14467
rect 4019 14433 4028 14467
rect 3976 14424 4028 14433
rect 6828 14424 6880 14476
rect 7380 14424 7432 14476
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 4068 14356 4120 14408
rect 5540 14356 5592 14408
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 11336 14399 11388 14408
rect 11336 14365 11343 14399
rect 11343 14365 11388 14399
rect 11336 14356 11388 14365
rect 940 14288 992 14340
rect 3792 14288 3844 14340
rect 5632 14331 5684 14340
rect 5632 14297 5641 14331
rect 5641 14297 5675 14331
rect 5675 14297 5684 14331
rect 5632 14288 5684 14297
rect 8208 14288 8260 14340
rect 10784 14288 10836 14340
rect 12808 14356 12860 14408
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 28632 14492 28684 14544
rect 33416 14492 33468 14544
rect 14924 14356 14976 14408
rect 17500 14356 17552 14408
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 24952 14356 25004 14408
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 26240 14356 26292 14408
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 27712 14424 27764 14476
rect 29000 14424 29052 14476
rect 31392 14424 31444 14476
rect 40224 14492 40276 14544
rect 26608 14356 26660 14365
rect 8300 14220 8352 14272
rect 11152 14220 11204 14272
rect 12164 14220 12216 14272
rect 12256 14220 12308 14272
rect 13636 14288 13688 14340
rect 16304 14288 16356 14340
rect 16488 14331 16540 14340
rect 16488 14297 16522 14331
rect 16522 14297 16540 14331
rect 16488 14288 16540 14297
rect 16580 14288 16632 14340
rect 15108 14220 15160 14272
rect 21916 14288 21968 14340
rect 30104 14356 30156 14408
rect 30564 14356 30616 14408
rect 30748 14356 30800 14408
rect 35624 14356 35676 14408
rect 37004 14356 37056 14408
rect 38844 14356 38896 14408
rect 27528 14331 27580 14340
rect 27528 14297 27537 14331
rect 27537 14297 27571 14331
rect 27571 14297 27580 14331
rect 27528 14288 27580 14297
rect 25320 14220 25372 14272
rect 26608 14220 26660 14272
rect 27252 14220 27304 14272
rect 27896 14331 27948 14340
rect 27896 14297 27905 14331
rect 27905 14297 27939 14331
rect 27939 14297 27948 14331
rect 27896 14288 27948 14297
rect 29828 14288 29880 14340
rect 34520 14288 34572 14340
rect 40040 14288 40092 14340
rect 40132 14331 40184 14340
rect 40132 14297 40141 14331
rect 40141 14297 40175 14331
rect 40175 14297 40184 14331
rect 40132 14288 40184 14297
rect 27712 14263 27764 14272
rect 27712 14229 27721 14263
rect 27721 14229 27755 14263
rect 27755 14229 27764 14263
rect 27712 14220 27764 14229
rect 28816 14220 28868 14272
rect 30472 14220 30524 14272
rect 30564 14263 30616 14272
rect 30564 14229 30573 14263
rect 30573 14229 30607 14263
rect 30607 14229 30616 14263
rect 30564 14220 30616 14229
rect 34244 14220 34296 14272
rect 35808 14220 35860 14272
rect 36728 14220 36780 14272
rect 44180 14288 44232 14340
rect 40316 14263 40368 14272
rect 40316 14229 40325 14263
rect 40325 14229 40359 14263
rect 40359 14229 40368 14263
rect 40316 14220 40368 14229
rect 41604 14220 41656 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 5632 14016 5684 14068
rect 10600 14016 10652 14068
rect 12992 14016 13044 14068
rect 14096 14016 14148 14068
rect 14832 14016 14884 14068
rect 16488 14016 16540 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 21824 14016 21876 14068
rect 23020 14016 23072 14068
rect 27528 14016 27580 14068
rect 30196 14016 30248 14068
rect 30748 14059 30800 14068
rect 30748 14025 30757 14059
rect 30757 14025 30791 14059
rect 30791 14025 30800 14059
rect 30748 14016 30800 14025
rect 33784 14059 33836 14068
rect 33784 14025 33793 14059
rect 33793 14025 33827 14059
rect 33827 14025 33836 14059
rect 33784 14016 33836 14025
rect 3976 13948 4028 14000
rect 10232 13948 10284 14000
rect 1952 13923 2004 13932
rect 1952 13889 1986 13923
rect 1986 13889 2004 13923
rect 1952 13880 2004 13889
rect 4804 13880 4856 13932
rect 9128 13880 9180 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 12348 13948 12400 14000
rect 2596 13676 2648 13728
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 6828 13812 6880 13864
rect 11612 13812 11664 13864
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 13636 13880 13688 13932
rect 16580 13948 16632 14000
rect 14464 13880 14516 13932
rect 16212 13880 16264 13932
rect 18144 13948 18196 14000
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 18604 13880 18656 13932
rect 23756 13948 23808 14000
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 21548 13880 21600 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 23664 13880 23716 13932
rect 23940 13923 23992 13932
rect 23940 13889 23949 13923
rect 23949 13889 23983 13923
rect 23983 13889 23992 13923
rect 23940 13880 23992 13889
rect 24860 13880 24912 13932
rect 30288 13948 30340 14000
rect 33416 13991 33468 14000
rect 33416 13957 33425 13991
rect 33425 13957 33459 13991
rect 33459 13957 33468 13991
rect 33416 13948 33468 13957
rect 37740 13991 37792 14000
rect 37740 13957 37749 13991
rect 37749 13957 37783 13991
rect 37783 13957 37792 13991
rect 37740 13948 37792 13957
rect 29920 13880 29972 13932
rect 33140 13923 33192 13932
rect 20628 13812 20680 13864
rect 21088 13855 21140 13864
rect 21088 13821 21097 13855
rect 21097 13821 21131 13855
rect 21131 13821 21140 13855
rect 21088 13812 21140 13821
rect 23296 13812 23348 13864
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 4988 13744 5040 13796
rect 7656 13676 7708 13728
rect 12164 13744 12216 13796
rect 9404 13719 9456 13728
rect 9404 13685 9413 13719
rect 9413 13685 9447 13719
rect 9447 13685 9456 13719
rect 9404 13676 9456 13685
rect 12072 13676 12124 13728
rect 29000 13744 29052 13796
rect 17868 13676 17920 13728
rect 22468 13676 22520 13728
rect 28264 13676 28316 13728
rect 33140 13889 33149 13923
rect 33149 13889 33183 13923
rect 33183 13889 33192 13923
rect 33140 13880 33192 13889
rect 33324 13923 33376 13932
rect 33324 13889 33331 13923
rect 33331 13889 33376 13923
rect 33324 13880 33376 13889
rect 33508 13923 33560 13932
rect 33508 13889 33517 13923
rect 33517 13889 33551 13923
rect 33551 13889 33560 13923
rect 33508 13880 33560 13889
rect 33600 13923 33652 13932
rect 33600 13889 33614 13923
rect 33614 13889 33648 13923
rect 33648 13889 33652 13923
rect 33600 13880 33652 13889
rect 37464 13923 37516 13932
rect 37464 13889 37473 13923
rect 37473 13889 37507 13923
rect 37507 13889 37516 13923
rect 37464 13880 37516 13889
rect 37648 13923 37700 13932
rect 37648 13889 37657 13923
rect 37657 13889 37691 13923
rect 37691 13889 37700 13923
rect 37648 13880 37700 13889
rect 38108 14016 38160 14068
rect 40776 13948 40828 14000
rect 30472 13812 30524 13864
rect 36728 13812 36780 13864
rect 32036 13744 32088 13796
rect 32864 13744 32916 13796
rect 38936 13812 38988 13864
rect 31484 13676 31536 13728
rect 35992 13676 36044 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 2504 13472 2556 13524
rect 4988 13472 5040 13524
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 11888 13472 11940 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 8208 13404 8260 13456
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 7656 13336 7708 13388
rect 15384 13404 15436 13456
rect 12900 13336 12952 13388
rect 13176 13336 13228 13388
rect 16580 13404 16632 13456
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 16948 13472 17000 13524
rect 19156 13472 19208 13524
rect 21088 13472 21140 13524
rect 26700 13472 26752 13524
rect 26976 13472 27028 13524
rect 29920 13515 29972 13524
rect 29920 13481 29929 13515
rect 29929 13481 29963 13515
rect 29963 13481 29972 13515
rect 29920 13472 29972 13481
rect 30564 13472 30616 13524
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5908 13268 5960 13320
rect 6828 13268 6880 13320
rect 9036 13268 9088 13320
rect 10140 13268 10192 13320
rect 12348 13311 12400 13320
rect 12348 13277 12357 13311
rect 12357 13277 12391 13311
rect 12391 13277 12400 13311
rect 12348 13268 12400 13277
rect 16856 13336 16908 13388
rect 22560 13336 22612 13388
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 16672 13268 16724 13320
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 20812 13268 20864 13320
rect 21732 13268 21784 13320
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 22928 13404 22980 13456
rect 53104 13472 53156 13524
rect 29000 13336 29052 13388
rect 30196 13336 30248 13388
rect 34612 13404 34664 13456
rect 940 13200 992 13252
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 6368 13200 6420 13252
rect 12900 13200 12952 13252
rect 3056 13132 3108 13184
rect 3332 13175 3384 13184
rect 3332 13141 3341 13175
rect 3341 13141 3375 13175
rect 3375 13141 3384 13175
rect 3332 13132 3384 13141
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 9404 13132 9456 13184
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 10968 13132 11020 13184
rect 18512 13200 18564 13252
rect 18880 13175 18932 13184
rect 18880 13141 18889 13175
rect 18889 13141 18923 13175
rect 18923 13141 18932 13175
rect 18880 13132 18932 13141
rect 20996 13200 21048 13252
rect 23664 13268 23716 13320
rect 27252 13311 27304 13320
rect 27252 13277 27261 13311
rect 27261 13277 27295 13311
rect 27295 13277 27304 13311
rect 27252 13268 27304 13277
rect 27896 13268 27948 13320
rect 30748 13268 30800 13320
rect 32036 13311 32088 13320
rect 32036 13277 32045 13311
rect 32045 13277 32079 13311
rect 32079 13277 32088 13311
rect 32036 13268 32088 13277
rect 37464 13404 37516 13456
rect 37280 13336 37332 13388
rect 35992 13311 36044 13320
rect 35992 13277 36001 13311
rect 36001 13277 36035 13311
rect 36035 13277 36044 13311
rect 35992 13268 36044 13277
rect 23756 13200 23808 13252
rect 27988 13200 28040 13252
rect 31852 13243 31904 13252
rect 31852 13209 31861 13243
rect 31861 13209 31895 13243
rect 31895 13209 31904 13243
rect 31852 13200 31904 13209
rect 32496 13200 32548 13252
rect 35900 13243 35952 13252
rect 35900 13209 35909 13243
rect 35909 13209 35943 13243
rect 35943 13209 35952 13243
rect 35900 13200 35952 13209
rect 37096 13311 37148 13320
rect 37096 13277 37105 13311
rect 37105 13277 37139 13311
rect 37139 13277 37148 13311
rect 37096 13268 37148 13277
rect 40776 13268 40828 13320
rect 41328 13268 41380 13320
rect 41604 13268 41656 13320
rect 37556 13200 37608 13252
rect 27436 13132 27488 13184
rect 31576 13132 31628 13184
rect 36268 13175 36320 13184
rect 36268 13141 36277 13175
rect 36277 13141 36311 13175
rect 36311 13141 36320 13175
rect 36268 13132 36320 13141
rect 39856 13132 39908 13184
rect 43812 13132 43864 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 940 12928 992 12980
rect 4068 12928 4120 12980
rect 8944 12928 8996 12980
rect 1032 12860 1084 12912
rect 9588 12860 9640 12912
rect 6368 12792 6420 12844
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 10876 12928 10928 12980
rect 10416 12792 10468 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 11980 12835 12032 12844
rect 11980 12801 12014 12835
rect 12014 12801 12032 12835
rect 11980 12792 12032 12801
rect 12348 12928 12400 12980
rect 16672 12928 16724 12980
rect 16856 12928 16908 12980
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 18604 12928 18656 12980
rect 12164 12860 12216 12912
rect 18880 12903 18932 12912
rect 18880 12869 18889 12903
rect 18889 12869 18923 12903
rect 18923 12869 18932 12903
rect 18880 12860 18932 12869
rect 940 12724 992 12776
rect 3332 12724 3384 12776
rect 3056 12656 3108 12708
rect 8944 12656 8996 12708
rect 9312 12724 9364 12776
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 17224 12792 17276 12844
rect 21732 12928 21784 12980
rect 23940 12928 23992 12980
rect 24860 12971 24912 12980
rect 24860 12937 24869 12971
rect 24869 12937 24903 12971
rect 24903 12937 24912 12971
rect 24860 12928 24912 12937
rect 22100 12860 22152 12912
rect 22652 12860 22704 12912
rect 26424 12928 26476 12980
rect 27436 12928 27488 12980
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 19432 12724 19484 12776
rect 24584 12792 24636 12844
rect 25780 12792 25832 12844
rect 22560 12767 22612 12776
rect 22560 12733 22569 12767
rect 22569 12733 22603 12767
rect 22603 12733 22612 12767
rect 22560 12724 22612 12733
rect 22744 12724 22796 12776
rect 23480 12767 23532 12776
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 26332 12903 26384 12912
rect 26332 12869 26341 12903
rect 26341 12869 26375 12903
rect 26375 12869 26384 12903
rect 26332 12860 26384 12869
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 31852 12928 31904 12980
rect 34060 12928 34112 12980
rect 37280 12928 37332 12980
rect 37648 12928 37700 12980
rect 38108 12928 38160 12980
rect 40040 12928 40092 12980
rect 40776 12928 40828 12980
rect 43720 12860 43772 12912
rect 28264 12835 28316 12844
rect 28264 12801 28273 12835
rect 28273 12801 28307 12835
rect 28307 12801 28316 12835
rect 28264 12792 28316 12801
rect 28816 12792 28868 12844
rect 31576 12835 31628 12844
rect 31576 12801 31585 12835
rect 31585 12801 31619 12835
rect 31619 12801 31628 12835
rect 31576 12792 31628 12801
rect 33140 12835 33192 12844
rect 33140 12801 33149 12835
rect 33149 12801 33183 12835
rect 33183 12801 33192 12835
rect 33140 12792 33192 12801
rect 34244 12792 34296 12844
rect 35624 12835 35676 12844
rect 35624 12801 35658 12835
rect 35658 12801 35676 12835
rect 35624 12792 35676 12801
rect 39856 12792 39908 12844
rect 40040 12792 40092 12844
rect 40776 12792 40828 12844
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 9404 12588 9456 12640
rect 15292 12588 15344 12640
rect 16028 12588 16080 12640
rect 21364 12588 21416 12640
rect 22100 12588 22152 12640
rect 25044 12656 25096 12708
rect 26884 12656 26936 12708
rect 28816 12656 28868 12708
rect 31300 12724 31352 12776
rect 34060 12724 34112 12776
rect 35348 12767 35400 12776
rect 35348 12733 35357 12767
rect 35357 12733 35391 12767
rect 35391 12733 35400 12767
rect 35348 12724 35400 12733
rect 37280 12724 37332 12776
rect 38292 12724 38344 12776
rect 33600 12656 33652 12708
rect 26792 12588 26844 12640
rect 31852 12588 31904 12640
rect 34244 12588 34296 12640
rect 36728 12631 36780 12640
rect 36728 12597 36737 12631
rect 36737 12597 36771 12631
rect 36771 12597 36780 12631
rect 36728 12588 36780 12597
rect 41420 12588 41472 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3792 12384 3844 12436
rect 7380 12316 7432 12368
rect 2780 12248 2832 12300
rect 940 12180 992 12232
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 1032 12112 1084 12164
rect 3884 12112 3936 12164
rect 2688 12044 2740 12096
rect 3424 12044 3476 12096
rect 7288 12180 7340 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 8116 12180 8168 12232
rect 10048 12112 10100 12164
rect 10324 12155 10376 12164
rect 4344 12044 4396 12096
rect 4988 12044 5040 12096
rect 10324 12121 10333 12155
rect 10333 12121 10367 12155
rect 10367 12121 10376 12155
rect 10324 12112 10376 12121
rect 11980 12384 12032 12436
rect 13268 12384 13320 12436
rect 11612 12248 11664 12300
rect 16856 12384 16908 12436
rect 15476 12316 15528 12368
rect 22560 12384 22612 12436
rect 24584 12427 24636 12436
rect 24584 12393 24593 12427
rect 24593 12393 24627 12427
rect 24627 12393 24636 12427
rect 24584 12384 24636 12393
rect 27252 12316 27304 12368
rect 27896 12427 27948 12436
rect 27896 12393 27905 12427
rect 27905 12393 27939 12427
rect 27939 12393 27948 12427
rect 27896 12384 27948 12393
rect 27988 12384 28040 12436
rect 31208 12384 31260 12436
rect 35624 12384 35676 12436
rect 35900 12384 35952 12436
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 16488 12248 16540 12300
rect 11060 12180 11112 12232
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 14188 12180 14240 12232
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 15568 12112 15620 12164
rect 16580 12180 16632 12232
rect 16764 12180 16816 12232
rect 17776 12248 17828 12300
rect 20168 12112 20220 12164
rect 20352 12155 20404 12164
rect 20352 12121 20361 12155
rect 20361 12121 20395 12155
rect 20395 12121 20404 12155
rect 20352 12112 20404 12121
rect 21364 12223 21416 12232
rect 21364 12189 21398 12223
rect 21398 12189 21416 12223
rect 21364 12180 21416 12189
rect 23848 12180 23900 12232
rect 21640 12112 21692 12164
rect 24860 12180 24912 12232
rect 25044 12223 25096 12232
rect 25044 12189 25053 12223
rect 25053 12189 25087 12223
rect 25087 12189 25096 12223
rect 25044 12180 25096 12189
rect 25228 12112 25280 12164
rect 26332 12248 26384 12300
rect 27160 12248 27212 12300
rect 35992 12316 36044 12368
rect 31208 12248 31260 12300
rect 38108 12316 38160 12368
rect 26700 12223 26752 12232
rect 26700 12189 26709 12223
rect 26709 12189 26743 12223
rect 26743 12189 26752 12223
rect 26700 12180 26752 12189
rect 26792 12223 26844 12232
rect 26792 12189 26801 12223
rect 26801 12189 26835 12223
rect 26835 12189 26844 12223
rect 26792 12180 26844 12189
rect 26976 12223 27028 12232
rect 26976 12189 26985 12223
rect 26985 12189 27019 12223
rect 27019 12189 27028 12223
rect 26976 12180 27028 12189
rect 27344 12180 27396 12232
rect 28356 12223 28408 12232
rect 28356 12189 28365 12223
rect 28365 12189 28399 12223
rect 28399 12189 28408 12223
rect 28356 12180 28408 12189
rect 28448 12223 28500 12232
rect 28448 12189 28458 12223
rect 28458 12189 28492 12223
rect 28492 12189 28500 12223
rect 28448 12180 28500 12189
rect 28816 12223 28868 12232
rect 28816 12189 28830 12223
rect 28830 12189 28864 12223
rect 28864 12189 28868 12223
rect 28816 12180 28868 12189
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 31852 12180 31904 12232
rect 32496 12180 32548 12232
rect 37188 12291 37240 12300
rect 37188 12257 37197 12291
rect 37197 12257 37231 12291
rect 37231 12257 37240 12291
rect 37188 12248 37240 12257
rect 38752 12248 38804 12300
rect 44088 12316 44140 12368
rect 47952 12316 48004 12368
rect 10692 12044 10744 12096
rect 12348 12044 12400 12096
rect 15384 12044 15436 12096
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 16672 12044 16724 12096
rect 18420 12044 18472 12096
rect 19064 12044 19116 12096
rect 25964 12087 26016 12096
rect 25964 12053 25973 12087
rect 25973 12053 26007 12087
rect 26007 12053 26016 12087
rect 25964 12044 26016 12053
rect 28540 12112 28592 12164
rect 28632 12155 28684 12164
rect 28632 12121 28641 12155
rect 28641 12121 28675 12155
rect 28675 12121 28684 12155
rect 28632 12112 28684 12121
rect 28724 12155 28776 12164
rect 28724 12121 28733 12155
rect 28733 12121 28767 12155
rect 28767 12121 28776 12155
rect 28724 12112 28776 12121
rect 28908 12112 28960 12164
rect 30012 12044 30064 12096
rect 30656 12112 30708 12164
rect 36268 12180 36320 12232
rect 36728 12180 36780 12232
rect 38660 12223 38712 12232
rect 35532 12112 35584 12164
rect 38660 12189 38669 12223
rect 38669 12189 38703 12223
rect 38703 12189 38712 12223
rect 38660 12180 38712 12189
rect 39028 12223 39080 12232
rect 39028 12189 39037 12223
rect 39037 12189 39071 12223
rect 39071 12189 39080 12223
rect 39028 12180 39080 12189
rect 39212 12180 39264 12232
rect 33140 12087 33192 12096
rect 33140 12053 33149 12087
rect 33149 12053 33183 12087
rect 33183 12053 33192 12087
rect 33140 12044 33192 12053
rect 38936 12155 38988 12164
rect 38936 12121 38945 12155
rect 38945 12121 38979 12155
rect 38979 12121 38988 12155
rect 38936 12112 38988 12121
rect 41328 12223 41380 12232
rect 41328 12189 41337 12223
rect 41337 12189 41371 12223
rect 41371 12189 41380 12223
rect 41328 12180 41380 12189
rect 41420 12180 41472 12232
rect 42340 12112 42392 12164
rect 40224 12044 40276 12096
rect 40408 12087 40460 12096
rect 40408 12053 40417 12087
rect 40417 12053 40451 12087
rect 40451 12053 40460 12087
rect 40408 12044 40460 12053
rect 42432 12044 42484 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 3424 11883 3476 11892
rect 3424 11849 3433 11883
rect 3433 11849 3467 11883
rect 3467 11849 3476 11883
rect 3424 11840 3476 11849
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 1124 11772 1176 11824
rect 2780 11815 2832 11824
rect 2780 11781 2789 11815
rect 2789 11781 2823 11815
rect 2823 11781 2832 11815
rect 2780 11772 2832 11781
rect 3056 11772 3108 11824
rect 3700 11704 3752 11756
rect 4252 11704 4304 11756
rect 5356 11772 5408 11824
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 12072 11840 12124 11892
rect 15476 11840 15528 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 16580 11840 16632 11892
rect 17224 11883 17276 11892
rect 17224 11849 17233 11883
rect 17233 11849 17267 11883
rect 17267 11849 17276 11883
rect 17224 11840 17276 11849
rect 17500 11840 17552 11892
rect 17776 11840 17828 11892
rect 18144 11840 18196 11892
rect 940 11636 992 11688
rect 2504 11636 2556 11688
rect 2228 11500 2280 11552
rect 8024 11704 8076 11756
rect 8760 11772 8812 11824
rect 14188 11772 14240 11824
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 7380 11636 7432 11688
rect 7840 11636 7892 11688
rect 10508 11704 10560 11756
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 16488 11772 16540 11824
rect 16764 11704 16816 11756
rect 17868 11747 17920 11756
rect 17868 11713 17877 11747
rect 17877 11713 17911 11747
rect 17911 11713 17920 11747
rect 17868 11704 17920 11713
rect 20352 11840 20404 11892
rect 20628 11840 20680 11892
rect 21640 11840 21692 11892
rect 22284 11840 22336 11892
rect 25964 11840 26016 11892
rect 28448 11840 28500 11892
rect 29368 11840 29420 11892
rect 30012 11840 30064 11892
rect 20168 11815 20220 11824
rect 20168 11781 20177 11815
rect 20177 11781 20211 11815
rect 20211 11781 20220 11815
rect 20168 11772 20220 11781
rect 24492 11772 24544 11824
rect 25596 11772 25648 11824
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 14188 11636 14240 11688
rect 21364 11636 21416 11688
rect 5540 11568 5592 11620
rect 10324 11568 10376 11620
rect 20996 11568 21048 11620
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 30288 11772 30340 11824
rect 39028 11772 39080 11824
rect 39856 11815 39908 11824
rect 39856 11781 39865 11815
rect 39865 11781 39899 11815
rect 39899 11781 39908 11815
rect 39856 11772 39908 11781
rect 40132 11883 40184 11892
rect 40132 11849 40141 11883
rect 40141 11849 40175 11883
rect 40175 11849 40184 11883
rect 40132 11840 40184 11849
rect 55956 11772 56008 11824
rect 27252 11704 27304 11756
rect 28540 11704 28592 11756
rect 29000 11704 29052 11756
rect 29460 11704 29512 11756
rect 29736 11747 29788 11756
rect 29736 11713 29745 11747
rect 29745 11713 29779 11747
rect 29779 11713 29788 11747
rect 29736 11704 29788 11713
rect 32864 11704 32916 11756
rect 33324 11704 33376 11756
rect 38568 11747 38620 11756
rect 38568 11713 38577 11747
rect 38577 11713 38611 11747
rect 38611 11713 38620 11747
rect 38568 11704 38620 11713
rect 21640 11636 21692 11688
rect 25688 11679 25740 11688
rect 25688 11645 25697 11679
rect 25697 11645 25731 11679
rect 25731 11645 25740 11679
rect 25688 11636 25740 11645
rect 7472 11500 7524 11552
rect 8116 11543 8168 11552
rect 8116 11509 8125 11543
rect 8125 11509 8159 11543
rect 8159 11509 8168 11543
rect 8116 11500 8168 11509
rect 9496 11500 9548 11552
rect 16672 11500 16724 11552
rect 18604 11500 18656 11552
rect 19984 11500 20036 11552
rect 21548 11568 21600 11620
rect 25596 11568 25648 11620
rect 25964 11679 26016 11688
rect 25964 11645 25973 11679
rect 25973 11645 26007 11679
rect 26007 11645 26016 11679
rect 25964 11636 26016 11645
rect 27160 11679 27212 11688
rect 27160 11645 27169 11679
rect 27169 11645 27203 11679
rect 27203 11645 27212 11679
rect 27160 11636 27212 11645
rect 30380 11636 30432 11688
rect 38844 11747 38896 11756
rect 38844 11713 38853 11747
rect 38853 11713 38887 11747
rect 38887 11713 38896 11747
rect 38844 11704 38896 11713
rect 39120 11636 39172 11688
rect 39948 11747 40000 11756
rect 39948 11713 39957 11747
rect 39957 11713 39991 11747
rect 39991 11713 40000 11747
rect 39948 11704 40000 11713
rect 42432 11636 42484 11688
rect 40040 11568 40092 11620
rect 28080 11500 28132 11552
rect 31484 11500 31536 11552
rect 37924 11500 37976 11552
rect 38660 11500 38712 11552
rect 43260 11500 43312 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4988 11339 5040 11348
rect 4988 11305 4997 11339
rect 4997 11305 5031 11339
rect 5031 11305 5040 11339
rect 4988 11296 5040 11305
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 3056 11271 3108 11280
rect 3056 11237 3065 11271
rect 3065 11237 3099 11271
rect 3099 11237 3108 11271
rect 3056 11228 3108 11237
rect 3700 11228 3752 11280
rect 6460 11228 6512 11280
rect 3884 11160 3936 11212
rect 5356 11160 5408 11212
rect 8300 11296 8352 11348
rect 12900 11296 12952 11348
rect 16304 11296 16356 11348
rect 17868 11296 17920 11348
rect 19340 11296 19392 11348
rect 21364 11296 21416 11348
rect 23664 11296 23716 11348
rect 27712 11296 27764 11348
rect 28632 11296 28684 11348
rect 29736 11296 29788 11348
rect 38568 11296 38620 11348
rect 8392 11228 8444 11280
rect 8760 11160 8812 11212
rect 10140 11228 10192 11280
rect 9496 11160 9548 11212
rect 24676 11228 24728 11280
rect 3976 11092 4028 11144
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7288 11092 7340 11144
rect 1952 11067 2004 11076
rect 1952 11033 1986 11067
rect 1986 11033 2004 11067
rect 1952 11024 2004 11033
rect 5264 11024 5316 11076
rect 7932 11092 7984 11144
rect 8024 11092 8076 11144
rect 7564 11024 7616 11076
rect 9956 11092 10008 11144
rect 10968 11160 11020 11212
rect 13820 11160 13872 11212
rect 16580 11160 16632 11212
rect 10508 11092 10560 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 9864 11024 9916 11076
rect 14188 11092 14240 11144
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15108 11092 15160 11144
rect 12256 11024 12308 11076
rect 15016 11024 15068 11076
rect 16212 11135 16264 11144
rect 16212 11101 16221 11135
rect 16221 11101 16255 11135
rect 16255 11101 16264 11135
rect 16212 11092 16264 11101
rect 17132 11092 17184 11144
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 30012 11160 30064 11212
rect 33968 11228 34020 11280
rect 38936 11228 38988 11280
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 18052 11024 18104 11076
rect 22284 11024 22336 11076
rect 25044 11092 25096 11144
rect 26608 11092 26660 11144
rect 28264 11092 28316 11144
rect 28908 11092 28960 11144
rect 38016 11160 38068 11212
rect 32772 11135 32824 11144
rect 32772 11101 32781 11135
rect 32781 11101 32815 11135
rect 32815 11101 32824 11135
rect 32772 11092 32824 11101
rect 32864 11135 32916 11144
rect 32864 11101 32873 11135
rect 32873 11101 32907 11135
rect 32907 11101 32916 11135
rect 32864 11092 32916 11101
rect 37648 11135 37700 11144
rect 37648 11101 37657 11135
rect 37657 11101 37691 11135
rect 37691 11101 37700 11135
rect 37648 11092 37700 11101
rect 38752 11092 38804 11144
rect 39120 11135 39172 11144
rect 39120 11101 39129 11135
rect 39129 11101 39163 11135
rect 39163 11101 39172 11135
rect 39120 11092 39172 11101
rect 39304 11092 39356 11144
rect 39948 11092 40000 11144
rect 40684 11092 40736 11144
rect 41328 11135 41380 11144
rect 41328 11101 41337 11135
rect 41337 11101 41371 11135
rect 41371 11101 41380 11135
rect 41328 11092 41380 11101
rect 44272 11203 44324 11212
rect 44272 11169 44281 11203
rect 44281 11169 44315 11203
rect 44315 11169 44324 11203
rect 44272 11160 44324 11169
rect 43352 11092 43404 11144
rect 25320 11024 25372 11076
rect 29920 11024 29972 11076
rect 7380 10956 7432 11008
rect 9772 10956 9824 11008
rect 17960 10956 18012 11008
rect 18880 10956 18932 11008
rect 21272 10956 21324 11008
rect 24768 10999 24820 11008
rect 24768 10965 24777 10999
rect 24777 10965 24811 10999
rect 24811 10965 24820 10999
rect 24768 10956 24820 10965
rect 25136 10999 25188 11008
rect 25136 10965 25145 10999
rect 25145 10965 25179 10999
rect 25179 10965 25188 10999
rect 25136 10956 25188 10965
rect 29644 10956 29696 11008
rect 32588 11067 32640 11076
rect 32588 11033 32597 11067
rect 32597 11033 32631 11067
rect 32631 11033 32640 11067
rect 32588 11024 32640 11033
rect 33232 11024 33284 11076
rect 35440 11024 35492 11076
rect 35532 11024 35584 11076
rect 37924 11067 37976 11076
rect 37924 11033 37959 11067
rect 37959 11033 37976 11067
rect 37924 11024 37976 11033
rect 38108 11024 38160 11076
rect 38476 11024 38528 11076
rect 38936 11024 38988 11076
rect 39028 11067 39080 11076
rect 39028 11033 39037 11067
rect 39037 11033 39071 11067
rect 39071 11033 39080 11067
rect 39028 11024 39080 11033
rect 42984 11024 43036 11076
rect 43536 11024 43588 11076
rect 31024 10956 31076 11008
rect 36728 10956 36780 11008
rect 37464 10999 37516 11008
rect 37464 10965 37473 10999
rect 37473 10965 37507 10999
rect 37507 10965 37516 10999
rect 37464 10956 37516 10965
rect 43168 10956 43220 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 1952 10795 2004 10804
rect 1952 10761 1961 10795
rect 1961 10761 1995 10795
rect 1995 10761 2004 10795
rect 1952 10752 2004 10761
rect 3056 10752 3108 10804
rect 2504 10684 2556 10736
rect 6000 10752 6052 10804
rect 9772 10752 9824 10804
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 12900 10752 12952 10804
rect 15292 10752 15344 10804
rect 18236 10752 18288 10804
rect 19340 10752 19392 10804
rect 22560 10752 22612 10804
rect 7288 10684 7340 10736
rect 7840 10684 7892 10736
rect 940 10548 992 10600
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 2412 10480 2464 10532
rect 3056 10548 3108 10600
rect 6828 10616 6880 10668
rect 7104 10548 7156 10600
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 14372 10684 14424 10736
rect 15844 10684 15896 10736
rect 16488 10684 16540 10736
rect 18328 10684 18380 10736
rect 24768 10684 24820 10736
rect 25136 10752 25188 10804
rect 25688 10795 25740 10804
rect 25688 10761 25697 10795
rect 25697 10761 25731 10795
rect 25731 10761 25740 10795
rect 25688 10752 25740 10761
rect 29920 10752 29972 10804
rect 30380 10752 30432 10804
rect 32588 10752 32640 10804
rect 37648 10752 37700 10804
rect 42984 10795 43036 10804
rect 42984 10761 42993 10795
rect 42993 10761 43027 10795
rect 43027 10761 43036 10795
rect 42984 10752 43036 10761
rect 44272 10795 44324 10804
rect 44272 10761 44281 10795
rect 44281 10761 44315 10795
rect 44315 10761 44324 10795
rect 44272 10752 44324 10761
rect 14464 10659 14516 10668
rect 12716 10616 12768 10625
rect 2688 10480 2740 10532
rect 4068 10480 4120 10532
rect 4620 10480 4672 10532
rect 13820 10548 13872 10600
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 18420 10659 18472 10668
rect 18420 10625 18454 10659
rect 18454 10625 18472 10659
rect 18420 10616 18472 10625
rect 23480 10616 23532 10668
rect 24676 10616 24728 10668
rect 14924 10548 14976 10600
rect 17868 10548 17920 10600
rect 25136 10616 25188 10668
rect 31024 10684 31076 10736
rect 29644 10616 29696 10668
rect 2964 10412 3016 10464
rect 7472 10412 7524 10464
rect 9772 10412 9824 10464
rect 10600 10412 10652 10464
rect 24584 10412 24636 10464
rect 30012 10548 30064 10600
rect 31300 10659 31352 10668
rect 31300 10625 31309 10659
rect 31309 10625 31343 10659
rect 31343 10625 31352 10659
rect 31300 10616 31352 10625
rect 31668 10616 31720 10668
rect 31208 10548 31260 10600
rect 35532 10684 35584 10736
rect 35992 10684 36044 10736
rect 33968 10659 34020 10668
rect 33968 10625 33977 10659
rect 33977 10625 34011 10659
rect 34011 10625 34020 10659
rect 33968 10616 34020 10625
rect 34520 10616 34572 10668
rect 38016 10616 38068 10668
rect 40408 10684 40460 10736
rect 42340 10684 42392 10736
rect 32496 10591 32548 10600
rect 32496 10557 32505 10591
rect 32505 10557 32539 10591
rect 32539 10557 32548 10591
rect 32496 10548 32548 10557
rect 36728 10548 36780 10600
rect 38384 10591 38436 10600
rect 38384 10557 38393 10591
rect 38393 10557 38427 10591
rect 38427 10557 38436 10591
rect 38384 10548 38436 10557
rect 40684 10591 40736 10600
rect 40684 10557 40693 10591
rect 40693 10557 40727 10591
rect 40727 10557 40736 10591
rect 40684 10548 40736 10557
rect 43168 10659 43220 10668
rect 43168 10625 43177 10659
rect 43177 10625 43211 10659
rect 43211 10625 43220 10659
rect 43168 10616 43220 10625
rect 43260 10659 43312 10668
rect 43260 10625 43269 10659
rect 43269 10625 43303 10659
rect 43303 10625 43312 10659
rect 43260 10616 43312 10625
rect 43444 10659 43496 10668
rect 43444 10625 43479 10659
rect 43479 10625 43496 10659
rect 43444 10616 43496 10625
rect 33048 10480 33100 10532
rect 31944 10412 31996 10464
rect 33968 10455 34020 10464
rect 33968 10421 33977 10455
rect 33977 10421 34011 10455
rect 34011 10421 34020 10455
rect 33968 10412 34020 10421
rect 37096 10412 37148 10464
rect 42524 10412 42576 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2596 10140 2648 10192
rect 4068 10140 4120 10192
rect 11060 10140 11112 10192
rect 16580 10183 16632 10192
rect 16580 10149 16589 10183
rect 16589 10149 16623 10183
rect 16623 10149 16632 10183
rect 16580 10140 16632 10149
rect 18420 10183 18472 10192
rect 18420 10149 18429 10183
rect 18429 10149 18463 10183
rect 18463 10149 18472 10183
rect 18420 10140 18472 10149
rect 22284 10208 22336 10260
rect 23940 10208 23992 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 26700 10208 26752 10260
rect 35992 10208 36044 10260
rect 36728 10251 36780 10260
rect 36728 10217 36737 10251
rect 36737 10217 36771 10251
rect 36771 10217 36780 10251
rect 36728 10208 36780 10217
rect 40224 10208 40276 10260
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3056 10115 3108 10124
rect 3056 10081 3065 10115
rect 3065 10081 3099 10115
rect 3099 10081 3108 10115
rect 3056 10072 3108 10081
rect 7564 10072 7616 10124
rect 5908 10004 5960 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 8208 10004 8260 10056
rect 9864 10072 9916 10124
rect 11612 10072 11664 10124
rect 16488 10072 16540 10124
rect 17132 10072 17184 10124
rect 17868 10072 17920 10124
rect 25320 10072 25372 10124
rect 31300 10140 31352 10192
rect 39856 10140 39908 10192
rect 30288 10072 30340 10124
rect 31760 10072 31812 10124
rect 35348 10115 35400 10124
rect 35348 10081 35357 10115
rect 35357 10081 35391 10115
rect 35391 10081 35400 10115
rect 35348 10072 35400 10081
rect 38384 10072 38436 10124
rect 940 9936 992 9988
rect 2412 9868 2464 9920
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 8300 9936 8352 9988
rect 9772 9979 9824 9988
rect 9772 9945 9781 9979
rect 9781 9945 9815 9979
rect 9815 9945 9824 9979
rect 9772 9936 9824 9945
rect 10324 9936 10376 9988
rect 11796 10004 11848 10056
rect 12348 9936 12400 9988
rect 14924 10004 14976 10056
rect 16672 9936 16724 9988
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 17316 10004 17368 10056
rect 17776 9936 17828 9988
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 21272 10047 21324 10056
rect 19248 9936 19300 9988
rect 21272 10013 21306 10047
rect 21306 10013 21324 10047
rect 21272 10004 21324 10013
rect 24676 10004 24728 10056
rect 6644 9868 6696 9920
rect 9680 9868 9732 9920
rect 9956 9868 10008 9920
rect 16764 9868 16816 9920
rect 22100 9936 22152 9988
rect 20076 9868 20128 9920
rect 20996 9868 21048 9920
rect 26148 10004 26200 10056
rect 27068 10004 27120 10056
rect 27344 10047 27396 10056
rect 27344 10013 27353 10047
rect 27353 10013 27387 10047
rect 27387 10013 27396 10047
rect 27344 10004 27396 10013
rect 25044 9936 25096 9988
rect 27712 9936 27764 9988
rect 28908 10004 28960 10056
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 31944 10004 31996 10056
rect 29000 9936 29052 9988
rect 26332 9868 26384 9920
rect 31576 9868 31628 9920
rect 31760 9868 31812 9920
rect 34520 10004 34572 10056
rect 37188 10047 37240 10056
rect 37188 10013 37197 10047
rect 37197 10013 37231 10047
rect 37231 10013 37240 10047
rect 37188 10004 37240 10013
rect 37464 10047 37516 10056
rect 37464 10013 37498 10047
rect 37498 10013 37516 10047
rect 37464 10004 37516 10013
rect 38844 10004 38896 10056
rect 33968 9936 34020 9988
rect 39028 9979 39080 9988
rect 39028 9945 39037 9979
rect 39037 9945 39071 9979
rect 39071 9945 39080 9979
rect 39028 9936 39080 9945
rect 39212 9979 39264 9988
rect 39212 9945 39221 9979
rect 39221 9945 39255 9979
rect 39255 9945 39264 9979
rect 39212 9936 39264 9945
rect 33692 9868 33744 9920
rect 33876 9868 33928 9920
rect 38016 9868 38068 9920
rect 42524 9868 42576 9920
rect 43536 9911 43588 9920
rect 43536 9877 43545 9911
rect 43545 9877 43579 9911
rect 43579 9877 43588 9911
rect 43536 9868 43588 9877
rect 43628 9911 43680 9920
rect 43628 9877 43637 9911
rect 43637 9877 43671 9911
rect 43671 9877 43680 9911
rect 43628 9868 43680 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 6460 9664 6512 9716
rect 2412 9571 2464 9580
rect 2412 9537 2446 9571
rect 2446 9537 2464 9571
rect 2412 9528 2464 9537
rect 6552 9596 6604 9648
rect 8300 9664 8352 9716
rect 9956 9664 10008 9716
rect 16580 9664 16632 9716
rect 17684 9664 17736 9716
rect 9496 9596 9548 9648
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 5448 9528 5500 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 7840 9528 7892 9580
rect 8208 9528 8260 9580
rect 8392 9460 8444 9512
rect 5908 9392 5960 9444
rect 2872 9324 2924 9376
rect 3884 9324 3936 9376
rect 8484 9392 8536 9444
rect 9864 9596 9916 9648
rect 11060 9596 11112 9648
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10508 9528 10560 9580
rect 16948 9596 17000 9648
rect 18328 9596 18380 9648
rect 21088 9596 21140 9648
rect 10600 9460 10652 9512
rect 15200 9528 15252 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 17408 9528 17460 9580
rect 19984 9528 20036 9580
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 22284 9596 22336 9648
rect 22560 9528 22612 9580
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26240 9528 26292 9537
rect 26424 9664 26476 9716
rect 27068 9664 27120 9716
rect 30012 9664 30064 9716
rect 31852 9664 31904 9716
rect 39028 9664 39080 9716
rect 43260 9664 43312 9716
rect 43996 9664 44048 9716
rect 26700 9596 26752 9648
rect 26608 9571 26660 9580
rect 26608 9537 26617 9571
rect 26617 9537 26651 9571
rect 26651 9537 26660 9571
rect 26608 9528 26660 9537
rect 28356 9596 28408 9648
rect 11060 9392 11112 9444
rect 15108 9392 15160 9444
rect 16488 9392 16540 9444
rect 22284 9503 22336 9512
rect 22284 9469 22293 9503
rect 22293 9469 22327 9503
rect 22327 9469 22336 9503
rect 22284 9460 22336 9469
rect 27344 9460 27396 9512
rect 27712 9571 27764 9580
rect 27712 9537 27721 9571
rect 27721 9537 27755 9571
rect 27755 9537 27764 9571
rect 27712 9528 27764 9537
rect 27804 9571 27856 9580
rect 27804 9537 27813 9571
rect 27813 9537 27847 9571
rect 27847 9537 27856 9571
rect 27804 9528 27856 9537
rect 28816 9596 28868 9648
rect 29000 9639 29052 9648
rect 29000 9605 29009 9639
rect 29009 9605 29043 9639
rect 29043 9605 29052 9639
rect 29000 9596 29052 9605
rect 30104 9639 30156 9648
rect 30104 9605 30113 9639
rect 30113 9605 30147 9639
rect 30147 9605 30156 9639
rect 30104 9596 30156 9605
rect 36452 9596 36504 9648
rect 37188 9596 37240 9648
rect 28632 9571 28684 9580
rect 28632 9537 28641 9571
rect 28641 9537 28675 9571
rect 28675 9537 28684 9571
rect 28632 9528 28684 9537
rect 30840 9528 30892 9580
rect 31484 9571 31536 9580
rect 31484 9537 31493 9571
rect 31493 9537 31527 9571
rect 31527 9537 31536 9571
rect 31484 9528 31536 9537
rect 31760 9528 31812 9580
rect 32128 9528 32180 9580
rect 31944 9460 31996 9512
rect 32220 9460 32272 9512
rect 33692 9528 33744 9580
rect 38660 9528 38712 9580
rect 39028 9571 39080 9580
rect 39028 9537 39037 9571
rect 39037 9537 39071 9571
rect 39071 9537 39080 9571
rect 39028 9528 39080 9537
rect 33968 9460 34020 9512
rect 34060 9503 34112 9512
rect 34060 9469 34069 9503
rect 34069 9469 34103 9503
rect 34103 9469 34112 9503
rect 34060 9460 34112 9469
rect 36084 9460 36136 9512
rect 23480 9392 23532 9444
rect 24676 9392 24728 9444
rect 28080 9435 28132 9444
rect 28080 9401 28089 9435
rect 28089 9401 28123 9435
rect 28123 9401 28132 9435
rect 28080 9392 28132 9401
rect 28632 9392 28684 9444
rect 36544 9392 36596 9444
rect 8116 9324 8168 9376
rect 8852 9324 8904 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 11704 9324 11756 9376
rect 12900 9324 12952 9376
rect 16028 9324 16080 9376
rect 17132 9324 17184 9376
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 21272 9324 21324 9376
rect 21456 9324 21508 9376
rect 25412 9324 25464 9376
rect 31484 9367 31536 9376
rect 31484 9333 31493 9367
rect 31493 9333 31527 9367
rect 31527 9333 31536 9367
rect 31484 9324 31536 9333
rect 32956 9324 33008 9376
rect 33048 9324 33100 9376
rect 39212 9571 39264 9580
rect 39212 9537 39221 9571
rect 39221 9537 39255 9571
rect 39255 9537 39264 9571
rect 39212 9528 39264 9537
rect 39856 9571 39908 9580
rect 39856 9537 39865 9571
rect 39865 9537 39899 9571
rect 39899 9537 39908 9571
rect 39856 9528 39908 9537
rect 40776 9528 40828 9580
rect 40684 9503 40736 9512
rect 40684 9469 40693 9503
rect 40693 9469 40727 9503
rect 40727 9469 40736 9503
rect 40684 9460 40736 9469
rect 40960 9324 41012 9376
rect 43628 9392 43680 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 7104 9120 7156 9172
rect 8116 9163 8168 9172
rect 8116 9129 8125 9163
rect 8125 9129 8159 9163
rect 8159 9129 8168 9163
rect 8116 9120 8168 9129
rect 8300 9120 8352 9172
rect 9588 9120 9640 9172
rect 12164 9120 12216 9172
rect 12348 9120 12400 9172
rect 28632 9120 28684 9172
rect 10508 9052 10560 9104
rect 1124 8984 1176 9036
rect 940 8916 992 8968
rect 5724 8916 5776 8968
rect 6552 8916 6604 8968
rect 1032 8848 1084 8900
rect 7196 8848 7248 8900
rect 7472 8891 7524 8900
rect 7472 8857 7497 8891
rect 7497 8857 7524 8891
rect 7748 8916 7800 8968
rect 7472 8848 7524 8857
rect 8668 8848 8720 8900
rect 5908 8780 5960 8832
rect 8300 8780 8352 8832
rect 9956 8984 10008 9036
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 11520 8916 11572 8968
rect 14280 9052 14332 9104
rect 16948 9052 17000 9104
rect 17224 9052 17276 9104
rect 17500 9052 17552 9104
rect 12900 8984 12952 9036
rect 19156 9052 19208 9104
rect 30656 9120 30708 9172
rect 36544 9120 36596 9172
rect 42248 9120 42300 9172
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 10968 8848 11020 8900
rect 16120 8916 16172 8968
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 12072 8848 12124 8900
rect 16028 8848 16080 8900
rect 17132 8916 17184 8968
rect 20352 8984 20404 9036
rect 21456 9027 21508 9036
rect 21456 8993 21465 9027
rect 21465 8993 21499 9027
rect 21499 8993 21508 9027
rect 21456 8984 21508 8993
rect 21640 9027 21692 9036
rect 21640 8993 21649 9027
rect 21649 8993 21683 9027
rect 21683 8993 21692 9027
rect 21640 8984 21692 8993
rect 19156 8916 19208 8968
rect 16764 8848 16816 8900
rect 12164 8780 12216 8832
rect 12256 8780 12308 8832
rect 12532 8780 12584 8832
rect 12624 8780 12676 8832
rect 17684 8848 17736 8900
rect 21548 8959 21600 8968
rect 21548 8925 21557 8959
rect 21557 8925 21591 8959
rect 21591 8925 21600 8959
rect 21548 8916 21600 8925
rect 25320 8984 25372 9036
rect 25964 8916 26016 8968
rect 26608 8984 26660 9036
rect 32864 9052 32916 9104
rect 36636 9052 36688 9104
rect 38844 9052 38896 9104
rect 37188 9027 37240 9036
rect 37188 8993 37197 9027
rect 37197 8993 37231 9027
rect 37231 8993 37240 9027
rect 37188 8984 37240 8993
rect 19340 8848 19392 8900
rect 22100 8848 22152 8900
rect 22560 8848 22612 8900
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 30288 8916 30340 8968
rect 31392 8916 31444 8968
rect 32864 8916 32916 8968
rect 26608 8848 26660 8900
rect 28908 8848 28960 8900
rect 29276 8848 29328 8900
rect 31484 8848 31536 8900
rect 26148 8780 26200 8832
rect 26240 8780 26292 8832
rect 29644 8780 29696 8832
rect 32220 8848 32272 8900
rect 33232 8848 33284 8900
rect 36452 8959 36504 8968
rect 36452 8925 36461 8959
rect 36461 8925 36495 8959
rect 36495 8925 36504 8959
rect 36452 8916 36504 8925
rect 37556 8916 37608 8968
rect 40132 8916 40184 8968
rect 39212 8848 39264 8900
rect 40316 8848 40368 8900
rect 32128 8780 32180 8832
rect 34612 8780 34664 8832
rect 34796 8780 34848 8832
rect 37556 8780 37608 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 7748 8576 7800 8628
rect 9496 8576 9548 8628
rect 10968 8576 11020 8628
rect 12072 8619 12124 8628
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 12164 8576 12216 8628
rect 16672 8576 16724 8628
rect 17132 8576 17184 8628
rect 17684 8576 17736 8628
rect 19432 8576 19484 8628
rect 1032 8508 1084 8560
rect 5172 8440 5224 8492
rect 5632 8440 5684 8492
rect 7196 8440 7248 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 940 8372 992 8424
rect 5080 8415 5132 8424
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 7472 8372 7524 8424
rect 10324 8508 10376 8560
rect 11244 8440 11296 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 13728 8440 13780 8492
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 22376 8576 22428 8628
rect 22928 8576 22980 8628
rect 14188 8440 14240 8449
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8116 8372 8168 8424
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 5448 8347 5500 8356
rect 5448 8313 5457 8347
rect 5457 8313 5491 8347
rect 5491 8313 5500 8347
rect 5448 8304 5500 8313
rect 8392 8304 8444 8356
rect 8944 8304 8996 8356
rect 9956 8304 10008 8356
rect 10508 8372 10560 8424
rect 10968 8372 11020 8424
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 14924 8440 14976 8492
rect 22560 8508 22612 8560
rect 16212 8372 16264 8424
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 19892 8440 19944 8492
rect 20352 8483 20404 8492
rect 20352 8449 20361 8483
rect 20361 8449 20395 8483
rect 20395 8449 20404 8483
rect 20352 8440 20404 8449
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 22376 8440 22428 8492
rect 16488 8304 16540 8356
rect 19984 8372 20036 8424
rect 17408 8304 17460 8356
rect 20168 8415 20220 8424
rect 20168 8381 20177 8415
rect 20177 8381 20211 8415
rect 20211 8381 20220 8415
rect 20168 8372 20220 8381
rect 10324 8236 10376 8288
rect 11704 8236 11756 8288
rect 14004 8236 14056 8288
rect 20812 8236 20864 8288
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 22008 8372 22060 8424
rect 22744 8440 22796 8492
rect 31852 8508 31904 8560
rect 32864 8551 32916 8560
rect 32864 8517 32873 8551
rect 32873 8517 32907 8551
rect 32907 8517 32916 8551
rect 32864 8508 32916 8517
rect 33048 8508 33100 8560
rect 34796 8576 34848 8628
rect 25412 8483 25464 8492
rect 25412 8449 25446 8483
rect 25446 8449 25464 8483
rect 25412 8440 25464 8449
rect 25872 8440 25924 8492
rect 31944 8440 31996 8492
rect 32128 8440 32180 8492
rect 33324 8483 33376 8492
rect 33324 8449 33333 8483
rect 33333 8449 33367 8483
rect 33367 8449 33376 8483
rect 33324 8440 33376 8449
rect 31760 8372 31812 8424
rect 32496 8372 32548 8424
rect 32772 8372 32824 8424
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35900 8508 35952 8560
rect 35992 8508 36044 8560
rect 35716 8440 35768 8492
rect 37740 8508 37792 8560
rect 36636 8483 36688 8492
rect 36636 8449 36645 8483
rect 36645 8449 36679 8483
rect 36679 8449 36688 8483
rect 36636 8440 36688 8449
rect 22100 8304 22152 8356
rect 26332 8304 26384 8356
rect 35900 8372 35952 8424
rect 36176 8372 36228 8424
rect 36728 8372 36780 8424
rect 37556 8372 37608 8424
rect 39488 8619 39540 8628
rect 39488 8585 39497 8619
rect 39497 8585 39531 8619
rect 39531 8585 39540 8619
rect 39488 8576 39540 8585
rect 40408 8508 40460 8560
rect 38844 8440 38896 8492
rect 38016 8372 38068 8424
rect 43444 8576 43496 8628
rect 40776 8508 40828 8560
rect 40868 8483 40920 8492
rect 40868 8449 40877 8483
rect 40877 8449 40911 8483
rect 40911 8449 40920 8483
rect 40868 8440 40920 8449
rect 40040 8415 40092 8424
rect 40040 8381 40049 8415
rect 40049 8381 40083 8415
rect 40083 8381 40092 8415
rect 40040 8372 40092 8381
rect 40132 8372 40184 8424
rect 41512 8372 41564 8424
rect 40684 8304 40736 8356
rect 21640 8236 21692 8288
rect 22192 8236 22244 8288
rect 25780 8236 25832 8288
rect 33876 8236 33928 8288
rect 35348 8236 35400 8288
rect 37832 8279 37884 8288
rect 37832 8245 37841 8279
rect 37841 8245 37875 8279
rect 37875 8245 37884 8279
rect 37832 8236 37884 8245
rect 40592 8236 40644 8288
rect 54116 8236 54168 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2320 8032 2372 8084
rect 5080 8032 5132 8084
rect 5172 8032 5224 8084
rect 9956 8032 10008 8084
rect 10968 8032 11020 8084
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 12348 8032 12400 8084
rect 15016 8032 15068 8084
rect 16488 8032 16540 8084
rect 10232 8007 10284 8016
rect 10232 7973 10241 8007
rect 10241 7973 10275 8007
rect 10275 7973 10284 8007
rect 10232 7964 10284 7973
rect 10600 7964 10652 8016
rect 13544 7964 13596 8016
rect 1768 7828 1820 7880
rect 4620 7828 4672 7880
rect 7196 7828 7248 7880
rect 8116 7828 8168 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 11152 7896 11204 7948
rect 11612 7896 11664 7948
rect 14280 7964 14332 8016
rect 17776 7964 17828 8016
rect 20720 8032 20772 8084
rect 21180 8032 21232 8084
rect 21640 8075 21692 8084
rect 21640 8041 21649 8075
rect 21649 8041 21683 8075
rect 21683 8041 21692 8075
rect 21640 8032 21692 8041
rect 22744 8032 22796 8084
rect 14004 7896 14056 7948
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 14188 7828 14240 7880
rect 14924 7896 14976 7948
rect 17868 7896 17920 7948
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 22560 7964 22612 8016
rect 26240 8032 26292 8084
rect 27344 8032 27396 8084
rect 40592 8032 40644 8084
rect 30748 7964 30800 8016
rect 25872 7939 25924 7948
rect 25872 7905 25881 7939
rect 25881 7905 25915 7939
rect 25915 7905 25924 7939
rect 25872 7896 25924 7905
rect 1952 7803 2004 7812
rect 1952 7769 1986 7803
rect 1986 7769 2004 7803
rect 1952 7760 2004 7769
rect 4528 7760 4580 7812
rect 7104 7760 7156 7812
rect 7748 7760 7800 7812
rect 11244 7760 11296 7812
rect 4712 7692 4764 7744
rect 8852 7692 8904 7744
rect 11152 7692 11204 7744
rect 14096 7692 14148 7744
rect 15292 7828 15344 7880
rect 18328 7828 18380 7880
rect 15752 7760 15804 7812
rect 17408 7760 17460 7812
rect 17776 7760 17828 7812
rect 19340 7828 19392 7880
rect 19984 7828 20036 7880
rect 22560 7871 22612 7880
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 22560 7828 22612 7837
rect 23112 7828 23164 7880
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 26148 7871 26200 7880
rect 26148 7837 26182 7871
rect 26182 7837 26200 7871
rect 19156 7760 19208 7812
rect 20904 7760 20956 7812
rect 22928 7760 22980 7812
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 22100 7692 22152 7744
rect 26148 7828 26200 7837
rect 31576 7871 31628 7880
rect 31576 7837 31585 7871
rect 31585 7837 31619 7871
rect 31619 7837 31628 7871
rect 31576 7828 31628 7837
rect 31668 7871 31720 7880
rect 31668 7837 31677 7871
rect 31677 7837 31711 7871
rect 31711 7837 31720 7871
rect 33232 7964 33284 8016
rect 33600 7964 33652 8016
rect 32404 7896 32456 7948
rect 32864 7896 32916 7948
rect 35348 7939 35400 7948
rect 35348 7905 35357 7939
rect 35357 7905 35391 7939
rect 35391 7905 35400 7939
rect 35348 7896 35400 7905
rect 31668 7828 31720 7837
rect 32404 7760 32456 7812
rect 33048 7828 33100 7880
rect 33140 7828 33192 7880
rect 34060 7828 34112 7880
rect 34796 7828 34848 7880
rect 33232 7760 33284 7812
rect 33784 7760 33836 7812
rect 40316 7896 40368 7948
rect 35992 7871 36044 7880
rect 35992 7837 36001 7871
rect 36001 7837 36035 7871
rect 36035 7837 36044 7871
rect 35992 7828 36044 7837
rect 37832 7828 37884 7880
rect 40040 7871 40092 7880
rect 40040 7837 40049 7871
rect 40049 7837 40083 7871
rect 40083 7837 40092 7871
rect 40040 7828 40092 7837
rect 41052 7828 41104 7880
rect 41512 7871 41564 7880
rect 41512 7837 41546 7871
rect 41546 7837 41564 7871
rect 41512 7828 41564 7837
rect 40132 7760 40184 7812
rect 40224 7803 40276 7812
rect 40224 7769 40233 7803
rect 40233 7769 40267 7803
rect 40267 7769 40276 7803
rect 40224 7760 40276 7769
rect 33140 7692 33192 7744
rect 33416 7692 33468 7744
rect 34336 7692 34388 7744
rect 35624 7692 35676 7744
rect 38660 7692 38712 7744
rect 40408 7692 40460 7744
rect 43260 7692 43312 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 1952 7531 2004 7540
rect 1952 7497 1961 7531
rect 1961 7497 1995 7531
rect 1995 7497 2004 7531
rect 1952 7488 2004 7497
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5172 7488 5224 7540
rect 9772 7488 9824 7540
rect 13360 7488 13412 7540
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 20812 7488 20864 7540
rect 940 7420 992 7472
rect 11152 7420 11204 7472
rect 11704 7463 11756 7472
rect 11704 7429 11713 7463
rect 11713 7429 11747 7463
rect 11747 7429 11756 7463
rect 11704 7420 11756 7429
rect 14096 7420 14148 7472
rect 5724 7352 5776 7404
rect 7196 7352 7248 7404
rect 10324 7352 10376 7404
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 2412 7284 2464 7336
rect 2596 7284 2648 7336
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11060 7284 11112 7336
rect 12072 7284 12124 7336
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 17776 7420 17828 7472
rect 20260 7420 20312 7472
rect 27344 7488 27396 7540
rect 32404 7531 32456 7540
rect 32404 7497 32413 7531
rect 32413 7497 32447 7531
rect 32447 7497 32456 7531
rect 32404 7488 32456 7497
rect 22560 7420 22612 7472
rect 33324 7488 33376 7540
rect 37740 7531 37792 7540
rect 37740 7497 37749 7531
rect 37749 7497 37783 7531
rect 37783 7497 37792 7531
rect 37740 7488 37792 7497
rect 42616 7420 42668 7472
rect 16672 7352 16724 7404
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 19616 7395 19668 7404
rect 19616 7361 19625 7395
rect 19625 7361 19659 7395
rect 19659 7361 19668 7395
rect 19616 7352 19668 7361
rect 20076 7352 20128 7404
rect 24676 7352 24728 7404
rect 30380 7352 30432 7404
rect 31300 7352 31352 7404
rect 32404 7352 32456 7404
rect 32680 7395 32732 7404
rect 32680 7361 32689 7395
rect 32689 7361 32723 7395
rect 32723 7361 32732 7395
rect 32680 7352 32732 7361
rect 17040 7284 17092 7336
rect 23020 7327 23072 7336
rect 23020 7293 23029 7327
rect 23029 7293 23063 7327
rect 23063 7293 23072 7327
rect 23020 7284 23072 7293
rect 23112 7327 23164 7336
rect 23112 7293 23121 7327
rect 23121 7293 23155 7327
rect 23155 7293 23164 7327
rect 23112 7284 23164 7293
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 10232 7148 10284 7200
rect 10508 7148 10560 7200
rect 17224 7216 17276 7268
rect 30840 7284 30892 7336
rect 32864 7284 32916 7336
rect 33416 7395 33468 7404
rect 33416 7361 33425 7395
rect 33425 7361 33459 7395
rect 33459 7361 33468 7395
rect 33416 7352 33468 7361
rect 33876 7352 33928 7404
rect 34336 7352 34388 7404
rect 38660 7352 38712 7404
rect 39212 7352 39264 7404
rect 42800 7395 42852 7404
rect 42800 7361 42809 7395
rect 42809 7361 42843 7395
rect 42843 7361 42852 7395
rect 42800 7352 42852 7361
rect 33692 7284 33744 7336
rect 38200 7327 38252 7336
rect 38200 7293 38209 7327
rect 38209 7293 38243 7327
rect 38243 7293 38252 7327
rect 38200 7284 38252 7293
rect 38384 7327 38436 7336
rect 38384 7293 38393 7327
rect 38393 7293 38427 7327
rect 38427 7293 38436 7327
rect 38384 7284 38436 7293
rect 41696 7284 41748 7336
rect 11980 7148 12032 7200
rect 14556 7148 14608 7200
rect 33048 7216 33100 7268
rect 33232 7216 33284 7268
rect 39028 7216 39080 7268
rect 40224 7216 40276 7268
rect 22744 7191 22796 7200
rect 22744 7157 22753 7191
rect 22753 7157 22787 7191
rect 22787 7157 22796 7191
rect 22744 7148 22796 7157
rect 32036 7148 32088 7200
rect 32772 7148 32824 7200
rect 32956 7148 33008 7200
rect 33416 7148 33468 7200
rect 42984 7191 43036 7200
rect 42984 7157 42993 7191
rect 42993 7157 43027 7191
rect 43027 7157 43036 7191
rect 42984 7148 43036 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12440 6944 12492 6996
rect 13452 6944 13504 6996
rect 16672 6987 16724 6996
rect 16672 6953 16681 6987
rect 16681 6953 16715 6987
rect 16715 6953 16724 6987
rect 16672 6944 16724 6953
rect 17224 6944 17276 6996
rect 33784 6944 33836 6996
rect 2596 6808 2648 6860
rect 4804 6808 4856 6860
rect 8392 6808 8444 6860
rect 11060 6876 11112 6928
rect 10876 6808 10928 6860
rect 22008 6851 22060 6860
rect 22008 6817 22017 6851
rect 22017 6817 22051 6851
rect 22051 6817 22060 6851
rect 22008 6808 22060 6817
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 30012 6851 30064 6860
rect 30012 6817 30021 6851
rect 30021 6817 30055 6851
rect 30055 6817 30064 6851
rect 30012 6808 30064 6817
rect 32864 6876 32916 6928
rect 940 6740 992 6792
rect 8024 6740 8076 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 13452 6740 13504 6792
rect 15108 6740 15160 6792
rect 17408 6740 17460 6792
rect 17500 6740 17552 6792
rect 19248 6740 19300 6792
rect 19616 6740 19668 6792
rect 22744 6740 22796 6792
rect 24492 6740 24544 6792
rect 26424 6740 26476 6792
rect 29276 6740 29328 6792
rect 29920 6783 29972 6792
rect 29920 6749 29929 6783
rect 29929 6749 29963 6783
rect 29963 6749 29972 6783
rect 29920 6740 29972 6749
rect 30104 6783 30156 6792
rect 30104 6749 30113 6783
rect 30113 6749 30147 6783
rect 30147 6749 30156 6783
rect 30104 6740 30156 6749
rect 30288 6783 30340 6792
rect 30288 6749 30297 6783
rect 30297 6749 30331 6783
rect 30331 6749 30340 6783
rect 30288 6740 30340 6749
rect 30840 6740 30892 6792
rect 31208 6783 31260 6792
rect 31208 6749 31217 6783
rect 31217 6749 31251 6783
rect 31251 6749 31260 6783
rect 31208 6740 31260 6749
rect 31392 6783 31444 6792
rect 31392 6749 31401 6783
rect 31401 6749 31435 6783
rect 31435 6749 31444 6783
rect 31392 6740 31444 6749
rect 31760 6808 31812 6860
rect 8300 6672 8352 6724
rect 9036 6672 9088 6724
rect 10876 6715 10928 6724
rect 10876 6681 10885 6715
rect 10885 6681 10919 6715
rect 10919 6681 10928 6715
rect 10876 6672 10928 6681
rect 11060 6672 11112 6724
rect 11612 6672 11664 6724
rect 11796 6715 11848 6724
rect 11796 6681 11830 6715
rect 11830 6681 11848 6715
rect 11796 6672 11848 6681
rect 17224 6672 17276 6724
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 3424 6604 3476 6656
rect 9864 6604 9916 6656
rect 11704 6604 11756 6656
rect 12164 6604 12216 6656
rect 16672 6604 16724 6656
rect 22100 6604 22152 6656
rect 30472 6647 30524 6656
rect 30472 6613 30481 6647
rect 30481 6613 30515 6647
rect 30515 6613 30524 6647
rect 30472 6604 30524 6613
rect 32036 6783 32088 6792
rect 32036 6749 32045 6783
rect 32045 6749 32079 6783
rect 32079 6749 32088 6783
rect 32036 6740 32088 6749
rect 32496 6740 32548 6792
rect 32312 6715 32364 6724
rect 32312 6681 32321 6715
rect 32321 6681 32355 6715
rect 32355 6681 32364 6715
rect 32312 6672 32364 6681
rect 31944 6604 31996 6656
rect 35716 6808 35768 6860
rect 33140 6783 33192 6792
rect 33140 6749 33174 6783
rect 33174 6749 33192 6783
rect 33140 6740 33192 6749
rect 35532 6783 35584 6792
rect 35532 6749 35541 6783
rect 35541 6749 35575 6783
rect 35575 6749 35584 6783
rect 35532 6740 35584 6749
rect 35624 6783 35676 6792
rect 35624 6749 35633 6783
rect 35633 6749 35667 6783
rect 35667 6749 35676 6783
rect 35624 6740 35676 6749
rect 34520 6604 34572 6656
rect 35808 6647 35860 6656
rect 35808 6613 35817 6647
rect 35817 6613 35851 6647
rect 35851 6613 35860 6647
rect 35808 6604 35860 6613
rect 36452 6715 36504 6724
rect 36452 6681 36461 6715
rect 36461 6681 36495 6715
rect 36495 6681 36504 6715
rect 36452 6672 36504 6681
rect 36728 6672 36780 6724
rect 41052 6740 41104 6792
rect 42984 6740 43036 6792
rect 36544 6604 36596 6656
rect 38384 6604 38436 6656
rect 42156 6672 42208 6724
rect 44272 6740 44324 6792
rect 42892 6604 42944 6656
rect 43076 6604 43128 6656
rect 43996 6604 44048 6656
rect 44364 6604 44416 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 2504 6400 2556 6452
rect 2136 6375 2188 6384
rect 2136 6341 2170 6375
rect 2170 6341 2188 6375
rect 2136 6332 2188 6341
rect 8392 6400 8444 6452
rect 8944 6400 8996 6452
rect 9036 6400 9088 6452
rect 7288 6375 7340 6384
rect 7288 6341 7297 6375
rect 7297 6341 7331 6375
rect 7331 6341 7340 6375
rect 7288 6332 7340 6341
rect 8024 6332 8076 6384
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 11060 6400 11112 6452
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 1768 6196 1820 6248
rect 5816 6264 5868 6316
rect 7564 6264 7616 6316
rect 13176 6332 13228 6384
rect 6552 6196 6604 6248
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 11336 6264 11388 6316
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12164 6307 12216 6316
rect 12164 6273 12173 6307
rect 12173 6273 12207 6307
rect 12207 6273 12216 6307
rect 12164 6264 12216 6273
rect 14004 6332 14056 6384
rect 14096 6375 14148 6384
rect 14096 6341 14121 6375
rect 14121 6341 14148 6375
rect 17408 6400 17460 6452
rect 14096 6332 14148 6341
rect 14740 6332 14792 6384
rect 17500 6332 17552 6384
rect 26148 6332 26200 6384
rect 13544 6264 13596 6316
rect 20444 6264 20496 6316
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 22100 6307 22152 6316
rect 22100 6273 22110 6307
rect 22110 6273 22144 6307
rect 22144 6273 22152 6307
rect 22100 6264 22152 6273
rect 1584 6060 1636 6112
rect 9680 6128 9732 6180
rect 22560 6264 22612 6316
rect 25320 6307 25372 6316
rect 25320 6273 25329 6307
rect 25329 6273 25363 6307
rect 25363 6273 25372 6307
rect 25320 6264 25372 6273
rect 25412 6264 25464 6316
rect 25596 6307 25648 6316
rect 25596 6273 25605 6307
rect 25605 6273 25639 6307
rect 25639 6273 25648 6307
rect 25596 6264 25648 6273
rect 29736 6332 29788 6384
rect 29920 6332 29972 6384
rect 32680 6332 32732 6384
rect 30472 6264 30524 6316
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 10876 6128 10928 6180
rect 11428 6128 11480 6180
rect 12532 6128 12584 6180
rect 12624 6060 12676 6112
rect 14004 6060 14056 6112
rect 17224 6196 17276 6248
rect 18788 6196 18840 6248
rect 19156 6239 19208 6248
rect 19156 6205 19165 6239
rect 19165 6205 19199 6239
rect 19199 6205 19208 6239
rect 19156 6196 19208 6205
rect 19248 6239 19300 6248
rect 19248 6205 19257 6239
rect 19257 6205 19291 6239
rect 19291 6205 19300 6239
rect 19248 6196 19300 6205
rect 22376 6196 22428 6248
rect 23112 6196 23164 6248
rect 30656 6196 30708 6248
rect 33140 6196 33192 6248
rect 33600 6196 33652 6248
rect 34520 6400 34572 6452
rect 35624 6400 35676 6452
rect 34152 6332 34204 6384
rect 34336 6264 34388 6316
rect 35532 6264 35584 6316
rect 37648 6307 37700 6316
rect 37648 6273 37657 6307
rect 37657 6273 37691 6307
rect 37691 6273 37700 6307
rect 37648 6264 37700 6273
rect 37832 6307 37884 6316
rect 37832 6273 37841 6307
rect 37841 6273 37875 6307
rect 37875 6273 37884 6307
rect 37832 6264 37884 6273
rect 38016 6307 38068 6316
rect 38016 6273 38025 6307
rect 38025 6273 38059 6307
rect 38059 6273 38068 6307
rect 38016 6264 38068 6273
rect 42800 6400 42852 6452
rect 42892 6400 42944 6452
rect 42156 6332 42208 6384
rect 40132 6264 40184 6316
rect 43076 6307 43128 6316
rect 43076 6273 43085 6307
rect 43085 6273 43119 6307
rect 43119 6273 43128 6307
rect 43076 6264 43128 6273
rect 44088 6400 44140 6452
rect 44272 6443 44324 6452
rect 44272 6409 44281 6443
rect 44281 6409 44315 6443
rect 44315 6409 44324 6443
rect 44272 6400 44324 6409
rect 45284 6264 45336 6316
rect 14832 6128 14884 6180
rect 22192 6128 22244 6180
rect 22652 6171 22704 6180
rect 22652 6137 22661 6171
rect 22661 6137 22695 6171
rect 22695 6137 22704 6171
rect 22652 6128 22704 6137
rect 14464 6060 14516 6112
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 25136 6060 25188 6069
rect 26608 6060 26660 6112
rect 29920 6060 29972 6112
rect 30288 6060 30340 6112
rect 32680 6128 32732 6180
rect 34152 6060 34204 6112
rect 35992 6196 36044 6248
rect 36360 6196 36412 6248
rect 40040 6103 40092 6112
rect 40040 6069 40049 6103
rect 40049 6069 40083 6103
rect 40083 6069 40092 6103
rect 40040 6060 40092 6069
rect 40316 6060 40368 6112
rect 43076 6128 43128 6180
rect 43628 6060 43680 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 940 5720 992 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 3424 5856 3476 5908
rect 6920 5856 6972 5908
rect 7104 5856 7156 5908
rect 9864 5856 9916 5908
rect 11520 5856 11572 5908
rect 12348 5899 12400 5908
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 18788 5899 18840 5908
rect 18788 5865 18797 5899
rect 18797 5865 18831 5899
rect 18831 5865 18840 5899
rect 18788 5856 18840 5865
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 9312 5788 9364 5840
rect 11244 5788 11296 5840
rect 11336 5788 11388 5840
rect 11980 5788 12032 5840
rect 20444 5788 20496 5840
rect 26608 5856 26660 5908
rect 29276 5856 29328 5908
rect 30656 5856 30708 5908
rect 37832 5856 37884 5908
rect 33048 5788 33100 5840
rect 4160 5720 4212 5772
rect 6920 5720 6972 5772
rect 8668 5720 8720 5772
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 7012 5652 7064 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10876 5720 10928 5772
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11152 5695 11204 5704
rect 11152 5661 11162 5695
rect 11162 5661 11196 5695
rect 11196 5661 11204 5695
rect 11152 5652 11204 5661
rect 11428 5695 11480 5704
rect 2596 5584 2648 5636
rect 3424 5584 3476 5636
rect 4804 5627 4856 5636
rect 4804 5593 4813 5627
rect 4813 5593 4847 5627
rect 4847 5593 4856 5627
rect 4804 5584 4856 5593
rect 6828 5584 6880 5636
rect 9680 5584 9732 5636
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 19432 5763 19484 5772
rect 19432 5729 19441 5763
rect 19441 5729 19475 5763
rect 19475 5729 19484 5763
rect 19432 5720 19484 5729
rect 20812 5720 20864 5772
rect 22008 5720 22060 5772
rect 25504 5720 25556 5772
rect 25872 5720 25924 5772
rect 35808 5720 35860 5772
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 18512 5652 18564 5704
rect 18880 5652 18932 5704
rect 22100 5652 22152 5704
rect 23388 5652 23440 5704
rect 25136 5652 25188 5704
rect 31944 5652 31996 5704
rect 11336 5627 11388 5636
rect 11336 5593 11345 5627
rect 11345 5593 11379 5627
rect 11379 5593 11388 5627
rect 11336 5584 11388 5593
rect 12072 5584 12124 5636
rect 12348 5627 12400 5636
rect 12348 5593 12373 5627
rect 12373 5593 12400 5627
rect 12348 5584 12400 5593
rect 14648 5627 14700 5636
rect 14648 5593 14657 5627
rect 14657 5593 14691 5627
rect 14691 5593 14700 5627
rect 14648 5584 14700 5593
rect 18696 5584 18748 5636
rect 4712 5516 4764 5568
rect 7932 5559 7984 5568
rect 7932 5525 7950 5559
rect 7950 5525 7984 5559
rect 7932 5516 7984 5525
rect 10600 5516 10652 5568
rect 11980 5516 12032 5568
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 22744 5584 22796 5636
rect 25320 5584 25372 5636
rect 29736 5584 29788 5636
rect 27344 5559 27396 5568
rect 27344 5525 27353 5559
rect 27353 5525 27387 5559
rect 27387 5525 27396 5559
rect 27344 5516 27396 5525
rect 30288 5516 30340 5568
rect 30380 5516 30432 5568
rect 33232 5559 33284 5568
rect 33232 5525 33241 5559
rect 33241 5525 33275 5559
rect 33275 5525 33284 5559
rect 33232 5516 33284 5525
rect 33600 5695 33652 5704
rect 33600 5661 33609 5695
rect 33609 5661 33643 5695
rect 33643 5661 33652 5695
rect 33600 5652 33652 5661
rect 34796 5652 34848 5704
rect 35900 5652 35952 5704
rect 36360 5695 36412 5704
rect 36360 5661 36369 5695
rect 36369 5661 36403 5695
rect 36403 5661 36412 5695
rect 36360 5652 36412 5661
rect 40040 5695 40092 5704
rect 40040 5661 40049 5695
rect 40049 5661 40083 5695
rect 40083 5661 40092 5695
rect 40040 5652 40092 5661
rect 40224 5695 40276 5704
rect 40224 5661 40233 5695
rect 40233 5661 40267 5695
rect 40267 5661 40276 5695
rect 40224 5652 40276 5661
rect 40408 5695 40460 5704
rect 40408 5661 40417 5695
rect 40417 5661 40451 5695
rect 40451 5661 40460 5695
rect 40408 5652 40460 5661
rect 34336 5584 34388 5636
rect 40316 5627 40368 5636
rect 40316 5593 40325 5627
rect 40325 5593 40359 5627
rect 40359 5593 40368 5627
rect 40316 5584 40368 5593
rect 35992 5516 36044 5568
rect 36452 5516 36504 5568
rect 44272 5856 44324 5908
rect 41052 5720 41104 5772
rect 43628 5763 43680 5772
rect 43628 5729 43637 5763
rect 43637 5729 43671 5763
rect 43671 5729 43680 5763
rect 43628 5720 43680 5729
rect 42892 5652 42944 5704
rect 43444 5695 43496 5704
rect 43444 5661 43479 5695
rect 43479 5661 43496 5695
rect 43444 5652 43496 5661
rect 41144 5516 41196 5568
rect 42340 5516 42392 5568
rect 42800 5516 42852 5568
rect 43628 5584 43680 5636
rect 43996 5516 44048 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 940 5244 992 5296
rect 3424 5244 3476 5296
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 940 5108 992 5160
rect 1032 5040 1084 5092
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 5540 5244 5592 5296
rect 7564 5312 7616 5364
rect 8668 5312 8720 5364
rect 3056 5108 3108 5160
rect 5080 5176 5132 5228
rect 7288 5176 7340 5228
rect 8116 5244 8168 5296
rect 8300 5244 8352 5296
rect 10508 5244 10560 5296
rect 10876 5312 10928 5364
rect 11888 5312 11940 5364
rect 12348 5312 12400 5364
rect 14096 5312 14148 5364
rect 10600 5176 10652 5228
rect 4620 5108 4672 5160
rect 6276 5108 6328 5160
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 6828 5108 6880 5160
rect 7196 5108 7248 5160
rect 7656 5108 7708 5160
rect 10784 5108 10836 5160
rect 13360 5176 13412 5228
rect 14280 5176 14332 5228
rect 14648 5355 14700 5364
rect 14648 5321 14657 5355
rect 14657 5321 14691 5355
rect 14691 5321 14700 5355
rect 14648 5312 14700 5321
rect 19156 5312 19208 5364
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 27344 5312 27396 5364
rect 16488 5244 16540 5296
rect 18972 5244 19024 5296
rect 23296 5244 23348 5296
rect 23388 5244 23440 5296
rect 23848 5244 23900 5296
rect 27528 5312 27580 5364
rect 27620 5312 27672 5364
rect 27896 5312 27948 5364
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 18512 5176 18564 5228
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 3884 4972 3936 5024
rect 8300 4972 8352 5024
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 10508 5015 10560 5024
rect 10508 4981 10517 5015
rect 10517 4981 10551 5015
rect 10551 4981 10560 5015
rect 10508 4972 10560 4981
rect 15936 5083 15988 5092
rect 15936 5049 15945 5083
rect 15945 5049 15979 5083
rect 15979 5049 15988 5083
rect 15936 5040 15988 5049
rect 17868 5040 17920 5092
rect 18696 5108 18748 5160
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 24032 5219 24084 5228
rect 24032 5185 24041 5219
rect 24041 5185 24075 5219
rect 24075 5185 24084 5219
rect 24032 5176 24084 5185
rect 24492 5219 24544 5228
rect 24492 5185 24501 5219
rect 24501 5185 24535 5219
rect 24535 5185 24544 5219
rect 24492 5176 24544 5185
rect 25504 5176 25556 5228
rect 27344 5219 27396 5228
rect 27344 5185 27351 5219
rect 27351 5185 27396 5219
rect 27344 5176 27396 5185
rect 27528 5219 27580 5226
rect 27528 5185 27537 5219
rect 27537 5185 27571 5219
rect 27571 5185 27580 5219
rect 27528 5174 27580 5185
rect 25596 5040 25648 5092
rect 14004 4972 14056 5024
rect 14740 4972 14792 5024
rect 16212 4972 16264 5024
rect 18236 4972 18288 5024
rect 22192 4972 22244 5024
rect 22560 4972 22612 5024
rect 29276 5176 29328 5228
rect 30012 5244 30064 5296
rect 30288 5312 30340 5364
rect 33600 5312 33652 5364
rect 33968 5312 34020 5364
rect 37832 5312 37884 5364
rect 38200 5312 38252 5364
rect 38384 5312 38436 5364
rect 30104 5219 30156 5228
rect 30104 5185 30113 5219
rect 30113 5185 30147 5219
rect 30147 5185 30156 5219
rect 30104 5176 30156 5185
rect 30380 5176 30432 5228
rect 33232 5244 33284 5296
rect 41144 5244 41196 5296
rect 41696 5312 41748 5364
rect 42800 5312 42852 5364
rect 49700 5312 49752 5364
rect 42340 5244 42392 5296
rect 56968 5244 57020 5296
rect 30012 5151 30064 5160
rect 30012 5117 30021 5151
rect 30021 5117 30055 5151
rect 30055 5117 30064 5151
rect 30012 5108 30064 5117
rect 33876 5108 33928 5160
rect 36360 5151 36412 5160
rect 36360 5117 36369 5151
rect 36369 5117 36403 5151
rect 36403 5117 36412 5151
rect 36360 5108 36412 5117
rect 36544 5151 36596 5160
rect 36544 5117 36553 5151
rect 36553 5117 36587 5151
rect 36587 5117 36596 5151
rect 36544 5108 36596 5117
rect 35992 5040 36044 5092
rect 40040 5040 40092 5092
rect 41420 5219 41472 5228
rect 41420 5185 41429 5219
rect 41429 5185 41463 5219
rect 41463 5185 41472 5219
rect 41420 5176 41472 5185
rect 41788 5219 41840 5228
rect 41788 5185 41797 5219
rect 41797 5185 41831 5219
rect 41831 5185 41840 5219
rect 41788 5176 41840 5185
rect 43444 5108 43496 5160
rect 29736 4972 29788 5024
rect 38292 4972 38344 5024
rect 38752 4972 38804 5024
rect 44180 5151 44232 5160
rect 44180 5117 44189 5151
rect 44189 5117 44223 5151
rect 44223 5117 44232 5151
rect 44180 5108 44232 5117
rect 44640 5108 44692 5160
rect 45284 5151 45336 5160
rect 45284 5117 45293 5151
rect 45293 5117 45327 5151
rect 45327 5117 45336 5151
rect 45284 5108 45336 5117
rect 44824 5015 44876 5024
rect 44824 4981 44833 5015
rect 44833 4981 44867 5015
rect 44867 4981 44876 5015
rect 44824 4972 44876 4981
rect 51632 4972 51684 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4768 1636 4820
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 5724 4768 5776 4820
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 11428 4768 11480 4820
rect 15936 4768 15988 4820
rect 19800 4700 19852 4752
rect 20076 4700 20128 4752
rect 5172 4632 5224 4684
rect 1768 4564 1820 4616
rect 2504 4564 2556 4616
rect 4252 4564 4304 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 3700 4496 3752 4548
rect 4068 4539 4120 4548
rect 4068 4505 4077 4539
rect 4077 4505 4111 4539
rect 4111 4505 4120 4539
rect 4068 4496 4120 4505
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 22652 4768 22704 4820
rect 25136 4768 25188 4820
rect 29828 4768 29880 4820
rect 30012 4768 30064 4820
rect 36544 4768 36596 4820
rect 22836 4700 22888 4752
rect 23664 4700 23716 4752
rect 23756 4632 23808 4684
rect 6920 4564 6972 4616
rect 10508 4607 10560 4616
rect 10508 4573 10542 4607
rect 10542 4573 10560 4607
rect 10508 4564 10560 4573
rect 10784 4564 10836 4616
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 5632 4496 5684 4548
rect 6276 4539 6328 4548
rect 6276 4505 6285 4539
rect 6285 4505 6319 4539
rect 6319 4505 6328 4539
rect 6276 4496 6328 4505
rect 8392 4496 8444 4548
rect 15292 4496 15344 4548
rect 16488 4496 16540 4548
rect 17408 4496 17460 4548
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 6368 4471 6420 4480
rect 6368 4437 6377 4471
rect 6377 4437 6411 4471
rect 6411 4437 6420 4471
rect 6368 4428 6420 4437
rect 7564 4428 7616 4480
rect 14832 4428 14884 4480
rect 16120 4428 16172 4480
rect 17960 4539 18012 4548
rect 17960 4505 17969 4539
rect 17969 4505 18003 4539
rect 18003 4505 18012 4539
rect 17960 4496 18012 4505
rect 18236 4539 18288 4548
rect 18236 4505 18245 4539
rect 18245 4505 18279 4539
rect 18279 4505 18288 4539
rect 18236 4496 18288 4505
rect 19340 4564 19392 4616
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 19984 4564 20036 4616
rect 18512 4496 18564 4548
rect 23848 4564 23900 4616
rect 19984 4428 20036 4480
rect 21824 4428 21876 4480
rect 23940 4496 23992 4548
rect 23756 4428 23808 4480
rect 37648 4700 37700 4752
rect 38016 4700 38068 4752
rect 38384 4700 38436 4752
rect 25872 4632 25924 4684
rect 29920 4675 29972 4684
rect 29920 4641 29929 4675
rect 29929 4641 29963 4675
rect 29963 4641 29972 4675
rect 29920 4632 29972 4641
rect 41420 4768 41472 4820
rect 41696 4768 41748 4820
rect 42892 4768 42944 4820
rect 43996 4768 44048 4820
rect 31208 4564 31260 4616
rect 38016 4607 38068 4616
rect 38016 4573 38025 4607
rect 38025 4573 38059 4607
rect 38059 4573 38068 4607
rect 38016 4564 38068 4573
rect 38108 4607 38160 4616
rect 38108 4573 38143 4607
rect 38143 4573 38160 4607
rect 38108 4564 38160 4573
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 30012 4496 30064 4548
rect 36268 4496 36320 4548
rect 43076 4700 43128 4752
rect 43996 4632 44048 4684
rect 41696 4607 41748 4616
rect 41696 4573 41705 4607
rect 41705 4573 41739 4607
rect 41739 4573 41748 4607
rect 41696 4564 41748 4573
rect 41788 4607 41840 4616
rect 41788 4573 41797 4607
rect 41797 4573 41831 4607
rect 41831 4573 41840 4607
rect 41788 4564 41840 4573
rect 42064 4607 42116 4616
rect 42064 4573 42073 4607
rect 42073 4573 42107 4607
rect 42107 4573 42116 4607
rect 42064 4564 42116 4573
rect 30840 4428 30892 4480
rect 38292 4428 38344 4480
rect 39120 4471 39172 4480
rect 39120 4437 39129 4471
rect 39129 4437 39163 4471
rect 39163 4437 39172 4471
rect 39120 4428 39172 4437
rect 40224 4428 40276 4480
rect 41420 4471 41472 4480
rect 41420 4437 41429 4471
rect 41429 4437 41463 4471
rect 41463 4437 41472 4471
rect 41420 4428 41472 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4068 4224 4120 4276
rect 3056 4156 3108 4208
rect 4252 4199 4304 4208
rect 4252 4165 4261 4199
rect 4261 4165 4295 4199
rect 4295 4165 4304 4199
rect 4252 4156 4304 4165
rect 940 4020 992 4072
rect 3608 4088 3660 4140
rect 3976 4088 4028 4140
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4712 4131 4764 4140
rect 4712 4097 4721 4131
rect 4721 4097 4755 4131
rect 4755 4097 4764 4131
rect 4712 4088 4764 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5356 4156 5408 4208
rect 11704 4224 11756 4276
rect 17592 4224 17644 4276
rect 29368 4224 29420 4276
rect 30748 4224 30800 4276
rect 30840 4224 30892 4276
rect 42064 4224 42116 4276
rect 1124 3952 1176 4004
rect 2320 4020 2372 4072
rect 4160 4020 4212 4072
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 11152 4156 11204 4208
rect 10232 4088 10284 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 5172 4020 5224 4072
rect 7656 4020 7708 4072
rect 12072 4020 12124 4072
rect 12532 4088 12584 4140
rect 17040 4156 17092 4208
rect 17868 4199 17920 4208
rect 17868 4165 17877 4199
rect 17877 4165 17911 4199
rect 17911 4165 17920 4199
rect 17868 4156 17920 4165
rect 24860 4156 24912 4208
rect 30380 4156 30432 4208
rect 14740 4088 14792 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 14924 4088 14976 4140
rect 17960 4088 18012 4140
rect 19248 4088 19300 4140
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 20904 4088 20956 4140
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 23940 4088 23992 4140
rect 29368 4088 29420 4140
rect 29460 4131 29512 4140
rect 29460 4097 29469 4131
rect 29469 4097 29503 4131
rect 29503 4097 29512 4131
rect 29460 4088 29512 4097
rect 29828 4131 29880 4140
rect 29828 4097 29837 4131
rect 29837 4097 29871 4131
rect 29871 4097 29880 4131
rect 29828 4088 29880 4097
rect 30012 4131 30064 4140
rect 30012 4097 30021 4131
rect 30021 4097 30055 4131
rect 30055 4097 30064 4131
rect 30012 4088 30064 4097
rect 15384 4020 15436 4072
rect 20260 4020 20312 4072
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 28908 4020 28960 4072
rect 30104 4020 30156 4072
rect 6828 3952 6880 4004
rect 28540 3952 28592 4004
rect 1952 3884 2004 3936
rect 5080 3884 5132 3936
rect 5816 3884 5868 3936
rect 7932 3884 7984 3936
rect 8392 3884 8444 3936
rect 12440 3884 12492 3936
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 12624 3884 12676 3936
rect 13544 3884 13596 3936
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 16580 3884 16632 3936
rect 24032 3884 24084 3936
rect 27620 3884 27672 3936
rect 29276 3884 29328 3936
rect 31208 4131 31260 4140
rect 31208 4097 31217 4131
rect 31217 4097 31251 4131
rect 31251 4097 31260 4131
rect 31208 4088 31260 4097
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 31760 4156 31812 4208
rect 34520 4156 34572 4208
rect 38660 4156 38712 4208
rect 41788 4156 41840 4208
rect 43628 4224 43680 4276
rect 43996 4267 44048 4276
rect 43996 4233 44005 4267
rect 44005 4233 44039 4267
rect 44039 4233 44048 4267
rect 43996 4224 44048 4233
rect 43076 4199 43128 4208
rect 43076 4165 43111 4199
rect 43111 4165 43128 4199
rect 43076 4156 43128 4165
rect 44364 4199 44416 4208
rect 44364 4165 44373 4199
rect 44373 4165 44407 4199
rect 44407 4165 44416 4199
rect 44364 4156 44416 4165
rect 38936 4088 38988 4140
rect 33140 4020 33192 4072
rect 34704 4020 34756 4072
rect 36360 4020 36412 4072
rect 39120 4020 39172 4072
rect 34612 3952 34664 4004
rect 42892 4131 42944 4140
rect 42892 4097 42901 4131
rect 42901 4097 42935 4131
rect 42935 4097 42944 4131
rect 42892 4088 42944 4097
rect 46848 4156 46900 4208
rect 42984 4020 43036 4072
rect 43352 4020 43404 4072
rect 44640 4063 44692 4072
rect 44640 4029 44649 4063
rect 44649 4029 44683 4063
rect 44683 4029 44692 4063
rect 44640 4020 44692 4029
rect 33968 3884 34020 3936
rect 42616 3927 42668 3936
rect 42616 3893 42625 3927
rect 42625 3893 42659 3927
rect 42659 3893 42668 3927
rect 42616 3884 42668 3893
rect 43260 3884 43312 3936
rect 54852 4088 54904 4140
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 4620 3680 4672 3732
rect 4896 3680 4948 3732
rect 940 3612 992 3664
rect 4068 3612 4120 3664
rect 5816 3612 5868 3664
rect 10692 3680 10744 3732
rect 12072 3680 12124 3732
rect 12440 3680 12492 3732
rect 13176 3680 13228 3732
rect 17316 3680 17368 3732
rect 18052 3680 18104 3732
rect 20168 3680 20220 3732
rect 28724 3680 28776 3732
rect 30932 3680 30984 3732
rect 31392 3680 31444 3732
rect 40040 3680 40092 3732
rect 43352 3680 43404 3732
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 3700 3476 3752 3528
rect 5172 3544 5224 3596
rect 6460 3544 6512 3596
rect 10416 3612 10468 3664
rect 12164 3612 12216 3664
rect 13360 3612 13412 3664
rect 16120 3612 16172 3664
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 4988 3476 5040 3528
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 1032 3408 1084 3460
rect 3608 3408 3660 3460
rect 4068 3408 4120 3460
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 9128 3476 9180 3528
rect 11520 3544 11572 3596
rect 11796 3544 11848 3596
rect 11888 3544 11940 3596
rect 6000 3408 6052 3460
rect 9404 3408 9456 3460
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 5816 3383 5868 3392
rect 5816 3349 5825 3383
rect 5825 3349 5859 3383
rect 5859 3349 5868 3383
rect 5816 3340 5868 3349
rect 11520 3408 11572 3460
rect 11796 3408 11848 3460
rect 12808 3476 12860 3528
rect 13176 3519 13228 3528
rect 13176 3485 13186 3519
rect 13186 3485 13220 3519
rect 13220 3485 13228 3519
rect 13176 3476 13228 3485
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13544 3476 13596 3528
rect 13636 3340 13688 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 14280 3408 14332 3460
rect 16304 3519 16356 3528
rect 16304 3485 16314 3519
rect 16314 3485 16348 3519
rect 16348 3485 16356 3519
rect 16580 3519 16632 3528
rect 16304 3476 16356 3485
rect 16580 3485 16597 3519
rect 16597 3485 16631 3519
rect 16631 3485 16632 3519
rect 16580 3476 16632 3485
rect 16764 3476 16816 3528
rect 17408 3519 17460 3528
rect 17408 3485 17418 3519
rect 17418 3485 17452 3519
rect 17452 3485 17460 3519
rect 17408 3476 17460 3485
rect 17868 3476 17920 3528
rect 16120 3408 16172 3460
rect 18972 3476 19024 3528
rect 19432 3476 19484 3528
rect 20812 3612 20864 3664
rect 27160 3655 27212 3664
rect 27160 3621 27169 3655
rect 27169 3621 27203 3655
rect 27203 3621 27212 3655
rect 27160 3612 27212 3621
rect 28908 3612 28960 3664
rect 20628 3544 20680 3596
rect 20536 3519 20588 3528
rect 20536 3485 20546 3519
rect 20546 3485 20580 3519
rect 20580 3485 20588 3519
rect 20536 3476 20588 3485
rect 22192 3544 22244 3596
rect 27620 3587 27672 3596
rect 27620 3553 27629 3587
rect 27629 3553 27663 3587
rect 27663 3553 27672 3587
rect 27620 3544 27672 3553
rect 30104 3612 30156 3664
rect 21088 3476 21140 3528
rect 23664 3476 23716 3528
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 25872 3476 25924 3528
rect 29460 3544 29512 3596
rect 28540 3519 28592 3528
rect 28540 3485 28549 3519
rect 28549 3485 28583 3519
rect 28583 3485 28592 3519
rect 28540 3476 28592 3485
rect 16764 3340 16816 3392
rect 19340 3408 19392 3460
rect 20996 3340 21048 3392
rect 21272 3340 21324 3392
rect 21640 3408 21692 3460
rect 22560 3408 22612 3460
rect 23848 3408 23900 3460
rect 23572 3383 23624 3392
rect 23572 3349 23581 3383
rect 23581 3349 23615 3383
rect 23615 3349 23624 3383
rect 23572 3340 23624 3349
rect 25412 3340 25464 3392
rect 28908 3519 28960 3528
rect 28908 3485 28917 3519
rect 28917 3485 28951 3519
rect 28951 3485 28960 3519
rect 28908 3476 28960 3485
rect 29920 3408 29972 3460
rect 30288 3408 30340 3460
rect 30012 3340 30064 3392
rect 30564 3476 30616 3528
rect 30748 3519 30800 3528
rect 30748 3485 30757 3519
rect 30757 3485 30791 3519
rect 30791 3485 30800 3519
rect 30748 3476 30800 3485
rect 30932 3519 30984 3528
rect 30932 3485 30941 3519
rect 30941 3485 30975 3519
rect 30975 3485 30984 3519
rect 30932 3476 30984 3485
rect 31484 3612 31536 3664
rect 40500 3612 40552 3664
rect 31944 3587 31996 3596
rect 31944 3553 31953 3587
rect 31953 3553 31987 3587
rect 31987 3553 31996 3587
rect 31944 3544 31996 3553
rect 33876 3544 33928 3596
rect 35900 3587 35952 3596
rect 35900 3553 35909 3587
rect 35909 3553 35943 3587
rect 35943 3553 35952 3587
rect 35900 3544 35952 3553
rect 30472 3408 30524 3460
rect 31392 3476 31444 3528
rect 31208 3408 31260 3460
rect 31760 3340 31812 3392
rect 32036 3340 32088 3392
rect 35532 3476 35584 3528
rect 38200 3476 38252 3528
rect 38752 3476 38804 3528
rect 41052 3519 41104 3528
rect 41052 3485 41061 3519
rect 41061 3485 41095 3519
rect 41095 3485 41104 3519
rect 41052 3476 41104 3485
rect 42616 3476 42668 3528
rect 44364 3476 44416 3528
rect 35348 3408 35400 3460
rect 40040 3408 40092 3460
rect 57060 3408 57112 3460
rect 34704 3340 34756 3392
rect 37280 3383 37332 3392
rect 37280 3349 37289 3383
rect 37289 3349 37323 3383
rect 37323 3349 37332 3383
rect 37280 3340 37332 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4896 3136 4948 3188
rect 5816 3136 5868 3188
rect 9772 3136 9824 3188
rect 9956 3136 10008 3188
rect 1860 3068 1912 3120
rect 6368 3068 6420 3120
rect 2228 3000 2280 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4436 3000 4488 3052
rect 5264 3000 5316 3052
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 8392 3068 8444 3120
rect 8668 3068 8720 3120
rect 10048 3111 10100 3120
rect 10048 3077 10057 3111
rect 10057 3077 10091 3111
rect 10091 3077 10100 3111
rect 10048 3068 10100 3077
rect 10784 3068 10836 3120
rect 5632 3000 5684 3009
rect 940 2932 992 2984
rect 3240 2932 3292 2984
rect 5816 2907 5868 2916
rect 5816 2873 5825 2907
rect 5825 2873 5859 2907
rect 5859 2873 5868 2907
rect 5816 2864 5868 2873
rect 8760 3000 8812 3052
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 13636 3068 13688 3120
rect 10968 3000 11020 3009
rect 13452 3000 13504 3052
rect 14648 3068 14700 3120
rect 19984 3068 20036 3120
rect 21548 3136 21600 3188
rect 23848 3136 23900 3188
rect 23940 3179 23992 3188
rect 23940 3145 23949 3179
rect 23949 3145 23983 3179
rect 23983 3145 23992 3179
rect 23940 3136 23992 3145
rect 26148 3136 26200 3188
rect 27804 3136 27856 3188
rect 29000 3136 29052 3188
rect 30012 3136 30064 3188
rect 30472 3136 30524 3188
rect 35716 3136 35768 3188
rect 39120 3136 39172 3188
rect 41236 3136 41288 3188
rect 43168 3136 43220 3188
rect 44456 3179 44508 3188
rect 44456 3145 44465 3179
rect 44465 3145 44499 3179
rect 44499 3145 44508 3179
rect 44456 3136 44508 3145
rect 44916 3136 44968 3188
rect 47952 3179 48004 3188
rect 47952 3145 47961 3179
rect 47961 3145 47995 3179
rect 47995 3145 48004 3179
rect 47952 3136 48004 3145
rect 54116 3179 54168 3188
rect 54116 3145 54125 3179
rect 54125 3145 54159 3179
rect 54159 3145 54168 3179
rect 54116 3136 54168 3145
rect 55956 3179 56008 3188
rect 55956 3145 55965 3179
rect 55965 3145 55999 3179
rect 55999 3145 56008 3179
rect 55956 3136 56008 3145
rect 6920 2932 6972 2984
rect 8484 2932 8536 2984
rect 9220 2864 9272 2916
rect 11244 2932 11296 2984
rect 12900 2932 12952 2984
rect 15660 2932 15712 2984
rect 13912 2864 13964 2916
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 17500 2932 17552 2984
rect 18420 2932 18472 2984
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 20904 3043 20956 3052
rect 20904 3009 20914 3043
rect 20914 3009 20948 3043
rect 20948 3009 20956 3043
rect 20904 3000 20956 3009
rect 20996 3000 21048 3052
rect 9772 2796 9824 2848
rect 15200 2796 15252 2848
rect 15292 2839 15344 2848
rect 15292 2805 15301 2839
rect 15301 2805 15335 2839
rect 15335 2805 15344 2839
rect 15292 2796 15344 2805
rect 17960 2796 18012 2848
rect 20536 2796 20588 2848
rect 22192 3000 22244 3052
rect 25872 3068 25924 3120
rect 23572 3000 23624 3052
rect 24952 3043 25004 3052
rect 24952 3009 24961 3043
rect 24961 3009 24995 3043
rect 24995 3009 25004 3043
rect 24952 3000 25004 3009
rect 27528 3000 27580 3052
rect 32588 3111 32640 3120
rect 32588 3077 32597 3111
rect 32597 3077 32631 3111
rect 32631 3077 32640 3111
rect 32588 3068 32640 3077
rect 33508 3068 33560 3120
rect 35900 3068 35952 3120
rect 30564 3043 30616 3052
rect 30564 3009 30573 3043
rect 30573 3009 30607 3043
rect 30607 3009 30616 3043
rect 30564 3000 30616 3009
rect 30748 3041 30800 3050
rect 30748 3007 30757 3041
rect 30757 3007 30791 3041
rect 30791 3007 30800 3041
rect 30748 2998 30800 3007
rect 24860 2932 24912 2984
rect 25872 2932 25924 2984
rect 31208 3000 31260 3052
rect 31760 3000 31812 3052
rect 33140 3000 33192 3052
rect 33876 3043 33928 3052
rect 33876 3009 33885 3043
rect 33885 3009 33919 3043
rect 33919 3009 33928 3043
rect 33876 3000 33928 3009
rect 33968 3000 34020 3052
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 38200 3043 38252 3052
rect 38200 3009 38209 3043
rect 38209 3009 38243 3043
rect 38243 3009 38252 3043
rect 38200 3000 38252 3009
rect 38292 3000 38344 3052
rect 41052 3068 41104 3120
rect 41512 3068 41564 3120
rect 45284 3068 45336 3120
rect 41420 3000 41472 3052
rect 42800 3000 42852 3052
rect 44180 3000 44232 3052
rect 45560 3000 45612 3052
rect 46940 3000 46992 3052
rect 56968 3111 57020 3120
rect 56968 3077 56977 3111
rect 56977 3077 57011 3111
rect 57011 3077 57020 3111
rect 56968 3068 57020 3077
rect 49700 3000 49752 3052
rect 51632 3043 51684 3052
rect 51632 3009 51641 3043
rect 51641 3009 51675 3043
rect 51675 3009 51684 3043
rect 51632 3000 51684 3009
rect 53840 3000 53892 3052
rect 54852 3043 54904 3052
rect 54852 3009 54861 3043
rect 54861 3009 54895 3043
rect 54895 3009 54904 3043
rect 54852 3000 54904 3009
rect 30748 2864 30800 2916
rect 31484 2932 31536 2984
rect 36360 2932 36412 2984
rect 48780 2932 48832 2984
rect 50160 2932 50212 2984
rect 51540 2932 51592 2984
rect 54300 2932 54352 2984
rect 56600 3000 56652 3052
rect 57980 2932 58032 2984
rect 24952 2796 25004 2848
rect 40224 2796 40276 2848
rect 44364 2864 44416 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 5448 2456 5500 2508
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 7104 2388 7156 2440
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 15292 2524 15344 2576
rect 2780 2320 2832 2372
rect 4068 2320 4120 2372
rect 4620 2320 4672 2372
rect 5080 2320 5132 2372
rect 7380 2320 7432 2372
rect 7840 2320 7892 2372
rect 10140 2320 10192 2372
rect 10600 2320 10652 2372
rect 3424 2252 3476 2304
rect 8576 2252 8628 2304
rect 9220 2252 9272 2304
rect 11980 2252 12032 2304
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 12440 2320 12492 2372
rect 13360 2320 13412 2372
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 17408 2388 17460 2440
rect 15200 2363 15252 2372
rect 15200 2329 15209 2363
rect 15209 2329 15243 2363
rect 15243 2329 15252 2363
rect 15200 2320 15252 2329
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 17868 2320 17920 2372
rect 21824 2524 21876 2576
rect 24768 2524 24820 2576
rect 24952 2524 25004 2576
rect 22468 2456 22520 2508
rect 18696 2363 18748 2372
rect 18696 2329 18705 2363
rect 18705 2329 18739 2363
rect 18739 2329 18748 2363
rect 18696 2320 18748 2329
rect 14740 2252 14792 2304
rect 22100 2388 22152 2440
rect 25136 2456 25188 2508
rect 20628 2320 20680 2372
rect 22008 2320 22060 2372
rect 23020 2320 23072 2372
rect 23480 2252 23532 2304
rect 23940 2388 23992 2440
rect 32312 2592 32364 2644
rect 33508 2592 33560 2644
rect 34244 2592 34296 2644
rect 35532 2635 35584 2644
rect 35532 2601 35541 2635
rect 35541 2601 35575 2635
rect 35575 2601 35584 2635
rect 35532 2592 35584 2601
rect 36912 2592 36964 2644
rect 40316 2592 40368 2644
rect 27436 2524 27488 2576
rect 30196 2524 30248 2576
rect 53104 2635 53156 2644
rect 53104 2601 53113 2635
rect 53113 2601 53147 2635
rect 53147 2601 53156 2635
rect 53104 2592 53156 2601
rect 24400 2320 24452 2372
rect 25320 2320 25372 2372
rect 26240 2320 26292 2372
rect 26700 2320 26752 2372
rect 26332 2252 26384 2304
rect 28264 2388 28316 2440
rect 29644 2388 29696 2440
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 28080 2320 28132 2372
rect 29460 2320 29512 2372
rect 30840 2320 30892 2372
rect 33508 2456 33560 2508
rect 33600 2456 33652 2508
rect 37280 2456 37332 2508
rect 42432 2456 42484 2508
rect 33692 2431 33744 2440
rect 33692 2397 33701 2431
rect 33701 2397 33735 2431
rect 33735 2397 33744 2431
rect 33692 2388 33744 2397
rect 34612 2388 34664 2440
rect 34980 2431 35032 2440
rect 34980 2397 34990 2431
rect 34990 2397 35024 2431
rect 35024 2397 35032 2431
rect 34980 2388 35032 2397
rect 35256 2431 35308 2440
rect 35256 2397 35265 2431
rect 35265 2397 35299 2431
rect 35299 2397 35308 2431
rect 35256 2388 35308 2397
rect 32220 2320 32272 2372
rect 33600 2320 33652 2372
rect 34060 2320 34112 2372
rect 32036 2252 32088 2304
rect 35624 2388 35676 2440
rect 37832 2431 37884 2440
rect 37832 2397 37841 2431
rect 37841 2397 37875 2431
rect 37875 2397 37884 2431
rect 37832 2388 37884 2397
rect 39212 2388 39264 2440
rect 40960 2431 41012 2440
rect 40960 2397 40969 2431
rect 40969 2397 41003 2431
rect 41003 2397 41012 2431
rect 40960 2388 41012 2397
rect 42524 2388 42576 2440
rect 43444 2388 43496 2440
rect 43812 2456 43864 2508
rect 36268 2363 36320 2372
rect 36268 2329 36277 2363
rect 36277 2329 36311 2363
rect 36311 2329 36320 2363
rect 36268 2320 36320 2329
rect 37740 2320 37792 2372
rect 38844 2363 38896 2372
rect 38844 2329 38853 2363
rect 38853 2329 38887 2363
rect 38887 2329 38896 2363
rect 38844 2320 38896 2329
rect 40316 2363 40368 2372
rect 40316 2329 40325 2363
rect 40325 2329 40359 2363
rect 40359 2329 40368 2363
rect 40316 2320 40368 2329
rect 40500 2320 40552 2372
rect 42892 2363 42944 2372
rect 42892 2329 42901 2363
rect 42901 2329 42935 2363
rect 42935 2329 42944 2363
rect 42892 2320 42944 2329
rect 43260 2320 43312 2372
rect 44640 2320 44692 2372
rect 46020 2320 46072 2372
rect 44272 2252 44324 2304
rect 55220 2388 55272 2440
rect 56416 2431 56468 2440
rect 56416 2397 56425 2431
rect 56425 2397 56459 2431
rect 56459 2397 56468 2431
rect 56416 2388 56468 2397
rect 47400 2320 47452 2372
rect 48320 2320 48372 2372
rect 49700 2320 49752 2372
rect 51080 2320 51132 2372
rect 52460 2320 52512 2372
rect 54116 2363 54168 2372
rect 54116 2329 54125 2363
rect 54125 2329 54159 2363
rect 54159 2329 54168 2363
rect 54116 2320 54168 2329
rect 55772 2363 55824 2372
rect 55772 2329 55781 2363
rect 55781 2329 55815 2363
rect 55815 2329 55824 2363
rect 55772 2320 55824 2329
rect 56692 2363 56744 2372
rect 56692 2329 56701 2363
rect 56701 2329 56735 2363
rect 56735 2329 56744 2363
rect 56692 2320 56744 2329
rect 48872 2295 48924 2304
rect 48872 2261 48881 2295
rect 48881 2261 48915 2295
rect 48915 2261 48924 2295
rect 48872 2252 48924 2261
rect 51448 2295 51500 2304
rect 51448 2261 51457 2295
rect 51457 2261 51491 2295
rect 51491 2261 51500 2295
rect 51448 2252 51500 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 22468 2048 22520 2100
rect 30472 2048 30524 2100
rect 2872 1980 2924 2032
rect 4804 1980 4856 2032
rect 5172 1980 5224 2032
rect 11336 1980 11388 2032
rect 12992 1980 13044 2032
rect 48872 1980 48924 2032
rect 2964 1912 3016 1964
rect 11152 1912 11204 1964
rect 15844 1912 15896 1964
rect 2044 1844 2096 1896
rect 11704 1844 11756 1896
rect 23480 1912 23532 1964
rect 27160 1912 27212 1964
rect 46848 1912 46900 1964
rect 56416 1912 56468 1964
rect 30748 1844 30800 1896
rect 35256 1844 35308 1896
rect 6092 1776 6144 1828
rect 51448 1776 51500 1828
rect 13268 1708 13320 1760
rect 31392 1708 31444 1760
rect 8852 1640 8904 1692
rect 55772 1640 55824 1692
rect 3332 1300 3384 1352
rect 21916 1300 21968 1352
rect 18696 892 18748 944
rect 19800 892 19852 944
rect 34980 892 35032 944
rect 36268 892 36320 944
rect 37280 892 37332 944
rect 38844 892 38896 944
rect 39120 892 39172 944
rect 40316 892 40368 944
rect 41880 892 41932 944
rect 42892 892 42944 944
rect 52920 892 52972 944
rect 54116 892 54168 944
rect 55680 892 55732 944
rect 56692 892 56744 944
<< metal2 >>
rect 3882 41200 3938 42000
rect 11334 41200 11390 42000
rect 18786 41200 18842 42000
rect 26238 41200 26294 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48594 41200 48650 42000
rect 56046 41200 56102 42000
rect 1122 41168 1178 41177
rect 3896 41138 3924 41200
rect 18800 41138 18828 41200
rect 1122 41103 1178 41112
rect 3884 41132 3936 41138
rect 1030 40352 1086 40361
rect 1030 40287 1086 40296
rect 938 39536 994 39545
rect 938 39471 940 39480
rect 992 39471 994 39480
rect 940 39442 992 39448
rect 1044 39370 1072 40287
rect 1032 39364 1084 39370
rect 1032 39306 1084 39312
rect 940 38888 992 38894
rect 940 38830 992 38836
rect 952 38729 980 38830
rect 1136 38826 1164 41103
rect 3884 41074 3936 41080
rect 4620 41132 4672 41138
rect 4620 41074 4672 41080
rect 18788 41132 18840 41138
rect 18788 41074 18840 41080
rect 19432 41132 19484 41138
rect 19432 41074 19484 41080
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4632 39506 4660 41074
rect 19444 39506 19472 41074
rect 26252 39506 26280 41200
rect 3424 39500 3476 39506
rect 3424 39442 3476 39448
rect 4620 39500 4672 39506
rect 4620 39442 4672 39448
rect 19432 39500 19484 39506
rect 19432 39442 19484 39448
rect 26240 39500 26292 39506
rect 26240 39442 26292 39448
rect 2504 39432 2556 39438
rect 2504 39374 2556 39380
rect 1124 38820 1176 38826
rect 1124 38762 1176 38768
rect 938 38720 994 38729
rect 938 38655 994 38664
rect 940 38276 992 38282
rect 940 38218 992 38224
rect 952 37913 980 38218
rect 938 37904 994 37913
rect 938 37839 994 37848
rect 2516 37670 2544 39374
rect 2504 37664 2556 37670
rect 2504 37606 2556 37612
rect 3436 37466 3464 39442
rect 33704 39438 33732 41200
rect 41156 41154 41184 41200
rect 41156 41126 41460 41154
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 41432 39642 41460 41126
rect 48608 39642 48636 41200
rect 41420 39636 41472 39642
rect 41420 39578 41472 39584
rect 48596 39636 48648 39642
rect 48596 39578 48648 39584
rect 56060 39506 56088 41200
rect 56048 39500 56100 39506
rect 56048 39442 56100 39448
rect 27160 39432 27212 39438
rect 27160 39374 27212 39380
rect 33692 39432 33744 39438
rect 33692 39374 33744 39380
rect 42156 39432 42208 39438
rect 42156 39374 42208 39380
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 7656 39024 7708 39030
rect 7656 38966 7708 38972
rect 6184 38956 6236 38962
rect 6184 38898 6236 38904
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 6196 37942 6224 38898
rect 6184 37936 6236 37942
rect 6184 37878 6236 37884
rect 6000 37664 6052 37670
rect 6000 37606 6052 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3424 37460 3476 37466
rect 3424 37402 3476 37408
rect 5356 37460 5408 37466
rect 5356 37402 5408 37408
rect 4068 37256 4120 37262
rect 4068 37198 4120 37204
rect 940 37188 992 37194
rect 940 37130 992 37136
rect 952 37097 980 37130
rect 938 37088 994 37097
rect 938 37023 994 37032
rect 940 36712 992 36718
rect 940 36654 992 36660
rect 952 36281 980 36654
rect 938 36272 994 36281
rect 938 36207 994 36216
rect 940 35624 992 35630
rect 940 35566 992 35572
rect 952 35465 980 35566
rect 938 35456 994 35465
rect 938 35391 994 35400
rect 940 35012 992 35018
rect 940 34954 992 34960
rect 952 34649 980 34954
rect 938 34640 994 34649
rect 938 34575 994 34584
rect 1032 34604 1084 34610
rect 1032 34546 1084 34552
rect 940 34536 992 34542
rect 940 34478 992 34484
rect 952 34241 980 34478
rect 938 34232 994 34241
rect 938 34167 994 34176
rect 1044 33833 1072 34546
rect 2688 34536 2740 34542
rect 2688 34478 2740 34484
rect 1124 33924 1176 33930
rect 1124 33866 1176 33872
rect 2136 33924 2188 33930
rect 2136 33866 2188 33872
rect 1030 33824 1086 33833
rect 1030 33759 1086 33768
rect 940 33448 992 33454
rect 938 33416 940 33425
rect 992 33416 994 33425
rect 938 33351 994 33360
rect 1136 33017 1164 33866
rect 1122 33008 1178 33017
rect 1122 32943 1178 32952
rect 940 32836 992 32842
rect 940 32778 992 32784
rect 952 32609 980 32778
rect 938 32600 994 32609
rect 938 32535 994 32544
rect 940 32360 992 32366
rect 940 32302 992 32308
rect 952 32201 980 32302
rect 938 32192 994 32201
rect 938 32127 994 32136
rect 1032 31884 1084 31890
rect 1032 31826 1084 31832
rect 940 31816 992 31822
rect 1044 31793 1072 31826
rect 940 31758 992 31764
rect 1030 31784 1086 31793
rect 952 31385 980 31758
rect 1030 31719 1086 31728
rect 938 31376 994 31385
rect 938 31311 994 31320
rect 940 31272 992 31278
rect 940 31214 992 31220
rect 952 30977 980 31214
rect 938 30968 994 30977
rect 938 30903 994 30912
rect 940 30660 992 30666
rect 940 30602 992 30608
rect 952 30569 980 30602
rect 1860 30592 1912 30598
rect 938 30560 994 30569
rect 1860 30534 1912 30540
rect 938 30495 994 30504
rect 940 30184 992 30190
rect 940 30126 992 30132
rect 1030 30152 1086 30161
rect 952 29753 980 30126
rect 1030 30087 1032 30096
rect 1084 30087 1086 30096
rect 1032 30058 1084 30064
rect 938 29744 994 29753
rect 938 29679 994 29688
rect 940 29572 992 29578
rect 940 29514 992 29520
rect 952 29345 980 29514
rect 938 29336 994 29345
rect 938 29271 994 29280
rect 1032 29096 1084 29102
rect 1032 29038 1084 29044
rect 940 29028 992 29034
rect 940 28970 992 28976
rect 952 28937 980 28970
rect 938 28928 994 28937
rect 938 28863 994 28872
rect 1044 28529 1072 29038
rect 1030 28520 1086 28529
rect 940 28484 992 28490
rect 1030 28455 1086 28464
rect 940 28426 992 28432
rect 952 28121 980 28426
rect 938 28112 994 28121
rect 938 28047 994 28056
rect 940 28008 992 28014
rect 940 27950 992 27956
rect 952 27713 980 27950
rect 1032 27940 1084 27946
rect 1032 27882 1084 27888
rect 938 27704 994 27713
rect 938 27639 994 27648
rect 940 27396 992 27402
rect 940 27338 992 27344
rect 952 26897 980 27338
rect 1044 27305 1072 27882
rect 1030 27296 1086 27305
rect 1030 27231 1086 27240
rect 1032 27056 1084 27062
rect 1032 26998 1084 27004
rect 938 26888 994 26897
rect 938 26823 994 26832
rect 1044 26489 1072 26998
rect 1124 26920 1176 26926
rect 1124 26862 1176 26868
rect 1030 26480 1086 26489
rect 1030 26415 1086 26424
rect 940 26308 992 26314
rect 940 26250 992 26256
rect 952 25673 980 26250
rect 1136 26081 1164 26862
rect 1122 26072 1178 26081
rect 1122 26007 1178 26016
rect 1124 25968 1176 25974
rect 1124 25910 1176 25916
rect 1032 25832 1084 25838
rect 1032 25774 1084 25780
rect 938 25664 994 25673
rect 938 25599 994 25608
rect 1044 24857 1072 25774
rect 1136 25265 1164 25910
rect 1122 25256 1178 25265
rect 1122 25191 1178 25200
rect 1030 24848 1086 24857
rect 940 24812 992 24818
rect 1030 24783 1086 24792
rect 940 24754 992 24760
rect 952 24449 980 24754
rect 1032 24744 1084 24750
rect 1032 24686 1084 24692
rect 938 24440 994 24449
rect 938 24375 994 24384
rect 1044 24041 1072 24686
rect 1676 24200 1728 24206
rect 1676 24142 1728 24148
rect 1030 24032 1086 24041
rect 1030 23967 1086 23976
rect 940 23724 992 23730
rect 940 23666 992 23672
rect 952 23225 980 23666
rect 1030 23624 1086 23633
rect 1030 23559 1086 23568
rect 938 23216 994 23225
rect 1044 23186 1072 23559
rect 938 23151 994 23160
rect 1032 23180 1084 23186
rect 1032 23122 1084 23128
rect 940 22976 992 22982
rect 940 22918 992 22924
rect 952 22817 980 22918
rect 938 22808 994 22817
rect 938 22743 994 22752
rect 1030 22400 1086 22409
rect 1030 22335 1086 22344
rect 938 21992 994 22001
rect 938 21927 940 21936
rect 992 21927 994 21936
rect 940 21898 992 21904
rect 940 21684 992 21690
rect 940 21626 992 21632
rect 952 21593 980 21626
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 1044 21486 1072 22335
rect 1688 22030 1716 24142
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 1032 21480 1084 21486
rect 1032 21422 1084 21428
rect 940 21412 992 21418
rect 940 21354 992 21360
rect 952 21185 980 21354
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 1688 20942 1716 21966
rect 1872 21350 1900 30534
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 1964 27130 1992 27270
rect 1952 27124 2004 27130
rect 1952 27066 2004 27072
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 2056 24750 2084 25230
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 1952 24404 2004 24410
rect 1952 24346 2004 24352
rect 1964 23866 1992 24346
rect 2056 24206 2084 24686
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 1964 22030 1992 22374
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1030 20768 1086 20777
rect 1030 20703 1086 20712
rect 940 20392 992 20398
rect 938 20360 940 20369
rect 992 20360 994 20369
rect 938 20295 994 20304
rect 938 19952 994 19961
rect 938 19887 940 19896
rect 992 19887 994 19896
rect 940 19858 992 19864
rect 1044 19854 1072 20703
rect 1688 20466 1716 20878
rect 2148 20602 2176 33866
rect 2504 32836 2556 32842
rect 2504 32778 2556 32784
rect 2412 29572 2464 29578
rect 2412 29514 2464 29520
rect 2320 26240 2372 26246
rect 2320 26182 2372 26188
rect 2332 25294 2360 26182
rect 2320 25288 2372 25294
rect 2320 25230 2372 25236
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 2240 21894 2268 24550
rect 2424 23338 2452 29514
rect 2516 26450 2544 32778
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2608 24614 2636 31758
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2516 23866 2544 24074
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2332 23310 2452 23338
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2240 20534 2268 20742
rect 2228 20528 2280 20534
rect 2228 20470 2280 20476
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 2332 20262 2360 23310
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2424 22778 2452 22918
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2608 21010 2636 22510
rect 2596 21004 2648 21010
rect 2596 20946 2648 20952
rect 2504 20528 2556 20534
rect 2504 20470 2556 20476
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2516 19854 2544 20470
rect 1032 19848 1084 19854
rect 1032 19790 1084 19796
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 940 19780 992 19786
rect 940 19722 992 19728
rect 952 19553 980 19722
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 938 19544 994 19553
rect 938 19479 994 19488
rect 940 19236 992 19242
rect 940 19178 992 19184
rect 952 19145 980 19178
rect 938 19136 994 19145
rect 938 19071 994 19080
rect 1768 18760 1820 18766
rect 938 18728 994 18737
rect 1768 18702 1820 18708
rect 938 18663 994 18672
rect 952 18358 980 18663
rect 1032 18420 1084 18426
rect 1032 18362 1084 18368
rect 940 18352 992 18358
rect 940 18294 992 18300
rect 1044 17921 1072 18362
rect 1122 18320 1178 18329
rect 1122 18255 1178 18264
rect 1030 17912 1086 17921
rect 1030 17847 1086 17856
rect 940 17672 992 17678
rect 940 17614 992 17620
rect 952 17513 980 17614
rect 1136 17610 1164 18255
rect 1780 17746 1808 18702
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1124 17604 1176 17610
rect 1124 17546 1176 17552
rect 938 17504 994 17513
rect 938 17439 994 17448
rect 940 17264 992 17270
rect 940 17206 992 17212
rect 952 17105 980 17206
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 938 16688 994 16697
rect 1780 16658 1808 17682
rect 938 16623 994 16632
rect 1768 16652 1820 16658
rect 952 16590 980 16623
rect 1768 16594 1820 16600
rect 940 16584 992 16590
rect 940 16526 992 16532
rect 938 16280 994 16289
rect 938 16215 994 16224
rect 952 16182 980 16215
rect 940 16176 992 16182
rect 1964 16153 1992 19654
rect 2700 19394 2728 34478
rect 4080 31958 4108 37198
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4620 34672 4672 34678
rect 4620 34614 4672 34620
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4068 31952 4120 31958
rect 4068 31894 4120 31900
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28490 4660 34614
rect 4620 28484 4672 28490
rect 4620 28426 4672 28432
rect 4068 28144 4120 28150
rect 4068 28086 4120 28092
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 2780 26852 2832 26858
rect 2780 26794 2832 26800
rect 2792 23866 2820 26794
rect 3424 26240 3476 26246
rect 3424 26182 3476 26188
rect 3436 25158 3464 26182
rect 3884 25696 3936 25702
rect 3884 25638 3936 25644
rect 3608 25288 3660 25294
rect 3608 25230 3660 25236
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2964 23656 3016 23662
rect 2964 23598 3016 23604
rect 2976 23186 3004 23598
rect 3436 23254 3464 25094
rect 3620 24750 3648 25230
rect 3896 24818 3924 25638
rect 3884 24812 3936 24818
rect 3884 24754 3936 24760
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3516 24676 3568 24682
rect 3516 24618 3568 24624
rect 3528 23866 3556 24618
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2976 22574 3004 23122
rect 3620 22642 3648 24686
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 3068 22234 3096 22578
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3252 21690 3280 22578
rect 3332 22432 3384 22438
rect 3332 22374 3384 22380
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3344 20874 3372 22374
rect 3988 21690 4016 26930
rect 4080 26926 4108 28086
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 4356 25838 4384 26386
rect 4632 26042 4660 27882
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 5276 26586 5304 26998
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 4988 25900 5040 25906
rect 4988 25842 5040 25848
rect 4344 25832 4396 25838
rect 4344 25774 4396 25780
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24206 4660 25706
rect 5000 24954 5028 25842
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4816 23662 4844 24006
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4436 22976 4488 22982
rect 4436 22918 4488 22924
rect 4448 22710 4476 22918
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4816 22098 4844 23598
rect 4908 22982 4936 24550
rect 5000 23798 5028 24890
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4804 22092 4856 22098
rect 4804 22034 4856 22040
rect 5000 21962 5028 23734
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 4988 21956 5040 21962
rect 4988 21898 5040 21904
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 5092 21554 5120 23462
rect 5184 23050 5212 23666
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5184 22778 5212 22986
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5184 22234 5212 22714
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3436 20806 3464 21422
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3436 20602 3464 20742
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 2976 20398 3004 20538
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3988 19514 4016 20198
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3240 19440 3292 19446
rect 2700 19366 2820 19394
rect 3240 19382 3292 19388
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 18766 2176 19110
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2424 16998 2452 17478
rect 2700 17134 2728 19246
rect 2792 18426 2820 19366
rect 3252 18970 3280 19382
rect 4080 18970 4108 21490
rect 5184 21350 5212 21966
rect 5276 21894 5304 21966
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2688 17128 2740 17134
rect 2608 17076 2688 17082
rect 2608 17070 2740 17076
rect 2608 17054 2728 17070
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2056 16658 2084 16934
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 940 16118 992 16124
rect 1950 16144 2006 16153
rect 1950 16079 2006 16088
rect 2608 16046 2636 17054
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 1122 15872 1178 15881
rect 1122 15807 1178 15816
rect 1030 15464 1086 15473
rect 940 15428 992 15434
rect 1030 15399 1086 15408
rect 940 15370 992 15376
rect 952 15065 980 15370
rect 1044 15366 1072 15399
rect 1032 15360 1084 15366
rect 1032 15302 1084 15308
rect 1136 15094 1164 15807
rect 1124 15088 1176 15094
rect 938 15056 994 15065
rect 1124 15030 1176 15036
rect 938 14991 994 15000
rect 938 14648 994 14657
rect 938 14583 994 14592
rect 952 14482 980 14583
rect 940 14476 992 14482
rect 940 14418 992 14424
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 940 14340 992 14346
rect 940 14282 992 14288
rect 952 13841 980 14282
rect 1030 14240 1086 14249
rect 1030 14175 1086 14184
rect 938 13832 994 13841
rect 938 13767 994 13776
rect 938 13424 994 13433
rect 938 13359 994 13368
rect 952 13258 980 13359
rect 940 13252 992 13258
rect 940 13194 992 13200
rect 938 13016 994 13025
rect 938 12951 940 12960
rect 992 12951 994 12960
rect 940 12922 992 12928
rect 1044 12918 1072 14175
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1964 13530 1992 13874
rect 2516 13530 2544 14350
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2608 13410 2636 13670
rect 2516 13394 2636 13410
rect 2516 13388 2648 13394
rect 2516 13382 2596 13388
rect 1032 12912 1084 12918
rect 1032 12854 1084 12860
rect 940 12776 992 12782
rect 940 12718 992 12724
rect 952 12617 980 12718
rect 938 12608 994 12617
rect 938 12543 994 12552
rect 940 12232 992 12238
rect 938 12200 940 12209
rect 992 12200 994 12209
rect 938 12135 994 12144
rect 1032 12164 1084 12170
rect 1032 12106 1084 12112
rect 1044 11801 1072 12106
rect 1124 11824 1176 11830
rect 1030 11792 1086 11801
rect 1124 11766 1176 11772
rect 1030 11727 1086 11736
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 952 11393 980 11630
rect 938 11384 994 11393
rect 938 11319 994 11328
rect 1136 10985 1164 11766
rect 2516 11694 2544 13382
rect 2596 13330 2648 13336
rect 2700 13274 2728 16934
rect 2792 16250 2820 18090
rect 3436 17338 3464 18294
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15094 3004 15846
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2608 13246 2728 13274
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1122 10976 1178 10985
rect 1122 10911 1178 10920
rect 1964 10810 1992 11018
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 940 10600 992 10606
rect 938 10568 940 10577
rect 992 10568 994 10577
rect 938 10503 994 10512
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 952 9761 980 9930
rect 938 9752 994 9761
rect 938 9687 994 9696
rect 1030 9344 1086 9353
rect 1030 9279 1086 9288
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 1044 8906 1072 9279
rect 1124 9036 1176 9042
rect 1124 8978 1176 8984
rect 938 8871 994 8880
rect 1032 8900 1084 8906
rect 1032 8842 1084 8848
rect 1032 8560 1084 8566
rect 1136 8537 1164 8978
rect 1032 8502 1084 8508
rect 1122 8528 1178 8537
rect 940 8424 992 8430
rect 940 8366 992 8372
rect 952 8129 980 8366
rect 938 8120 994 8129
rect 938 8055 994 8064
rect 1044 7721 1072 8502
rect 1122 8463 1178 8472
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1030 7712 1086 7721
rect 1030 7647 1086 7656
rect 940 7472 992 7478
rect 940 7414 992 7420
rect 952 7313 980 7414
rect 938 7304 994 7313
rect 938 7239 994 7248
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 952 6798 980 6831
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 938 6488 994 6497
rect 938 6423 994 6432
rect 952 5778 980 6423
rect 1780 6254 1808 7822
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7546 1992 7754
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6390 2176 6598
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1584 6112 1636 6118
rect 1030 6080 1086 6089
rect 1584 6054 1636 6060
rect 1030 6015 1086 6024
rect 940 5772 992 5778
rect 940 5714 992 5720
rect 940 5296 992 5302
rect 938 5264 940 5273
rect 992 5264 994 5273
rect 938 5199 994 5208
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4865 980 5102
rect 1044 5098 1072 6015
rect 1596 5710 1624 6054
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1032 5092 1084 5098
rect 1032 5034 1084 5040
rect 938 4856 994 4865
rect 1596 4826 1624 5170
rect 938 4791 994 4800
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1780 4622 1808 6190
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 938 4448 994 4457
rect 938 4383 994 4392
rect 952 4078 980 4383
rect 940 4072 992 4078
rect 940 4014 992 4020
rect 1124 4004 1176 4010
rect 1124 3946 1176 3952
rect 940 3664 992 3670
rect 938 3632 940 3641
rect 992 3632 994 3641
rect 938 3567 994 3576
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 940 2984 992 2990
rect 940 2926 992 2932
rect 952 2825 980 2926
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 1044 2417 1072 3402
rect 1030 2408 1086 2417
rect 1030 2343 1086 2352
rect 1136 785 1164 3946
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1964 3738 1992 3878
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1872 800 1900 3062
rect 2240 3058 2268 11494
rect 2516 10826 2544 11630
rect 2424 10798 2544 10826
rect 2424 10538 2452 10798
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2424 10010 2452 10474
rect 2332 9982 2452 10010
rect 2332 8242 2360 9982
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9586 2452 9862
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2516 9178 2544 10678
rect 2608 10198 2636 13246
rect 3068 13190 3096 13670
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 3068 12714 3096 13126
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2700 10538 2728 12038
rect 2792 11830 2820 12242
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3068 11286 3096 11766
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3068 10810 3096 11222
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2976 10130 3004 10406
rect 3068 10130 3096 10542
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9382 2912 9862
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 3252 9178 3280 17002
rect 3436 16590 3464 17274
rect 4540 17202 4568 17274
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 14822 4108 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3988 14482 4016 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 12782 3372 13126
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3804 12442 3832 14282
rect 3988 14006 4016 14418
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 14074 4108 14350
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3988 12238 4016 13942
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4080 12986 4108 13194
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11898 3464 12038
rect 3896 11898 3924 12106
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11286 3740 11698
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3896 9382 3924 11154
rect 3988 11150 4016 12174
rect 4344 12096 4396 12102
rect 4264 12056 4344 12084
rect 4264 11762 4292 12056
rect 4344 12038 4396 12044
rect 4632 11801 4660 19722
rect 4724 19310 4752 20334
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5184 17882 5212 18702
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5184 17678 5212 17818
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4988 17604 5040 17610
rect 4988 17546 5040 17552
rect 5000 17338 5028 17546
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4618 11792 4674 11801
rect 4252 11756 4304 11762
rect 4618 11727 4674 11736
rect 4252 11698 4304 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4080 10198 4108 10474
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4632 9586 4660 10474
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 2332 8214 2452 8242
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2332 7546 2360 8026
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2424 7342 2452 8214
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7886 4660 9522
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4528 7812 4580 7818
rect 4528 7754 4580 7760
rect 4540 7546 4568 7754
rect 4724 7750 4752 17274
rect 5184 16658 5212 17614
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2608 6866 2636 7278
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4816 6866 4844 13874
rect 4908 11150 4936 14758
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5000 13530 5028 13738
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11354 5028 12038
rect 5276 11354 5304 19110
rect 5368 17882 5396 37402
rect 6012 35894 6040 37606
rect 7668 35894 7696 38966
rect 10324 38344 10376 38350
rect 10324 38286 10376 38292
rect 6012 35866 6132 35894
rect 7668 35866 7788 35894
rect 5540 35080 5592 35086
rect 5540 35022 5592 35028
rect 5552 32502 5580 35022
rect 5540 32496 5592 32502
rect 5540 32438 5592 32444
rect 6000 26240 6052 26246
rect 6000 26182 6052 26188
rect 6012 25226 6040 26182
rect 6000 25220 6052 25226
rect 6000 25162 6052 25168
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5460 19854 5488 21286
rect 5552 19922 5580 21490
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5368 17134 5396 17818
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5460 16574 5488 19654
rect 5552 19446 5580 19858
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 6012 19514 6040 19790
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 5540 19440 5592 19446
rect 6104 19394 6132 35866
rect 6184 31952 6236 31958
rect 6184 31894 6236 31900
rect 6196 20262 6224 31894
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6460 29028 6512 29034
rect 6460 28970 6512 28976
rect 6472 26450 6500 28970
rect 6460 26444 6512 26450
rect 6460 26386 6512 26392
rect 6656 26382 6684 31826
rect 6644 26376 6696 26382
rect 6644 26318 6696 26324
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 6368 26240 6420 26246
rect 6368 26182 6420 26188
rect 7472 26240 7524 26246
rect 7472 26182 7524 26188
rect 6380 25498 6408 26182
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 6736 25696 6788 25702
rect 6736 25638 6788 25644
rect 6368 25492 6420 25498
rect 6368 25434 6420 25440
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6564 23730 6592 25230
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6564 23202 6592 23462
rect 6656 23322 6684 23666
rect 6644 23316 6696 23322
rect 6644 23258 6696 23264
rect 6564 23174 6684 23202
rect 6656 22982 6684 23174
rect 6748 23050 6776 25638
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7208 23322 7236 25434
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6472 19922 6500 21830
rect 6656 21350 6684 22918
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6644 20868 6696 20874
rect 6644 20810 6696 20816
rect 6656 20602 6684 20810
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 5540 19382 5592 19388
rect 6012 19366 6132 19394
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5644 16590 5672 17206
rect 5920 17066 5948 18634
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5920 16590 5948 17002
rect 6012 16590 6040 19366
rect 6196 18034 6224 19382
rect 6288 19378 6316 19654
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6380 18766 6408 19450
rect 6564 19378 6592 19994
rect 6656 19530 6684 20198
rect 6748 19854 6776 22374
rect 7208 21486 7236 23258
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6840 20262 6868 20402
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 7208 19718 7236 21286
rect 7300 20398 7328 23122
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 6656 19502 6776 19530
rect 6748 19446 6776 19502
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6748 18970 6776 19382
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6840 18834 6868 19314
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6104 18006 6224 18034
rect 5368 16546 5488 16574
rect 5632 16584 5684 16590
rect 5368 13326 5396 16546
rect 5632 16526 5684 16532
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5644 15638 5672 16526
rect 5828 16250 5856 16526
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5632 15632 5684 15638
rect 5632 15574 5684 15580
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 14414 5580 15370
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5644 14074 5672 14282
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5368 11830 5396 13262
rect 5920 12434 5948 13262
rect 5828 12406 5948 12434
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6458 2544 6598
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2608 5642 2636 6802
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5914 3464 6598
rect 3790 6352 3846 6361
rect 3790 6287 3792 6296
rect 3844 6287 3846 6296
rect 3792 6258 3844 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3436 5302 3464 5578
rect 3424 5296 3476 5302
rect 4172 5250 4200 5714
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 3424 5238 3476 5244
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4080 5222 4200 5250
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4826 3096 5102
rect 3896 5030 3924 5170
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 1902 2084 2382
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 2332 800 2360 4014
rect 2516 3534 2544 4558
rect 3068 4214 3096 4762
rect 3712 4554 3740 4966
rect 4080 4706 4108 5222
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3988 4678 4108 4706
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3988 4146 4016 4678
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 4282 4108 4490
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 3620 3466 3648 4082
rect 4080 3670 4108 4082
rect 4172 4078 4200 4422
rect 4264 4214 4292 4558
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3738 4660 5102
rect 4724 4146 4752 5510
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3620 3058 3648 3402
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2792 800 2820 2314
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 2884 1601 2912 1974
rect 2976 1970 3004 2382
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 3252 800 3280 2926
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 2009 3464 2246
rect 3422 2000 3478 2009
rect 3422 1935 3478 1944
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 1193 3372 1294
rect 3330 1184 3386 1193
rect 3330 1119 3386 1128
rect 3712 800 3740 3470
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 3233 4108 3402
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4066 3224 4122 3233
rect 4066 3159 4122 3168
rect 4448 3058 4476 3334
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4080 898 4108 2314
rect 4080 870 4200 898
rect 4172 800 4200 870
rect 4632 800 4660 2314
rect 4816 2038 4844 5578
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3738 4936 4082
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5000 3534 5028 11290
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5092 8090 5120 8366
rect 5184 8090 5212 8434
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5184 7546 5212 8026
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5092 3942 5120 5170
rect 5184 4690 5212 6054
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4078 5212 4626
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5184 3602 5212 4014
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4908 3194 4936 3470
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5276 3058 5304 11018
rect 5368 9058 5396 11154
rect 5552 10674 5580 11562
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5460 9178 5488 9522
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5368 9030 5488 9058
rect 5460 8362 5488 9030
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4214 5396 4558
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5460 2514 5488 8298
rect 5552 5302 5580 10610
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5552 4622 5580 5238
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5644 4554 5672 8434
rect 5736 7410 5764 8910
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5828 6322 5856 12406
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6012 10062 6040 10746
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5920 9450 5948 9998
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5920 8838 5948 9386
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 4826 5764 5646
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5644 3534 5672 4490
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5828 3942 5856 4082
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3670 5856 3878
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 3058 5672 3470
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5828 3194 5856 3334
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5814 2952 5870 2961
rect 5814 2887 5816 2896
rect 5868 2887 5870 2896
rect 5816 2858 5868 2864
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 5092 800 5120 2314
rect 5184 2038 5212 2382
rect 5172 2032 5224 2038
rect 5172 1974 5224 1980
rect 6012 800 6040 3402
rect 6104 1834 6132 18006
rect 6656 17054 6868 17082
rect 6656 16998 6684 17054
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6196 15570 6224 16662
rect 6644 16584 6696 16590
rect 6748 16572 6776 16934
rect 6696 16544 6776 16572
rect 6644 16526 6696 16532
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6380 12850 6408 13194
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6472 9722 6500 11222
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6564 9654 6592 16050
rect 6748 16046 6776 16544
rect 6840 16522 6868 17054
rect 6828 16516 6880 16522
rect 6828 16458 6880 16464
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14482 6868 14894
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6840 13870 6868 14418
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13326 6868 13806
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 10674 6868 13262
rect 6932 11150 6960 19246
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7024 16590 7052 16730
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7208 16114 7236 17614
rect 7300 17338 7328 20334
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14618 7144 14962
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7300 12434 7328 17138
rect 7392 14482 7420 25842
rect 7484 25294 7512 26182
rect 7472 25288 7524 25294
rect 7472 25230 7524 25236
rect 7668 25158 7696 26250
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7668 23186 7696 25094
rect 7760 23594 7788 35866
rect 10336 27606 10364 38286
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 14280 37936 14332 37942
rect 14280 37878 14332 37884
rect 11980 36780 12032 36786
rect 11980 36722 12032 36728
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 10416 30320 10468 30326
rect 10416 30262 10468 30268
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 8036 26042 8064 26386
rect 8024 26036 8076 26042
rect 8024 25978 8076 25984
rect 8036 25838 8064 25978
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 10232 25696 10284 25702
rect 10232 25638 10284 25644
rect 10244 24886 10272 25638
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10232 24880 10284 24886
rect 10232 24822 10284 24828
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9692 24206 9720 24686
rect 10336 24206 10364 25094
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 9692 23474 9720 24142
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9416 23446 9720 23474
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 7760 21146 7788 23054
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8220 22642 8248 22918
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7760 20602 7788 21082
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7024 12406 7328 12434
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6564 8974 6592 9590
rect 6656 9586 6684 9862
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6564 5166 6592 6190
rect 7024 5930 7052 12406
rect 7392 12374 7420 13126
rect 7484 12434 7512 19926
rect 8220 19854 8248 20334
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7760 15706 7788 16050
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 13734 7696 14418
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13394 7696 13670
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7484 12406 7604 12434
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7300 11898 7328 12174
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7300 11150 7328 11834
rect 7392 11694 7420 12310
rect 7576 12238 7604 12406
rect 7852 12238 7880 19722
rect 8220 19378 8248 19790
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7944 15638 7972 18702
rect 8220 17678 8248 19314
rect 8496 17814 8524 21558
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8588 20534 8616 21286
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8680 19922 8708 20198
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8496 17270 8524 17750
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8956 17338 8984 17546
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 8036 15910 8064 17206
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7944 13954 7972 15574
rect 8036 15570 8064 15846
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 7944 13926 8064 13954
rect 8036 12434 8064 13926
rect 8220 13462 8248 14282
rect 8312 14278 8340 14758
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 9048 13326 9076 22578
rect 9416 22574 9444 23446
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9416 20942 9444 22510
rect 9692 22234 9720 22578
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9140 19786 9168 20810
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9508 19174 9536 21490
rect 9600 20806 9628 21490
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 19446 9628 20742
rect 9692 20602 9720 21626
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9876 19514 9904 23530
rect 10428 22506 10456 30262
rect 10784 30116 10836 30122
rect 10784 30058 10836 30064
rect 10692 28484 10744 28490
rect 10692 28426 10744 28432
rect 10704 26042 10732 28426
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10704 24614 10732 25842
rect 10796 25362 10824 30058
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10888 25362 10916 25774
rect 10784 25356 10836 25362
rect 10784 25298 10836 25304
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10060 21146 10088 21966
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9600 18970 9628 19382
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9600 17202 9628 18906
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9784 18154 9812 18838
rect 9876 18698 9904 19450
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10152 18970 10180 19314
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 9968 18766 9996 18906
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16998 9628 17138
rect 10336 17066 10364 21966
rect 10428 21894 10456 22442
rect 10704 22438 10732 24550
rect 10796 24070 10824 25094
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10796 22710 10824 24006
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10428 20058 10456 20402
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10520 20058 10548 20198
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15366 9352 15846
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9140 13530 9168 13874
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8956 12714 8984 12922
rect 9048 12850 9076 13262
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 9232 12646 9260 14758
rect 9324 12782 9352 15302
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 13190 9444 13670
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 8036 12406 8248 12434
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7300 10606 7328 10678
rect 7392 10606 7420 10950
rect 7484 10606 7512 11494
rect 7576 11082 7604 12174
rect 7852 11694 7880 12174
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7116 10062 7144 10542
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9178 7144 9998
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 8498 7236 8842
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 7886 7236 8434
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7116 7342 7144 7754
rect 7208 7410 7236 7822
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6932 5914 7052 5930
rect 7116 5914 7144 7278
rect 6920 5908 7052 5914
rect 6972 5902 7052 5908
rect 6920 5850 6972 5856
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 5166 6868 5578
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6288 4554 6316 5102
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 3126 6408 4422
rect 6840 4010 6868 5102
rect 6932 4622 6960 5714
rect 7024 5710 7052 5902
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7208 5166 7236 7346
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7300 6390 7328 7142
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7300 5234 7328 6326
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 4146 6960 4558
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 6472 800 6500 3538
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 800 6960 2926
rect 7392 2774 7420 10542
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 8906 7512 10406
rect 7576 10130 7604 11018
rect 7852 10742 7880 11630
rect 8036 11150 8064 11698
rect 8128 11558 8156 12174
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7852 9586 7880 10678
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 8430 7512 8842
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7760 8498 7788 8570
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7760 7818 7788 8434
rect 7944 8430 7972 11086
rect 8220 10146 8248 12406
rect 8772 11830 8800 12582
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8312 11354 8340 11698
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8036 10118 8248 10146
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 5370 7604 6258
rect 7944 5574 7972 8366
rect 8036 6798 8064 10118
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 9586 8248 9998
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8312 9722 8340 9930
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 9178 8156 9318
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8220 9058 8248 9522
rect 8404 9518 8432 11222
rect 8772 11218 8800 11766
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8128 9030 8248 9058
rect 8128 8430 8156 9030
rect 8312 8838 8340 9114
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8128 7886 8156 8366
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8404 6866 8432 8298
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6390 8064 6734
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7576 4486 7604 5306
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7668 4078 7696 5102
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7944 3942 7972 5510
rect 8128 5302 8156 6054
rect 8312 5302 8340 6666
rect 8404 6458 8432 6802
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8312 5030 8340 5238
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4554 8432 4966
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3126 8432 3878
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8496 2990 8524 9386
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8242 8708 8842
rect 8864 8430 8892 9318
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8956 8242 8984 8298
rect 8680 8214 8984 8242
rect 8680 6254 8708 8214
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8588 4826 8616 6190
rect 8680 5778 8708 6190
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7116 2746 7420 2774
rect 7116 2446 7144 2746
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 7392 800 7420 2314
rect 7852 800 7880 2314
rect 8588 2310 8616 3470
rect 8680 3126 8708 5306
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8772 800 8800 2994
rect 8864 1698 8892 7686
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8956 6458 8984 7142
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9048 6458 9076 6666
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 3058 9168 3470
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9232 2922 9260 12582
rect 9324 5846 9352 12718
rect 9416 12646 9444 13126
rect 9600 12918 9628 13126
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9416 3466 9444 12582
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 11218 9536 11494
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9692 9926 9720 17002
rect 10520 16794 10548 19994
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 12434 9812 16526
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9784 12406 9904 12434
rect 9876 11082 9904 12406
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9968 11150 9996 11630
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10810 9812 10950
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 9994 9812 10406
rect 9876 10130 9904 11018
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9508 8634 9536 9590
rect 9784 9466 9812 9930
rect 9876 9654 9904 10066
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 9722 9996 9862
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9784 9438 9996 9466
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 7342 9628 9114
rect 9784 7546 9812 9318
rect 9968 9042 9996 9438
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 10060 8974 10088 12106
rect 10152 11370 10180 13262
rect 10244 11898 10272 13942
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10336 11626 10364 12106
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10152 11342 10364 11370
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9876 6662 9904 8910
rect 10046 8392 10102 8401
rect 9956 8356 10008 8362
rect 10046 8327 10102 8336
rect 9956 8298 10008 8304
rect 9968 8090 9996 8298
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 7886 10088 8327
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5642 9720 6122
rect 9876 5914 9904 6598
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10152 5710 10180 11222
rect 10336 10146 10364 11342
rect 10244 10118 10364 10146
rect 10244 8022 10272 10118
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10336 9586 10364 9930
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10336 8294 10364 8502
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 10244 4146 10272 7142
rect 10336 6458 10364 7346
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10428 3670 10456 12786
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11150 10548 11698
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10612 10470 10640 14010
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9110 10548 9522
rect 10612 9518 10640 10406
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 7206 10548 8366
rect 10612 8022 10640 8842
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10704 7410 10732 12038
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10506 5400 10562 5409
rect 10506 5335 10562 5344
rect 10520 5302 10548 5335
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10612 5234 10640 5510
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4622 10548 4966
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10704 3738 10732 6258
rect 10796 5166 10824 14282
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10888 7342 10916 12922
rect 10980 11218 11008 13126
rect 11072 12238 11100 21286
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11164 14414 11192 19722
rect 11256 15162 11284 27542
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11348 17542 11376 24074
rect 11716 23526 11744 35634
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11900 21622 11928 21898
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 11440 19922 11468 20470
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11256 14550 11284 15098
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11348 14414 11376 14826
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11164 14278 11192 14350
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11072 9654 11100 10134
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8634 11008 8842
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 8090 11008 8366
rect 11072 8090 11100 9386
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7954 11192 14214
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10888 6866 10916 7278
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 6186 10916 6666
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10888 5370 10916 5714
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9772 3188 9824 3194
rect 9956 3188 10008 3194
rect 9824 3148 9956 3176
rect 9772 3130 9824 3136
rect 9956 3130 10008 3136
rect 10796 3126 10824 4558
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 2446 9812 2790
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8852 1692 8904 1698
rect 8852 1634 8904 1640
rect 9232 800 9260 2246
rect 9692 870 9812 898
rect 9692 800 9720 870
rect 1122 776 1178 785
rect 1122 711 1178 720
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 9784 762 9812 870
rect 10060 762 10088 3062
rect 10980 3058 11008 7822
rect 11256 7818 11284 8434
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 7478 11192 7686
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11072 6934 11100 7278
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11072 6458 11100 6666
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11072 5710 11100 6394
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11348 5846 11376 6258
rect 11440 6186 11468 18770
rect 11532 16454 11560 21490
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11624 19854 11652 20402
rect 11716 20262 11744 21286
rect 11992 21146 12020 36722
rect 12440 32428 12492 32434
rect 12440 32370 12492 32376
rect 12452 29646 12480 32370
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 13544 29232 13596 29238
rect 13544 29174 13596 29180
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12820 22778 12848 22986
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12912 22574 12940 23054
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 12912 21570 12940 22510
rect 12912 21554 13032 21570
rect 12912 21548 13044 21554
rect 12912 21542 12992 21548
rect 12992 21490 13044 21496
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 11992 20602 12020 21082
rect 13004 20942 13032 21490
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12360 20602 12388 20810
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12452 20482 12480 20742
rect 12268 20466 12480 20482
rect 13004 20466 13032 20878
rect 11796 20460 11848 20466
rect 12256 20460 12480 20466
rect 11848 20420 12112 20448
rect 11796 20402 11848 20408
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11716 18970 11744 20198
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11808 18766 11836 19994
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11900 18766 11928 19858
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11716 18426 11744 18634
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11716 17338 11744 17546
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11532 15366 11560 16118
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11624 13870 11652 17070
rect 11808 16590 11836 18702
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 17270 12020 17478
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 15706 11744 16390
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11716 12850 11744 15030
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14618 11836 14962
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11900 13954 11928 15642
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11808 13926 11928 13954
rect 11992 13938 12020 14554
rect 11980 13932 12032 13938
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12434 11744 12786
rect 11624 12406 11744 12434
rect 11624 12306 11652 12406
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11624 11150 11652 12242
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 10130 11652 11086
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11808 10062 11836 13926
rect 11980 13874 12032 13880
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 13530 11928 13806
rect 12084 13734 12112 20420
rect 12308 20454 12480 20460
rect 12992 20460 13044 20466
rect 12256 20402 12308 20408
rect 12992 20402 13044 20408
rect 12348 20392 12400 20398
rect 12400 20340 12480 20346
rect 12348 20334 12480 20340
rect 12360 20318 12480 20334
rect 12452 18970 12480 20318
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 20058 12940 20198
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12820 19514 12848 19994
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12164 18624 12216 18630
rect 12452 18578 12480 18906
rect 13096 18873 13124 22578
rect 13280 22098 13308 22578
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13188 20942 13216 22034
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13280 20806 13308 22034
rect 13268 20800 13320 20806
rect 13268 20742 13320 20748
rect 13280 19922 13308 20742
rect 13464 20602 13492 23462
rect 13556 23322 13584 29174
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13648 24818 13676 26250
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13556 22778 13584 23258
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 14108 21962 14136 26862
rect 14292 22094 14320 37878
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 27172 35894 27200 39374
rect 28264 39364 28316 39370
rect 28264 39306 28316 39312
rect 27172 35866 27292 35894
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 22836 32496 22888 32502
rect 22836 32438 22888 32444
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 14648 26988 14700 26994
rect 14648 26930 14700 26936
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 14660 26314 14688 26930
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14752 26518 14780 26726
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14740 26512 14792 26518
rect 14740 26454 14792 26460
rect 14740 26376 14792 26382
rect 14844 26364 14872 26522
rect 14792 26336 14872 26364
rect 14740 26318 14792 26324
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14752 25906 14780 26318
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14752 24614 14780 25842
rect 14936 25838 14964 26862
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 15028 25702 15056 26318
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15120 26042 15148 26182
rect 15108 26036 15160 26042
rect 15108 25978 15160 25984
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15028 24886 15056 25230
rect 15396 25226 15424 26726
rect 15948 26586 15976 26930
rect 15936 26580 15988 26586
rect 15936 26522 15988 26528
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 15672 26194 15700 26250
rect 15580 26166 15700 26194
rect 15844 26240 15896 26246
rect 15844 26182 15896 26188
rect 15384 25220 15436 25226
rect 15384 25162 15436 25168
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 15028 24614 15056 24822
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 14752 24274 14780 24550
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14200 22066 14320 22094
rect 14096 21956 14148 21962
rect 14096 21898 14148 21904
rect 14108 21418 14136 21898
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13464 19854 13492 20538
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13740 20058 13768 20402
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13648 19922 13676 19994
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13082 18864 13138 18873
rect 13082 18799 13138 18808
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12216 18572 12480 18578
rect 12164 18566 12480 18572
rect 12176 18550 12480 18566
rect 12452 15434 12480 18550
rect 12912 16697 12940 18634
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17134 13032 17614
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12898 16688 12954 16697
rect 12898 16623 12954 16632
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 14278 12296 14758
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12176 13938 12204 14214
rect 12360 14006 12388 15030
rect 12820 14414 12848 15370
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12912 13870 12940 16623
rect 13004 16182 13032 17070
rect 12992 16176 13044 16182
rect 13188 16130 13216 19790
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13372 18970 13400 19722
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 14200 16250 14228 22066
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14292 21622 14320 21830
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17270 14320 17478
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 12992 16118 13044 16124
rect 13004 16046 13032 16118
rect 13096 16102 13216 16130
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 12176 12918 12204 13738
rect 12912 13394 12940 13806
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 12986 12388 13262
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11992 12442 12020 12786
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11898 12112 12174
rect 12360 12102 12388 12922
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12912 11354 12940 13194
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12268 10810 12296 11018
rect 12912 10810 12940 11290
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 6798 11560 8910
rect 11716 8430 11744 9318
rect 12360 9178 12388 9930
rect 12164 9172 12216 9178
rect 12348 9172 12400 9178
rect 12216 9132 12296 9160
rect 12164 9114 12216 9120
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12084 8634 12112 8842
rect 12268 8838 12296 9132
rect 12348 9114 12400 9120
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12176 8634 12204 8774
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12544 8498 12572 8774
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11716 8294 11744 8366
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11624 6730 11652 7890
rect 11716 7478 11744 8230
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11716 6662 11744 7414
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11808 6458 11836 6666
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11992 6322 12020 7142
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11060 5704 11112 5710
rect 11152 5704 11204 5710
rect 11060 5646 11112 5652
rect 11150 5672 11152 5681
rect 11204 5672 11206 5681
rect 11150 5607 11206 5616
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10152 800 10180 2314
rect 10612 800 10640 2314
rect 11164 1970 11192 4150
rect 11256 2990 11284 5782
rect 11348 5642 11376 5782
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11440 4826 11468 5646
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11334 4720 11390 4729
rect 11334 4655 11390 4664
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11348 2038 11376 4655
rect 11532 3602 11560 5850
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11992 5574 12020 5782
rect 12084 5642 12112 7278
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6322 12204 6598
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12360 5914 12388 8026
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12360 5370 12388 5578
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11532 800 11560 3402
rect 11716 1902 11744 4218
rect 11900 4146 11928 5306
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11900 3602 11928 4082
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12084 3738 12112 4014
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12176 3670 12204 4082
rect 12452 4026 12480 6938
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12544 4146 12572 6122
rect 12636 6118 12664 8774
rect 12728 8498 12756 10610
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9042 12940 9318
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12532 4140 12584 4146
rect 12584 4100 12664 4128
rect 12532 4082 12584 4088
rect 12452 3998 12572 4026
rect 12544 3942 12572 3998
rect 12636 3942 12664 4100
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11808 3466 11836 3538
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 12820 2553 12848 3470
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12806 2544 12862 2553
rect 12806 2479 12862 2488
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 11992 800 12020 2246
rect 12452 800 12480 2314
rect 12912 800 12940 2926
rect 13096 2774 13124 16102
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14482 13492 14758
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 13938 13676 14282
rect 14108 14074 14136 15438
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13188 6390 13216 13330
rect 13268 12436 13320 12442
rect 14384 12434 14412 22646
rect 14660 17678 14688 22986
rect 15028 22642 15056 24550
rect 15580 24206 15608 26166
rect 15856 25906 15884 26182
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15856 25498 15884 25842
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 15844 25492 15896 25498
rect 15844 25434 15896 25440
rect 15948 24410 15976 25774
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16132 24410 16160 24754
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15580 23594 15608 24142
rect 15568 23588 15620 23594
rect 15568 23530 15620 23536
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15948 21622 15976 24346
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16592 23322 16620 24074
rect 17040 23792 17092 23798
rect 16960 23740 17040 23746
rect 16960 23734 17092 23740
rect 16960 23718 17080 23734
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16868 23118 16896 23462
rect 16960 23254 16988 23718
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16948 23248 17000 23254
rect 16948 23190 17000 23196
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16776 22166 16804 23054
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16868 22506 16896 22918
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 14832 20528 14884 20534
rect 14832 20470 14884 20476
rect 14844 19854 14872 20470
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19378 14872 19790
rect 15120 19786 15148 20810
rect 15304 20262 15332 20810
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14752 17678 14780 18226
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14476 16794 14504 17614
rect 14660 17066 14688 17614
rect 14752 17202 14780 17614
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 13530 14504 13874
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 13268 12378 13320 12384
rect 14292 12406 14412 12434
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13176 3732 13228 3738
rect 13280 3720 13308 12378
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14200 11830 14228 12174
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13832 10606 13860 11154
rect 14200 11150 14228 11630
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 14292 9110 14320 12406
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14384 10742 14412 12174
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14476 10674 14504 11086
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13372 7546 13400 7822
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13464 7002 13492 7822
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13360 5228 13412 5234
rect 13464 5216 13492 6734
rect 13556 6322 13584 7958
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13412 5188 13492 5216
rect 13360 5170 13412 5176
rect 13228 3692 13308 3720
rect 13176 3674 13228 3680
rect 13188 3534 13216 3674
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13372 3534 13400 3606
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13464 3058 13492 5188
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3534 13584 3878
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13740 3398 13768 8434
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 7954 14044 8230
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14016 6390 14044 7890
rect 14200 7886 14228 8434
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14292 8022 14320 8366
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7478 14136 7686
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14108 6390 14136 7414
rect 14568 7206 14596 16526
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14660 15502 14688 16186
rect 14752 15502 14780 17138
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14844 15706 14872 16050
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 15028 14958 15056 18158
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14844 13326 14872 14010
rect 14936 13326 14964 14350
rect 15120 14278 15148 19722
rect 15304 17746 15332 20198
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16132 19786 16160 19994
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16132 19514 16160 19722
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16500 19446 16528 19654
rect 16776 19514 16804 22102
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 16408 17202 16436 18702
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15212 16182 15240 16594
rect 15292 16584 15344 16590
rect 15290 16552 15292 16561
rect 15344 16552 15346 16561
rect 15290 16487 15346 16496
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14936 10606 14964 13262
rect 15120 11150 15148 14214
rect 15396 13462 15424 16594
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10062 14964 10542
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 15028 9674 15056 11018
rect 15304 10810 15332 12582
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15028 9646 15148 9674
rect 15120 9450 15148 9646
rect 15198 9616 15254 9625
rect 15198 9551 15200 9560
rect 15252 9551 15254 9560
rect 15292 9580 15344 9586
rect 15200 9522 15252 9528
rect 15292 9522 15344 9528
rect 15304 9489 15332 9522
rect 15290 9480 15346 9489
rect 15108 9444 15160 9450
rect 15290 9415 15346 9424
rect 15108 9386 15160 9392
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14936 7954 14964 8434
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15028 7410 15056 8026
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 15120 6798 15148 9386
rect 15304 7886 15332 9415
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5030 14044 6054
rect 14108 5370 14136 6326
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5710 14504 6054
rect 14752 5710 14780 6326
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14464 5704 14516 5710
rect 14740 5704 14792 5710
rect 14464 5646 14516 5652
rect 14646 5672 14702 5681
rect 14740 5646 14792 5652
rect 14646 5607 14648 5616
rect 14700 5607 14702 5616
rect 14648 5578 14700 5584
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14292 5234 14320 5510
rect 14660 5370 14688 5578
rect 14844 5409 14872 6122
rect 14830 5400 14886 5409
rect 14648 5364 14700 5370
rect 14830 5335 14886 5344
rect 14648 5306 14700 5312
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4146 14780 4966
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4146 14872 4422
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14002 3496 14058 3505
rect 14002 3431 14058 3440
rect 14280 3460 14332 3466
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13648 3126 13676 3334
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 14016 2938 14044 3431
rect 14280 3402 14332 3408
rect 13924 2922 14044 2938
rect 13912 2916 14044 2922
rect 13964 2910 14044 2916
rect 13912 2858 13964 2864
rect 13004 2746 13124 2774
rect 13004 2038 13032 2746
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 13280 1766 13308 2382
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 13268 1760 13320 1766
rect 13268 1702 13320 1708
rect 13372 800 13400 2314
rect 14292 800 14320 3402
rect 14660 3126 14688 3878
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14936 2446 14964 4082
rect 15198 3088 15254 3097
rect 15198 3023 15254 3032
rect 15212 2854 15240 3023
rect 15304 2854 15332 4490
rect 15396 4078 15424 12038
rect 15488 11898 15516 12310
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15580 11898 15608 12106
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15474 9616 15530 9625
rect 15474 9551 15476 9560
rect 15528 9551 15530 9560
rect 15476 9522 15528 9528
rect 15764 7818 15792 11698
rect 15856 10742 15884 17138
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 16250 16344 16390
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16408 16130 16436 17138
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16592 16590 16620 16934
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16316 16102 16436 16130
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16224 13938 16252 14486
rect 16316 14346 16344 16102
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16040 11762 16068 12582
rect 16316 12434 16344 14282
rect 16500 14074 16528 14282
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16592 14006 16620 14282
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16684 13784 16712 18158
rect 16592 13756 16712 13784
rect 16592 13462 16620 13756
rect 16776 13682 16804 19450
rect 16868 18222 16896 22442
rect 16960 22438 16988 23190
rect 17052 22642 17080 23190
rect 17144 23118 17172 23598
rect 17788 23526 17816 25774
rect 19076 24818 19104 27270
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27130 20024 27270
rect 20640 27130 20668 27406
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19260 25974 19288 26250
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 19352 25770 19380 27066
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 19536 26858 19564 26930
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19524 26852 19576 26858
rect 19524 26794 19576 26800
rect 19812 26790 19840 26862
rect 19800 26784 19852 26790
rect 19800 26726 19852 26732
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19628 25294 19656 25638
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19616 25288 19668 25294
rect 19616 25230 19668 25236
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 17880 24206 17908 24550
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17880 23730 17908 24142
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17788 23118 17816 23462
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17788 22642 17816 23054
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 17610 16896 18022
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16960 16114 16988 22374
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 20874 17724 21966
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17696 20330 17724 20810
rect 17788 20534 17816 21286
rect 17972 21146 18000 21558
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 18064 19922 18092 21830
rect 18432 20942 18460 22714
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18524 21146 18552 21354
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18524 20398 18552 21082
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17052 17338 17080 18226
rect 17144 17882 17172 18226
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17224 18148 17276 18154
rect 17276 18108 17356 18136
rect 17224 18090 17276 18096
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17038 16688 17094 16697
rect 17038 16623 17040 16632
rect 17092 16623 17094 16632
rect 17040 16594 17092 16600
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16684 13654 16804 13682
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16684 13326 16712 13654
rect 16960 13530 16988 16050
rect 17052 15638 17080 16458
rect 17144 16454 17172 17070
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17236 15042 17264 17546
rect 17328 17338 17356 18108
rect 17972 17678 18000 18158
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17420 17202 17448 17478
rect 17972 17202 18000 17614
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17144 15014 17264 15042
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16672 13320 16724 13326
rect 16224 12406 16344 12434
rect 16592 13280 16672 13308
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16224 11150 16252 12406
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16316 11354 16344 12242
rect 16500 12102 16528 12242
rect 16592 12238 16620 13280
rect 16672 13262 16724 13268
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11830 16528 12038
rect 16592 11898 16620 12174
rect 16684 12102 16712 12922
rect 16776 12238 16804 13466
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16868 12986 16896 13330
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 12442 16896 12786
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16684 11558 16712 12038
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16040 8906 16068 9318
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 16040 5234 16068 8842
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15948 4826 15976 5034
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16132 4486 16160 8910
rect 16224 8430 16252 11086
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16500 10130 16528 10678
rect 16592 10198 16620 11154
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16500 9353 16528 9386
rect 16486 9344 16542 9353
rect 16486 9279 16542 9288
rect 16592 8974 16620 9658
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16684 8634 16712 9930
rect 16776 9926 16804 11698
rect 17144 11150 17172 15014
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17236 11898 17264 12786
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 8906 16804 9862
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16212 8424 16264 8430
rect 16868 8401 16896 10610
rect 17144 10282 17172 11086
rect 17144 10254 17264 10282
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16960 9110 16988 9590
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 17052 8616 17080 9998
rect 17144 9382 17172 10066
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 8974 17172 9318
rect 17236 9110 17264 10254
rect 17328 10062 17356 16594
rect 17406 16552 17462 16561
rect 17406 16487 17462 16496
rect 17420 16454 17448 16487
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17512 15706 17540 17138
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17512 15570 17540 15642
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17512 14550 17540 14894
rect 17500 14544 17552 14550
rect 17420 14492 17500 14498
rect 17420 14486 17552 14492
rect 17420 14470 17540 14486
rect 17420 14074 17448 14470
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17512 13326 17540 14350
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17512 11898 17540 13262
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17420 9489 17448 9522
rect 17406 9480 17462 9489
rect 17406 9415 17462 9424
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17132 8628 17184 8634
rect 17052 8588 17132 8616
rect 16212 8366 16264 8372
rect 16854 8392 16910 8401
rect 16488 8356 16540 8362
rect 16854 8327 16910 8336
rect 16488 8298 16540 8304
rect 16500 8090 16528 8298
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16684 7002 16712 7346
rect 17052 7342 17080 8588
rect 17132 8570 17184 8576
rect 17512 8498 17540 9046
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17224 7268 17276 7274
rect 17224 7210 17276 7216
rect 17236 7002 17264 7210
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 16684 6662 16712 6938
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 17236 6254 17264 6666
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4622 16252 4966
rect 16212 4616 16264 4622
rect 16264 4576 16344 4604
rect 16212 4558 16264 4564
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16132 3466 16160 3606
rect 16316 3534 16344 4576
rect 16500 4554 16528 5238
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3534 16620 3878
rect 16762 3632 16818 3641
rect 16762 3567 16818 3576
rect 16776 3534 16804 3567
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16776 3398 16804 3470
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15304 2582 15332 2790
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 800 14780 2246
rect 15212 800 15240 2314
rect 15672 800 15700 2926
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15856 1970 15884 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15844 1964 15896 1970
rect 15844 1906 15896 1912
rect 16132 800 16160 2314
rect 17052 800 17080 4150
rect 17328 3738 17356 8434
rect 17420 8362 17448 8434
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17420 6798 17448 7754
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17420 6458 17448 6734
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17512 6390 17540 6734
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17420 3534 17448 4490
rect 17604 4282 17632 16118
rect 17696 9722 17724 16526
rect 17880 13734 17908 17002
rect 18248 16250 18276 17138
rect 18524 16250 18552 17274
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18616 16114 18644 20742
rect 18800 20466 18828 24550
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 18892 22778 18920 23462
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18892 16182 18920 22578
rect 19352 22574 19380 25094
rect 19444 24342 19472 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19432 24336 19484 24342
rect 19432 24278 19484 24284
rect 19628 24070 19656 24754
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19720 24070 19748 24210
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20088 23798 20116 26522
rect 20364 26382 20392 26930
rect 20444 26852 20496 26858
rect 20444 26794 20496 26800
rect 20456 26382 20484 26794
rect 20640 26790 20668 27066
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 20548 26602 20576 26726
rect 20548 26574 20760 26602
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20456 26042 20484 26318
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20456 24954 20484 25978
rect 20444 24948 20496 24954
rect 20444 24890 20496 24896
rect 20548 24698 20576 26574
rect 20628 26512 20680 26518
rect 20628 26454 20680 26460
rect 20640 26382 20668 26454
rect 20732 26382 20760 26574
rect 22020 26382 22048 26726
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20720 26376 20772 26382
rect 20720 26318 20772 26324
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 20640 24818 20668 26318
rect 21548 26240 21600 26246
rect 21548 26182 21600 26188
rect 21560 25294 21588 26182
rect 22296 25498 22324 26318
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20548 24670 20668 24698
rect 20916 24682 20944 25230
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19352 22234 19380 22510
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 19720 22166 19748 22374
rect 19708 22160 19760 22166
rect 19708 22102 19760 22108
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 19720 22030 19748 22102
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19260 19854 19288 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19352 20058 19380 20402
rect 19996 20346 20024 21422
rect 20088 20618 20116 22102
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20180 21622 20208 21966
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20088 20590 20208 20618
rect 20180 20534 20208 20590
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 19996 20318 20116 20346
rect 20180 20330 20208 20470
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19444 19854 19472 20198
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 17678 19380 18566
rect 19444 18408 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20088 18766 20116 20318
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20272 19854 20300 22986
rect 20364 22506 20392 24550
rect 20536 24132 20588 24138
rect 20536 24074 20588 24080
rect 20548 23798 20576 24074
rect 20536 23792 20588 23798
rect 20536 23734 20588 23740
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20456 23050 20484 23598
rect 20444 23044 20496 23050
rect 20444 22986 20496 22992
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 20364 21554 20392 22442
rect 20640 22094 20668 24670
rect 20904 24676 20956 24682
rect 20904 24618 20956 24624
rect 20916 24274 20944 24618
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21008 23730 21036 24006
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 20456 22066 20668 22094
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20456 21486 20484 22066
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20732 20398 20760 21830
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20824 19854 20852 23054
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 20942 21036 21286
rect 21376 20942 21404 22986
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 21622 22140 22918
rect 22204 22710 22232 23054
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22296 22030 22324 22578
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22100 21616 22152 21622
rect 22100 21558 22152 21564
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21376 19854 21404 20878
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18634
rect 19984 18420 20036 18426
rect 19444 18380 19564 18408
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 17882 19472 18226
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19536 17814 19564 18380
rect 19984 18362 20036 18368
rect 19524 17808 19576 17814
rect 19444 17756 19524 17762
rect 19444 17750 19576 17756
rect 19444 17734 19564 17750
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 16182 19012 16934
rect 19444 16658 19472 17734
rect 19996 17610 20024 18362
rect 20088 17678 20116 18702
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 20088 16454 20116 17614
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18064 15910 18092 15982
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 18616 15026 18644 16050
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18616 14550 18644 14962
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 18064 12434 18092 14350
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 17972 12406 18092 12434
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17788 11898 17816 12242
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 11354 17908 11698
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17972 11014 18000 12406
rect 18156 11898 18184 13942
rect 18616 13938 18644 14486
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 12986 18552 13194
rect 18616 12986 18644 13874
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18800 12434 18828 15846
rect 19812 15570 19840 15982
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12918 18920 13126
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18800 12406 19012 12434
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 10130 17908 10542
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17696 8634 17724 8842
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17788 8022 17816 9930
rect 17880 9353 17908 10066
rect 17866 9344 17922 9353
rect 17866 9279 17922 9288
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17788 7818 17816 7958
rect 17880 7954 17908 9279
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7478 17816 7754
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17880 4214 17908 5034
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17972 4146 18000 4490
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 17880 3534 17908 3567
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17406 2544 17462 2553
rect 17406 2479 17462 2488
rect 17420 2446 17448 2479
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17512 800 17540 2926
rect 17972 2854 18000 4082
rect 18064 3738 18092 11018
rect 18156 8498 18184 11834
rect 18432 11150 18460 12038
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 11150 18644 11494
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18236 10804 18288 10810
rect 18432 10792 18460 11086
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18432 10764 18552 10792
rect 18236 10746 18288 10752
rect 18248 8498 18276 10746
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18340 9654 18368 10678
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18432 10198 18460 10610
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18340 7886 18368 9590
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18524 5710 18552 10764
rect 18892 10062 18920 10950
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18800 5914 18828 6190
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18892 5710 18920 6054
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18524 5234 18552 5646
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4554 18276 4966
rect 18524 4554 18552 5170
rect 18708 5166 18736 5578
rect 18984 5302 19012 12406
rect 19076 12102 19104 15438
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19444 15162 19472 15370
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19892 15088 19944 15094
rect 19996 15076 20024 15302
rect 19944 15048 20024 15076
rect 19892 15030 19944 15036
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19168 9110 19196 13466
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19352 10810 19380 11290
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19156 8968 19208 8974
rect 19260 8922 19288 9930
rect 19208 8916 19288 8922
rect 19156 8910 19288 8916
rect 19168 8894 19288 8910
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19168 7546 19196 7754
rect 19260 7698 19288 8894
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19352 7886 19380 8842
rect 19444 8634 19472 12718
rect 20180 12434 20208 18838
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 18086 20760 18566
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 16046 20300 17478
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16114 20760 16662
rect 20824 16522 20852 19790
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20916 19514 20944 19654
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20916 18766 20944 19450
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 21008 18766 21036 19382
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 21008 16182 21036 18702
rect 21468 18630 21496 18702
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 18358 21496 18566
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21364 16720 21416 16726
rect 21364 16662 21416 16668
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 20720 16108 20772 16114
rect 20772 16068 20852 16096
rect 20720 16050 20772 16056
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15162 20760 15846
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20180 12406 20300 12434
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20180 11830 20208 12106
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9586 20024 11494
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19996 8514 20024 9522
rect 19904 8498 20024 8514
rect 19892 8492 20024 8498
rect 19944 8486 20024 8492
rect 19892 8434 19944 8440
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19260 7670 19380 7698
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19352 7410 19380 7670
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6254 19288 6734
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19168 5370 19196 6190
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 18972 5296 19024 5302
rect 19352 5273 19380 7346
rect 19444 5778 19472 7890
rect 19996 7886 20024 8366
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19628 6798 19656 7346
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 18972 5238 19024 5244
rect 19338 5264 19394 5273
rect 19338 5199 19394 5208
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 19340 4616 19392 4622
rect 19260 4564 19340 4570
rect 19260 4558 19392 4564
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 19260 4542 19380 4558
rect 19260 4146 19288 4542
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 19444 3534 19472 5714
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19812 4622 19840 4694
rect 19996 4622 20024 7822
rect 20088 7410 20116 9862
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20088 4758 20116 7346
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 18984 3058 19012 3470
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 17880 898 17908 2314
rect 17880 870 18000 898
rect 17972 800 18000 870
rect 18432 800 18460 2926
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18708 950 18736 2314
rect 18696 944 18748 950
rect 18696 886 18748 892
rect 19352 800 19380 3402
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3126 20024 4422
rect 20180 3738 20208 8366
rect 20272 7478 20300 12406
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20364 11898 20392 12106
rect 20640 11898 20668 13806
rect 20824 13326 20852 16068
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 21008 13258 21036 16118
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21100 15706 21128 15982
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21192 15570 21220 16526
rect 21376 16454 21404 16662
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21284 15570 21312 16050
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21284 15026 21312 15370
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 13938 21312 14962
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 21100 13530 21128 13806
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21376 12238 21404 12582
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 21008 9926 21036 11562
rect 21376 11354 21404 11630
rect 21560 11626 21588 13874
rect 21652 12170 21680 21286
rect 22204 21146 22232 21898
rect 22848 21894 22876 32438
rect 23768 22778 23796 33458
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24412 26450 24440 26726
rect 24400 26444 24452 26450
rect 24400 26386 24452 26392
rect 24596 26382 24624 26726
rect 24860 26512 24912 26518
rect 24860 26454 24912 26460
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24872 25294 24900 26454
rect 24964 26314 24992 26930
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24596 24886 24624 25230
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24596 24274 24624 24822
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 24780 24410 24808 24754
rect 25608 24614 25636 29582
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25976 25498 26004 26250
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24584 24268 24636 24274
rect 24584 24210 24636 24216
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23400 22234 23428 22578
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23768 22030 23796 22714
rect 24596 22642 24624 24210
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22296 21026 22324 21830
rect 22204 20998 22324 21026
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21744 16697 21772 18702
rect 22204 18426 22232 20998
rect 22572 20942 22600 21830
rect 23492 21146 23520 21966
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22296 18902 22324 19722
rect 22388 18970 22416 20878
rect 22928 19236 22980 19242
rect 22928 19178 22980 19184
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22652 18896 22704 18902
rect 22704 18856 22784 18884
rect 22652 18838 22704 18844
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22020 17678 22048 18022
rect 22112 17882 22140 18226
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22204 17678 22232 18362
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 21730 16688 21786 16697
rect 21730 16623 21786 16632
rect 21744 16114 21772 16623
rect 21732 16108 21784 16114
rect 21732 16050 21784 16056
rect 21836 14074 21864 17614
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 15450 21956 17478
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22020 15570 22048 15846
rect 22112 15706 22140 16050
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22204 15502 22232 16458
rect 22100 15496 22152 15502
rect 21928 15422 22048 15450
rect 22100 15438 22152 15444
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21744 12986 21772 13262
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21652 11694 21680 11834
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 11150 21404 11290
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21284 10062 21312 10950
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 21008 9586 21036 9862
rect 21560 9674 21588 11562
rect 21088 9648 21140 9654
rect 21560 9646 21680 9674
rect 21088 9590 21140 9596
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20364 8498 20392 8978
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20732 8090 20760 9318
rect 21100 8498 21128 9590
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 20812 8288 20864 8294
rect 20864 8236 20944 8242
rect 20812 8230 20944 8236
rect 20824 8214 20944 8230
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20916 7818 20944 8214
rect 21192 8090 21220 8366
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 7546 20852 7686
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20260 7472 20312 7478
rect 20260 7414 20312 7420
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20456 5846 20484 6258
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19800 944 19852 950
rect 19800 886 19852 892
rect 19812 800 19840 886
rect 20272 800 20300 4014
rect 20364 3505 20392 4082
rect 20824 3670 20852 5714
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20812 3664 20864 3670
rect 20626 3632 20682 3641
rect 20812 3606 20864 3612
rect 20626 3567 20628 3576
rect 20680 3567 20682 3576
rect 20628 3538 20680 3544
rect 20536 3528 20588 3534
rect 20350 3496 20406 3505
rect 20536 3470 20588 3476
rect 20350 3431 20406 3440
rect 20548 2854 20576 3470
rect 20824 3058 20852 3606
rect 20916 3058 20944 4082
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21008 3058 21036 3334
rect 21100 3097 21128 3470
rect 21284 3398 21312 9318
rect 21468 9042 21496 9318
rect 21652 9042 21680 9646
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21560 3194 21588 8910
rect 21652 8294 21680 8978
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 8090 21680 8230
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21640 3460 21692 3466
rect 21640 3402 21692 3408
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21086 3088 21142 3097
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 20996 3052 21048 3058
rect 21086 3023 21142 3032
rect 20996 2994 21048 3000
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 898 20668 2314
rect 20640 870 20760 898
rect 20732 800 20760 870
rect 21652 800 21680 3402
rect 21836 2582 21864 4422
rect 21824 2576 21876 2582
rect 21824 2518 21876 2524
rect 21928 1358 21956 14282
rect 22020 13938 22048 15422
rect 22112 15094 22140 15438
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22112 13326 22140 15030
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22112 12918 22140 13262
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22204 12850 22232 15438
rect 22756 15434 22784 18856
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22848 17882 22876 18702
rect 22940 18426 22968 19178
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 11150 22140 12582
rect 22296 11898 22324 12786
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22190 11792 22246 11801
rect 22190 11727 22192 11736
rect 22244 11727 22246 11736
rect 22192 11698 22244 11704
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22112 9994 22140 11086
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22296 10266 22324 11018
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22296 9654 22324 10202
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22020 6866 22048 8366
rect 22112 8362 22140 8842
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22112 7750 22140 8298
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 6322 22140 6598
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22020 5778 22048 6258
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22112 5710 22140 6258
rect 22204 6186 22232 8230
rect 22296 6361 22324 9454
rect 22480 8786 22508 13670
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22572 12782 22600 13330
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22572 12442 22600 12718
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22664 10826 22692 12854
rect 22756 12782 22784 15370
rect 23216 15026 23244 20946
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23584 19922 23612 20810
rect 23676 20058 23704 20878
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23492 19446 23520 19654
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23308 16522 23336 18702
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23308 14958 23336 16458
rect 23400 15706 23428 17682
rect 23584 17542 23612 19858
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23676 18086 23704 18770
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23492 16658 23520 16934
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23584 16454 23612 17138
rect 23676 17066 23704 18022
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23676 16590 23704 17002
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23768 16017 23796 20878
rect 24964 20058 24992 24142
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25056 22234 25084 22578
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 25240 22030 25268 24142
rect 25608 24138 25636 24550
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 26068 22778 26096 31282
rect 26148 24132 26200 24138
rect 26148 24074 26200 24080
rect 26160 23866 26188 24074
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 26332 23724 26384 23730
rect 26332 23666 26384 23672
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 25332 20806 25360 21966
rect 26068 21962 26096 22714
rect 26344 22098 26372 23666
rect 26516 23520 26568 23526
rect 26516 23462 26568 23468
rect 26528 23322 26556 23462
rect 26516 23316 26568 23322
rect 26516 23258 26568 23264
rect 26332 22092 26384 22098
rect 26332 22034 26384 22040
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 26344 21622 26372 22034
rect 26332 21616 26384 21622
rect 26332 21558 26384 21564
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25792 21078 25820 21286
rect 25780 21072 25832 21078
rect 25780 21014 25832 21020
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24400 19780 24452 19786
rect 24400 19722 24452 19728
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24320 19514 24348 19654
rect 24412 19514 24440 19722
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 24400 19508 24452 19514
rect 24400 19450 24452 19456
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18358 23980 19110
rect 24780 18834 24808 19790
rect 24872 19242 24900 19790
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24872 18766 24900 19178
rect 24860 18760 24912 18766
rect 24912 18720 24992 18748
rect 24860 18702 24912 18708
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 23952 17270 23980 18294
rect 24780 18222 24808 18634
rect 24964 18290 24992 18720
rect 25056 18426 25084 19790
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24780 18086 24808 18158
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24872 17898 24900 18226
rect 24596 17870 24900 17898
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23754 16008 23810 16017
rect 23754 15943 23810 15952
rect 23860 15892 23888 16458
rect 23676 15864 23888 15892
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 22928 14884 22980 14890
rect 22928 14826 22980 14832
rect 22940 13462 22968 14826
rect 23032 14074 23060 14894
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23308 13870 23336 14894
rect 23676 13938 23704 15864
rect 23952 15026 23980 17206
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 23676 13326 23704 13874
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23768 13258 23796 13942
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23386 11792 23442 11801
rect 23386 11727 23442 11736
rect 22572 10810 22692 10826
rect 22560 10804 22692 10810
rect 22612 10798 22692 10804
rect 22560 10746 22612 10752
rect 22572 9586 22600 10746
rect 23400 10033 23428 11727
rect 23492 11665 23520 12718
rect 23860 12238 23888 14758
rect 23940 13932 23992 13938
rect 24044 13920 24072 16730
rect 24136 15094 24164 17138
rect 24596 17134 24624 17870
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24676 17128 24728 17134
rect 24860 17128 24912 17134
rect 24676 17070 24728 17076
rect 24780 17076 24860 17082
rect 24780 17070 24912 17076
rect 24228 16590 24256 17070
rect 24688 16590 24716 17070
rect 24780 17054 24900 17070
rect 24780 16794 24808 17054
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24780 16522 24808 16730
rect 24964 16658 24992 16730
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 25056 16182 25084 16526
rect 25148 16250 25176 19926
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25608 18834 25636 19246
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25608 18222 25636 18770
rect 25884 18630 25912 21422
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25976 21010 26004 21286
rect 25964 21004 26016 21010
rect 25964 20946 26016 20952
rect 26160 20942 26188 21422
rect 26252 20942 26280 21422
rect 27068 21412 27120 21418
rect 27068 21354 27120 21360
rect 27080 20942 27108 21354
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 26068 19938 26096 20878
rect 26160 20398 26188 20878
rect 26252 20398 26280 20878
rect 26792 20800 26844 20806
rect 26792 20742 26844 20748
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26148 20392 26200 20398
rect 26148 20334 26200 20340
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26332 20324 26384 20330
rect 26332 20266 26384 20272
rect 26068 19910 26188 19938
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26068 19514 26096 19790
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25964 19440 26016 19446
rect 25964 19382 26016 19388
rect 25976 19242 26004 19382
rect 25964 19236 26016 19242
rect 25964 19178 26016 19184
rect 26160 18970 26188 19910
rect 26344 19854 26372 20266
rect 26712 19922 26740 20538
rect 26804 20466 26832 20742
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26884 20392 26936 20398
rect 26884 20334 26936 20340
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25240 16590 25268 17478
rect 25318 16688 25374 16697
rect 25318 16623 25320 16632
rect 25372 16623 25374 16632
rect 25320 16594 25372 16600
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25608 16182 25636 18158
rect 25044 16176 25096 16182
rect 24674 16144 24730 16153
rect 24492 16108 24544 16114
rect 25044 16118 25096 16124
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25700 16114 25728 18226
rect 25884 18222 25912 18362
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 25884 16697 25912 18158
rect 26252 17610 26280 19790
rect 26344 18698 26372 19790
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26528 19174 26556 19246
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26424 18896 26476 18902
rect 26422 18864 26424 18873
rect 26476 18864 26478 18873
rect 26422 18799 26478 18808
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 26528 18426 26556 19110
rect 26896 18766 26924 20334
rect 26988 18902 27016 20878
rect 27080 20466 27108 20878
rect 27172 20602 27200 21490
rect 27264 21078 27292 35866
rect 28276 26450 28304 39306
rect 33324 39296 33376 39302
rect 33324 39238 33376 39244
rect 33336 35894 33364 39238
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 33244 35866 33364 35894
rect 31944 28416 31996 28422
rect 31944 28358 31996 28364
rect 28264 26444 28316 26450
rect 28264 26386 28316 26392
rect 28724 26444 28776 26450
rect 28724 26386 28776 26392
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 27724 24206 27752 24754
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 28264 23588 28316 23594
rect 28264 23530 28316 23536
rect 28276 23186 28304 23530
rect 28736 23254 28764 26386
rect 30288 25968 30340 25974
rect 30288 25910 30340 25916
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 29000 25832 29052 25838
rect 29000 25774 29052 25780
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 28920 24818 28948 25298
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28816 24744 28868 24750
rect 28816 24686 28868 24692
rect 28828 24614 28856 24686
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 29012 24410 29040 25774
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 29932 24818 29960 25638
rect 30012 25288 30064 25294
rect 30012 25230 30064 25236
rect 30024 24954 30052 25230
rect 30012 24948 30064 24954
rect 30012 24890 30064 24896
rect 30116 24886 30144 25842
rect 30104 24880 30156 24886
rect 30104 24822 30156 24828
rect 29920 24812 29972 24818
rect 29920 24754 29972 24760
rect 29736 24676 29788 24682
rect 29736 24618 29788 24624
rect 29368 24608 29420 24614
rect 29368 24550 29420 24556
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 29012 23526 29040 24346
rect 29380 23798 29408 24550
rect 29460 24336 29512 24342
rect 29460 24278 29512 24284
rect 29368 23792 29420 23798
rect 29368 23734 29420 23740
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 28724 23248 28776 23254
rect 28724 23190 28776 23196
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28736 23118 28764 23190
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28724 23112 28776 23118
rect 28724 23054 28776 23060
rect 28368 22982 28396 23054
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28460 22778 28488 23054
rect 29184 23044 29236 23050
rect 29184 22986 29236 22992
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 29104 22522 29132 22918
rect 29196 22710 29224 22986
rect 29184 22704 29236 22710
rect 29184 22646 29236 22652
rect 29104 22494 29224 22522
rect 29196 22234 29224 22494
rect 27528 22228 27580 22234
rect 27528 22170 27580 22176
rect 29184 22228 29236 22234
rect 29184 22170 29236 22176
rect 27540 22098 27568 22170
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 27252 21072 27304 21078
rect 27252 21014 27304 21020
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27356 20398 27384 21422
rect 27540 21146 27568 21422
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27632 20942 27660 21422
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28552 21010 28580 21286
rect 28644 21010 28672 21422
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28632 21004 28684 21010
rect 28632 20946 28684 20952
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27632 20398 27660 20878
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 27160 20392 27212 20398
rect 27160 20334 27212 20340
rect 27344 20392 27396 20398
rect 27344 20334 27396 20340
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27528 20392 27580 20398
rect 27528 20334 27580 20340
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27172 19378 27200 20334
rect 27448 19446 27476 20334
rect 27540 19990 27568 20334
rect 27528 19984 27580 19990
rect 27528 19926 27580 19932
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27448 19310 27476 19382
rect 27632 19310 27660 20334
rect 28736 19854 28764 20810
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 28816 20460 28868 20466
rect 28816 20402 28868 20408
rect 28828 20058 28856 20402
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27620 19304 27672 19310
rect 27620 19246 27672 19252
rect 27160 19236 27212 19242
rect 27160 19178 27212 19184
rect 26976 18896 27028 18902
rect 26976 18838 27028 18844
rect 27172 18834 27200 19178
rect 27356 18902 27384 19246
rect 27540 19174 27568 19246
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27344 18896 27396 18902
rect 27344 18838 27396 18844
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 28736 18766 28764 19790
rect 28920 19718 28948 20538
rect 29196 19718 29224 22170
rect 29368 19916 29420 19922
rect 29368 19858 29420 19864
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 28920 19378 28948 19654
rect 29196 19378 29224 19654
rect 29380 19378 29408 19858
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 26700 18760 26752 18766
rect 26700 18702 26752 18708
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 26712 18426 26740 18702
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 26896 18154 26924 18702
rect 26884 18148 26936 18154
rect 26884 18090 26936 18096
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27448 16794 27476 17138
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 25870 16688 25926 16697
rect 27540 16658 27568 17614
rect 25870 16623 25926 16632
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27540 16454 27568 16594
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 24492 16050 24544 16056
rect 24596 16088 24674 16096
rect 24596 16068 24676 16088
rect 24124 15088 24176 15094
rect 24124 15030 24176 15036
rect 23992 13892 24072 13920
rect 23940 13874 23992 13880
rect 23952 12986 23980 13874
rect 24136 13870 24164 15030
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23478 11656 23534 11665
rect 23478 11591 23534 11600
rect 23492 10674 23520 11591
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23386 10024 23442 10033
rect 23386 9959 23442 9968
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22572 8906 22600 9522
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22480 8758 22692 8786
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22388 8498 22416 8570
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22572 8022 22600 8502
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22572 7478 22600 7822
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22282 6352 22338 6361
rect 22282 6287 22338 6296
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22376 6248 22428 6254
rect 22374 6216 22376 6225
rect 22428 6216 22430 6225
rect 22192 6180 22244 6186
rect 22374 6151 22430 6160
rect 22192 6122 22244 6128
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22112 2446 22140 5646
rect 22572 5030 22600 6258
rect 22664 6186 22692 8758
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22756 8090 22784 8434
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22940 7818 22968 8570
rect 23492 7886 23520 9386
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 23124 7342 23152 7822
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22756 6798 22784 7142
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 23032 5914 23060 7278
rect 23124 6254 23152 7278
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 22756 5522 22784 5578
rect 22756 5494 22876 5522
rect 22848 5234 22876 5494
rect 23294 5400 23350 5409
rect 23294 5335 23350 5344
rect 23308 5302 23336 5335
rect 23400 5302 23428 5646
rect 23296 5296 23348 5302
rect 23296 5238 23348 5244
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22204 3602 22232 4966
rect 22664 4826 22692 5170
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22848 4758 22876 5170
rect 23676 4758 23704 11290
rect 23952 10266 23980 12922
rect 24504 11830 24532 16050
rect 24596 14362 24624 16068
rect 24728 16079 24730 16088
rect 25688 16108 25740 16114
rect 24676 16050 24728 16056
rect 25688 16050 25740 16056
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24688 15434 24716 15846
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24688 14550 24716 15370
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24780 14550 24808 14962
rect 24676 14544 24728 14550
rect 24676 14486 24728 14492
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24964 14414 24992 15370
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25320 14884 25372 14890
rect 25320 14826 25372 14832
rect 24952 14408 25004 14414
rect 24596 14334 24716 14362
rect 24952 14350 25004 14356
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24596 12442 24624 12786
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24688 11286 24716 14334
rect 25332 14278 25360 14826
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24872 12986 24900 13874
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24872 12238 24900 12922
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 25056 12238 25084 12650
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 25056 11150 25084 12174
rect 25228 12164 25280 12170
rect 25228 12106 25280 12112
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 24780 10742 24808 10950
rect 25148 10810 25176 10950
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 25148 10674 25176 10746
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24596 10266 24624 10406
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24688 10062 24716 10610
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24688 9450 24716 9998
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 24676 9444 24728 9450
rect 24676 9386 24728 9392
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24688 6866 24716 7346
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23848 5296 23900 5302
rect 23848 5238 23900 5244
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22204 3058 22232 3538
rect 23676 3534 23704 4694
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23768 4486 23796 4626
rect 23860 4622 23888 5238
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 4146 23796 4422
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23860 4078 23888 4558
rect 23952 4554 23980 5306
rect 24504 5234 24532 6734
rect 25056 6225 25084 9930
rect 25240 6304 25268 12106
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25332 10130 25360 11018
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25332 9586 25360 10066
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25332 8378 25360 8978
rect 25424 8498 25452 9318
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25332 8350 25452 8378
rect 25424 6322 25452 8350
rect 25320 6316 25372 6322
rect 25240 6276 25320 6304
rect 25320 6258 25372 6264
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25042 6216 25098 6225
rect 25042 6151 25098 6160
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 25148 5710 25176 6054
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 25332 5642 25360 6258
rect 25320 5636 25372 5642
rect 25320 5578 25372 5584
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 23940 4548 23992 4554
rect 23940 4490 23992 4496
rect 24044 4298 24072 5170
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 23952 4270 24072 4298
rect 23952 4146 23980 4270
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 21916 1352 21968 1358
rect 21916 1294 21968 1300
rect 22020 898 22048 2314
rect 22480 2106 22508 2450
rect 22468 2100 22520 2106
rect 22468 2042 22520 2048
rect 22020 870 22140 898
rect 22112 800 22140 870
rect 22572 800 22600 3402
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23584 3058 23612 3334
rect 23860 3194 23888 3402
rect 23952 3194 23980 4082
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24044 3534 24072 3878
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 24872 3074 24900 4150
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 24780 3046 24900 3074
rect 24952 3052 25004 3058
rect 24780 2582 24808 3046
rect 24952 2994 25004 3000
rect 24860 2984 24912 2990
rect 24964 2961 24992 2994
rect 24860 2926 24912 2932
rect 24950 2952 25006 2961
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 23032 800 23060 2314
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23492 1970 23520 2246
rect 23480 1964 23532 1970
rect 23480 1906 23532 1912
rect 23952 800 23980 2382
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 24412 800 24440 2314
rect 24872 800 24900 2926
rect 24950 2887 25006 2896
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 24964 2582 24992 2790
rect 24952 2576 25004 2582
rect 24952 2518 25004 2524
rect 25148 2514 25176 4762
rect 25424 3398 25452 6258
rect 25516 5778 25544 14962
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25608 11626 25636 11766
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25700 10810 25728 11630
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25792 8294 25820 12786
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25976 11898 26004 12038
rect 25964 11892 26016 11898
rect 25964 11834 26016 11840
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 25976 8974 26004 11630
rect 26160 10062 26188 16050
rect 27540 15570 27568 16390
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26700 15496 26752 15502
rect 26700 15438 26752 15444
rect 26240 14544 26292 14550
rect 26240 14486 26292 14492
rect 26252 14414 26280 14486
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26344 12918 26372 15438
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26436 12986 26464 14962
rect 26712 14550 26740 15438
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 26700 14544 26752 14550
rect 26700 14486 26752 14492
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26620 14278 26648 14350
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26712 13530 26740 14486
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26332 12912 26384 12918
rect 26332 12854 26384 12860
rect 26344 12306 26372 12854
rect 26896 12714 26924 14418
rect 27252 14272 27304 14278
rect 27252 14214 27304 14220
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26332 12300 26384 12306
rect 26332 12242 26384 12248
rect 26148 10056 26200 10062
rect 26148 9998 26200 10004
rect 26344 9926 26372 12242
rect 26804 12238 26832 12582
rect 26988 12238 27016 13466
rect 27264 13326 27292 14214
rect 27252 13320 27304 13326
rect 27080 13280 27252 13308
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26424 9716 26476 9722
rect 26424 9658 26476 9664
rect 26240 9580 26292 9586
rect 26292 9540 26372 9568
rect 26240 9522 26292 9528
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 25872 8492 25924 8498
rect 25872 8434 25924 8440
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25884 7954 25912 8434
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 25516 5234 25544 5714
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25608 5098 25636 6258
rect 25884 5778 25912 7890
rect 26160 7886 26188 8774
rect 26252 8090 26280 8774
rect 26344 8362 26372 9540
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 26148 6384 26200 6390
rect 26148 6326 26200 6332
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25596 5092 25648 5098
rect 25596 5034 25648 5040
rect 25884 4690 25912 5714
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 25884 3534 25912 4626
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 25884 3126 25912 3470
rect 26160 3194 26188 6326
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 25884 2990 25912 3062
rect 25872 2984 25924 2990
rect 25872 2926 25924 2932
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25320 2372 25372 2378
rect 25320 2314 25372 2320
rect 26240 2372 26292 2378
rect 26240 2314 26292 2320
rect 25332 800 25360 2314
rect 26252 800 26280 2314
rect 26344 2310 26372 8298
rect 26436 6798 26464 9658
rect 26620 9586 26648 11086
rect 26712 10266 26740 12174
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26712 9654 26740 10202
rect 27080 10062 27108 13280
rect 27252 13262 27304 13268
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27172 12306 27200 12786
rect 27356 12434 27384 14894
rect 27540 14346 27568 15370
rect 27632 14958 27660 17818
rect 28080 17808 28132 17814
rect 28080 17750 28132 17756
rect 27896 16992 27948 16998
rect 27896 16934 27948 16940
rect 27908 16590 27936 16934
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27804 15632 27856 15638
rect 27804 15574 27856 15580
rect 27712 15360 27764 15366
rect 27712 15302 27764 15308
rect 27620 14952 27672 14958
rect 27620 14894 27672 14900
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27540 14074 27568 14282
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27448 12986 27476 13126
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27356 12406 27476 12434
rect 27252 12368 27304 12374
rect 27252 12310 27304 12316
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27264 11762 27292 12310
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27160 11688 27212 11694
rect 27158 11656 27160 11665
rect 27212 11656 27214 11665
rect 27158 11591 27214 11600
rect 27356 10062 27384 12174
rect 27068 10056 27120 10062
rect 27068 9998 27120 10004
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27080 9722 27108 9998
rect 27068 9716 27120 9722
rect 27068 9658 27120 9664
rect 26700 9648 26752 9654
rect 26700 9590 26752 9596
rect 26608 9580 26660 9586
rect 26608 9522 26660 9528
rect 26620 9042 26648 9522
rect 27356 9518 27384 9998
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26620 6118 26648 8842
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27356 7546 27384 8026
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 26620 5914 26648 6054
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 27356 5370 27384 5510
rect 27344 5364 27396 5370
rect 27344 5306 27396 5312
rect 27356 5234 27384 5306
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27448 4185 27476 12406
rect 27526 6216 27582 6225
rect 27526 6151 27582 6160
rect 27540 5370 27568 6151
rect 27632 5370 27660 14758
rect 27724 14482 27752 15302
rect 27816 15026 27844 15574
rect 28092 15434 28120 17750
rect 29196 17202 29224 19314
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 28172 17128 28224 17134
rect 28172 17070 28224 17076
rect 28184 16726 28212 17070
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28920 16794 28948 16934
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28172 16720 28224 16726
rect 28172 16662 28224 16668
rect 29092 16652 29144 16658
rect 29092 16594 29144 16600
rect 29104 15706 29132 16594
rect 29196 16590 29224 17138
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29196 16182 29224 16526
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 28080 15428 28132 15434
rect 28080 15370 28132 15376
rect 28092 15094 28120 15370
rect 28080 15088 28132 15094
rect 28080 15030 28132 15036
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28632 14884 28684 14890
rect 28632 14826 28684 14832
rect 28644 14550 28672 14826
rect 28632 14544 28684 14550
rect 28632 14486 28684 14492
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27724 14278 27752 14418
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27908 13326 27936 14282
rect 28264 13728 28316 13734
rect 28264 13670 28316 13676
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27908 12442 27936 13262
rect 27988 13252 28040 13258
rect 27988 13194 28040 13200
rect 28000 12442 28028 13194
rect 28276 12850 28304 13670
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 27988 12436 28040 12442
rect 28276 12434 28304 12786
rect 28276 12406 28396 12434
rect 27988 12378 28040 12384
rect 28368 12238 28396 12406
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28448 12232 28500 12238
rect 28448 12174 28500 12180
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27724 9994 27752 11290
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27724 9586 27752 9930
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27528 5364 27580 5370
rect 27528 5306 27580 5312
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27528 5226 27580 5232
rect 27528 5168 27580 5174
rect 27434 4176 27490 4185
rect 27434 4111 27490 4120
rect 27540 4026 27568 5168
rect 27448 3998 27568 4026
rect 27160 3664 27212 3670
rect 27160 3606 27212 3612
rect 26700 2372 26752 2378
rect 26700 2314 26752 2320
rect 26332 2304 26384 2310
rect 26332 2246 26384 2252
rect 26712 800 26740 2314
rect 27172 1970 27200 3606
rect 27448 2582 27476 3998
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 3602 27660 3878
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27816 3194 27844 9522
rect 28092 9450 28120 11494
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28080 9444 28132 9450
rect 28080 9386 28132 9392
rect 27894 5400 27950 5409
rect 27894 5335 27896 5344
rect 27948 5335 27950 5344
rect 27896 5306 27948 5312
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 27160 1964 27212 1970
rect 27160 1906 27212 1912
rect 27540 898 27568 2994
rect 28276 2446 28304 11086
rect 28368 9654 28396 12174
rect 28460 11898 28488 12174
rect 28644 12170 28672 14486
rect 29012 14482 29040 14962
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28828 12850 28856 14214
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 29012 13394 29040 13738
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28816 12708 28868 12714
rect 28816 12650 28868 12656
rect 28828 12238 28856 12650
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28540 12164 28592 12170
rect 28540 12106 28592 12112
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28724 12164 28776 12170
rect 28724 12106 28776 12112
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28552 11762 28580 12106
rect 28540 11756 28592 11762
rect 28540 11698 28592 11704
rect 28644 11354 28672 12106
rect 28632 11348 28684 11354
rect 28632 11290 28684 11296
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28644 9450 28672 9522
rect 28632 9444 28684 9450
rect 28632 9386 28684 9392
rect 28644 9178 28672 9386
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 28540 4004 28592 4010
rect 28540 3946 28592 3952
rect 28552 3534 28580 3946
rect 28736 3738 28764 12106
rect 28828 9654 28856 12174
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 28920 11150 28948 12106
rect 29380 11898 29408 19314
rect 29472 17202 29500 24278
rect 29748 23322 29776 24618
rect 30208 23730 30236 25842
rect 30300 24818 30328 25910
rect 30840 25764 30892 25770
rect 30840 25706 30892 25712
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30392 24818 30420 25094
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 30024 22778 30052 23054
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 30208 22438 30236 23666
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30484 22250 30512 23666
rect 30576 23254 30604 24006
rect 30564 23248 30616 23254
rect 30564 23190 30616 23196
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30564 22432 30616 22438
rect 30564 22374 30616 22380
rect 30300 22234 30512 22250
rect 30288 22228 30512 22234
rect 30340 22222 30512 22228
rect 30288 22170 30340 22176
rect 30196 22024 30248 22030
rect 30196 21966 30248 21972
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 29748 21622 29776 21830
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 30116 21350 30144 21830
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29840 19378 29868 20198
rect 29932 19854 29960 20334
rect 30024 20262 30052 20402
rect 30208 20398 30236 21966
rect 30484 21894 30512 22222
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30576 21078 30604 22374
rect 30668 22166 30696 23054
rect 30852 22234 30880 25706
rect 31760 24268 31812 24274
rect 31760 24210 31812 24216
rect 31772 23866 31800 24210
rect 31760 23860 31812 23866
rect 31760 23802 31812 23808
rect 31760 23656 31812 23662
rect 31760 23598 31812 23604
rect 31208 23588 31260 23594
rect 31208 23530 31260 23536
rect 30840 22228 30892 22234
rect 30840 22170 30892 22176
rect 30656 22160 30708 22166
rect 30656 22102 30708 22108
rect 30668 21554 30696 22102
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30760 21842 30788 21898
rect 30760 21814 30880 21842
rect 30852 21622 30880 21814
rect 30840 21616 30892 21622
rect 30840 21558 30892 21564
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30852 21486 30880 21558
rect 31220 21486 31248 23530
rect 31392 23044 31444 23050
rect 31392 22986 31444 22992
rect 30840 21480 30892 21486
rect 30840 21422 30892 21428
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 30564 21072 30616 21078
rect 30564 21014 30616 21020
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30012 20256 30064 20262
rect 30012 20198 30064 20204
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 30024 19786 30052 20198
rect 30012 19780 30064 19786
rect 30012 19722 30064 19728
rect 30104 19780 30156 19786
rect 30104 19722 30156 19728
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 30116 18834 30144 19722
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30300 19530 30328 19654
rect 30300 19502 30420 19530
rect 30392 19446 30420 19502
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 30380 19440 30432 19446
rect 30380 19382 30432 19388
rect 30104 18828 30156 18834
rect 30104 18770 30156 18776
rect 30116 18698 30144 18770
rect 30104 18692 30156 18698
rect 30300 18680 30328 19382
rect 30380 18692 30432 18698
rect 30300 18652 30380 18680
rect 30104 18634 30156 18640
rect 30380 18634 30432 18640
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29472 15473 29500 16050
rect 29932 15502 29960 16050
rect 29920 15496 29972 15502
rect 29458 15464 29514 15473
rect 29920 15438 29972 15444
rect 29458 15399 29514 15408
rect 29368 11892 29420 11898
rect 29368 11834 29420 11840
rect 29472 11762 29500 15399
rect 29932 15026 29960 15438
rect 29920 15020 29972 15026
rect 29920 14962 29972 14968
rect 30116 14414 30144 18634
rect 30392 18222 30420 18634
rect 30484 18442 30512 20878
rect 30576 20874 30604 21014
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30484 18414 30604 18442
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30392 17270 30420 18158
rect 30484 17746 30512 18226
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30380 17264 30432 17270
rect 30380 17206 30432 17212
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30196 15904 30248 15910
rect 30196 15846 30248 15852
rect 30208 15502 30236 15846
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30300 15178 30328 17138
rect 30392 16794 30420 17206
rect 30472 17128 30524 17134
rect 30472 17070 30524 17076
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30484 16182 30512 17070
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30300 15150 30420 15178
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29828 14340 29880 14346
rect 29828 14282 29880 14288
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28920 8906 28948 9998
rect 29012 9994 29040 11698
rect 29748 11354 29776 11698
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29644 11008 29696 11014
rect 29644 10950 29696 10956
rect 29656 10674 29684 10950
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 29012 9654 29040 9930
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 29276 8900 29328 8906
rect 29276 8842 29328 8848
rect 29288 6798 29316 8842
rect 29656 8838 29684 10610
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29288 5914 29316 6734
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29288 5234 29316 5850
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28920 3670 28948 4014
rect 29288 3942 29316 5170
rect 29368 4276 29420 4282
rect 29368 4218 29420 4224
rect 29380 4146 29408 4218
rect 29368 4140 29420 4146
rect 29368 4082 29420 4088
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29276 3936 29328 3942
rect 29276 3878 29328 3884
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28920 3534 28948 3606
rect 29472 3602 29500 4082
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28080 2372 28132 2378
rect 28080 2314 28132 2320
rect 27540 870 27660 898
rect 27632 800 27660 870
rect 28092 800 28120 2314
rect 29012 800 29040 3130
rect 29656 2446 29684 8774
rect 29748 6390 29776 8910
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 29736 5636 29788 5642
rect 29736 5578 29788 5584
rect 29748 5030 29776 5578
rect 29736 5024 29788 5030
rect 29736 4966 29788 4972
rect 29840 4826 29868 14282
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 29932 13530 29960 13874
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 30012 12096 30064 12102
rect 30012 12038 30064 12044
rect 30024 11898 30052 12038
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 30012 11212 30064 11218
rect 30012 11154 30064 11160
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29932 10810 29960 11018
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 30024 10606 30052 11154
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 30024 9722 30052 10542
rect 30116 10062 30144 14350
rect 30208 14074 30236 14758
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30288 14000 30340 14006
rect 30288 13942 30340 13948
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 30116 9654 30144 9998
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 29932 6390 29960 6734
rect 29920 6384 29972 6390
rect 29920 6326 29972 6332
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29840 4146 29868 4762
rect 29932 4729 29960 6054
rect 30024 5302 30052 6802
rect 30104 6792 30156 6798
rect 30102 6760 30104 6769
rect 30156 6760 30158 6769
rect 30102 6695 30158 6704
rect 30012 5296 30064 5302
rect 30012 5238 30064 5244
rect 30116 5234 30144 6695
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 30024 4826 30052 5102
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 29918 4720 29974 4729
rect 29918 4655 29920 4664
rect 29972 4655 29974 4664
rect 29920 4626 29972 4632
rect 30012 4548 30064 4554
rect 30012 4490 30064 4496
rect 30024 4146 30052 4490
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 30116 4078 30144 5170
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 29918 3904 29974 3913
rect 29918 3839 29974 3848
rect 29932 3466 29960 3839
rect 30116 3670 30144 4014
rect 30104 3664 30156 3670
rect 30104 3606 30156 3612
rect 29920 3460 29972 3466
rect 29920 3402 29972 3408
rect 30012 3392 30064 3398
rect 30012 3334 30064 3340
rect 30024 3194 30052 3334
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 30024 3097 30052 3130
rect 30010 3088 30066 3097
rect 30010 3023 30066 3032
rect 30208 2582 30236 13330
rect 30300 11830 30328 13942
rect 30288 11824 30340 11830
rect 30288 11766 30340 11772
rect 30300 10130 30328 11766
rect 30392 11694 30420 15150
rect 30576 14414 30604 18414
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30668 17882 30696 18226
rect 30656 17876 30708 17882
rect 30656 17818 30708 17824
rect 30656 17604 30708 17610
rect 30656 17546 30708 17552
rect 30668 17134 30696 17546
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 30852 16946 30880 21422
rect 31220 21078 31248 21422
rect 31208 21072 31260 21078
rect 31208 21014 31260 21020
rect 30932 21004 30984 21010
rect 30932 20946 30984 20952
rect 30944 19922 30972 20946
rect 31404 20942 31432 22986
rect 31772 22778 31800 23598
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31024 20936 31076 20942
rect 31392 20936 31444 20942
rect 31076 20884 31392 20890
rect 31024 20878 31444 20884
rect 31036 20862 31432 20878
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 31392 19304 31444 19310
rect 31392 19246 31444 19252
rect 31208 19168 31260 19174
rect 31208 19110 31260 19116
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31036 18290 31064 18702
rect 31024 18284 31076 18290
rect 31024 18226 31076 18232
rect 31128 17610 31156 18702
rect 31220 18698 31248 19110
rect 31404 18970 31432 19246
rect 31392 18964 31444 18970
rect 31392 18906 31444 18912
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 31392 18148 31444 18154
rect 31392 18090 31444 18096
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 31312 17746 31340 18022
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 30668 16918 30880 16946
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30484 13870 30512 14214
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30576 13530 30604 14214
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30668 12170 30696 16918
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 16114 30788 16390
rect 31024 16244 31076 16250
rect 31024 16186 31076 16192
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30760 15570 30788 16050
rect 31036 15638 31064 16186
rect 31024 15632 31076 15638
rect 31024 15574 31076 15580
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30748 14408 30800 14414
rect 30748 14350 30800 14356
rect 30760 14074 30788 14350
rect 30748 14068 30800 14074
rect 30748 14010 30800 14016
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30380 11688 30432 11694
rect 30380 11630 30432 11636
rect 30380 10804 30432 10810
rect 30380 10746 30432 10752
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 30300 8974 30328 10066
rect 30288 8968 30340 8974
rect 30288 8910 30340 8916
rect 30392 7410 30420 10746
rect 30668 9178 30696 12106
rect 30656 9172 30708 9178
rect 30656 9114 30708 9120
rect 30760 8022 30788 13262
rect 31036 12434 31064 15574
rect 31312 15026 31340 16730
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31300 15020 31352 15026
rect 31300 14962 31352 14968
rect 31220 12442 31248 14962
rect 31404 14482 31432 18090
rect 31392 14476 31444 14482
rect 31392 14418 31444 14424
rect 31496 13734 31524 22170
rect 31956 19446 31984 28358
rect 32496 26444 32548 26450
rect 32496 26386 32548 26392
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32140 25906 32168 26318
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32140 23118 32168 25842
rect 32220 24608 32272 24614
rect 32324 24596 32352 26318
rect 32508 25906 32536 26386
rect 32680 26308 32732 26314
rect 32680 26250 32732 26256
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32508 24970 32536 25842
rect 32272 24568 32352 24596
rect 32220 24550 32272 24556
rect 32324 23730 32352 24568
rect 32416 24942 32536 24970
rect 32416 24342 32444 24942
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 32404 24336 32456 24342
rect 32404 24278 32456 24284
rect 32508 23866 32536 24754
rect 32600 24274 32628 24754
rect 32588 24268 32640 24274
rect 32588 24210 32640 24216
rect 32496 23860 32548 23866
rect 32496 23802 32548 23808
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32324 23526 32352 23666
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 32312 22432 32364 22438
rect 32312 22374 32364 22380
rect 32036 20392 32088 20398
rect 32036 20334 32088 20340
rect 31944 19440 31996 19446
rect 31944 19382 31996 19388
rect 31576 19236 31628 19242
rect 31576 19178 31628 19184
rect 31588 18766 31616 19178
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 32048 18698 32076 20334
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 31588 18290 31892 18306
rect 31576 18284 31892 18290
rect 31628 18278 31892 18284
rect 31576 18226 31628 18232
rect 31864 18086 31892 18278
rect 31852 18080 31904 18086
rect 31852 18022 31904 18028
rect 32048 17610 32076 18634
rect 32036 17604 32088 17610
rect 32036 17546 32088 17552
rect 32324 17202 32352 22374
rect 32494 19680 32550 19689
rect 32494 19615 32550 19624
rect 32508 19514 32536 19615
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32036 13796 32088 13802
rect 32036 13738 32088 13744
rect 31484 13728 31536 13734
rect 31484 13670 31536 13676
rect 32048 13326 32076 13738
rect 32036 13320 32088 13326
rect 32036 13262 32088 13268
rect 31852 13252 31904 13258
rect 31852 13194 31904 13200
rect 31576 13184 31628 13190
rect 31576 13126 31628 13132
rect 31588 12850 31616 13126
rect 31864 12986 31892 13194
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 31300 12776 31352 12782
rect 31300 12718 31352 12724
rect 31208 12436 31260 12442
rect 31036 12406 31156 12434
rect 31024 11008 31076 11014
rect 31024 10950 31076 10956
rect 31036 10742 31064 10950
rect 31024 10736 31076 10742
rect 31024 10678 31076 10684
rect 31128 10690 31156 12406
rect 31208 12378 31260 12384
rect 31220 12306 31248 12378
rect 31208 12300 31260 12306
rect 31208 12242 31260 12248
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30748 8016 30800 8022
rect 30748 7958 30800 7964
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30300 6118 30328 6734
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 6322 30512 6598
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30656 6248 30708 6254
rect 30656 6190 30708 6196
rect 30288 6112 30340 6118
rect 30288 6054 30340 6060
rect 30668 5914 30696 6190
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30288 5568 30340 5574
rect 30288 5510 30340 5516
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30300 5370 30328 5510
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 30392 5234 30420 5510
rect 30380 5228 30432 5234
rect 30380 5170 30432 5176
rect 30392 4214 30420 5170
rect 30760 4282 30788 7958
rect 30852 7342 30880 9522
rect 30840 7336 30892 7342
rect 30840 7278 30892 7284
rect 30852 6798 30880 7278
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30840 4480 30892 4486
rect 30840 4422 30892 4428
rect 30852 4282 30880 4422
rect 30748 4276 30800 4282
rect 30748 4218 30800 4224
rect 30840 4276 30892 4282
rect 30840 4218 30892 4224
rect 30380 4208 30432 4214
rect 30380 4150 30432 4156
rect 30760 3534 30788 4218
rect 30932 3732 30984 3738
rect 30932 3674 30984 3680
rect 30944 3534 30972 3674
rect 30564 3528 30616 3534
rect 30564 3470 30616 3476
rect 30748 3528 30800 3534
rect 30932 3528 30984 3534
rect 30748 3470 30800 3476
rect 30852 3488 30932 3516
rect 30288 3460 30340 3466
rect 30288 3402 30340 3408
rect 30472 3460 30524 3466
rect 30472 3402 30524 3408
rect 30196 2576 30248 2582
rect 30196 2518 30248 2524
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29460 2372 29512 2378
rect 29460 2314 29512 2320
rect 29472 800 29500 2314
rect 30300 898 30328 3402
rect 30484 3194 30512 3402
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30484 2106 30512 3130
rect 30576 3058 30604 3470
rect 30564 3052 30616 3058
rect 30564 2994 30616 3000
rect 30748 3050 30800 3056
rect 30852 3040 30880 3488
rect 30932 3470 30984 3476
rect 30800 3012 30880 3040
rect 30748 2992 30800 2998
rect 30748 2916 30800 2922
rect 30748 2858 30800 2864
rect 30472 2100 30524 2106
rect 30472 2042 30524 2048
rect 30760 1902 30788 2858
rect 31036 2774 31064 10678
rect 31128 10662 31248 10690
rect 31312 10674 31340 12718
rect 31852 12640 31904 12646
rect 31852 12582 31904 12588
rect 31864 12238 31892 12582
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31852 12232 31904 12238
rect 31852 12174 31904 12180
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 31220 10606 31248 10662
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 31312 10198 31340 10610
rect 31300 10192 31352 10198
rect 31300 10134 31352 10140
rect 31496 9586 31524 11494
rect 31668 10668 31720 10674
rect 31668 10610 31720 10616
rect 31576 9920 31628 9926
rect 31576 9862 31628 9868
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31392 8968 31444 8974
rect 31392 8910 31444 8916
rect 31300 7404 31352 7410
rect 31300 7346 31352 7352
rect 31208 6792 31260 6798
rect 31208 6734 31260 6740
rect 31220 4622 31248 6734
rect 31208 4616 31260 4622
rect 31208 4558 31260 4564
rect 31312 4468 31340 7346
rect 31404 6798 31432 8910
rect 31496 8906 31524 9318
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31588 7886 31616 9862
rect 31680 7886 31708 10610
rect 31772 10130 31800 12174
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 31956 10062 31984 10406
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31760 9920 31812 9926
rect 31760 9862 31812 9868
rect 31772 9586 31800 9862
rect 31852 9716 31904 9722
rect 31852 9658 31904 9664
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31864 8566 31892 9658
rect 32128 9580 32180 9586
rect 32128 9522 32180 9528
rect 31944 9512 31996 9518
rect 31944 9454 31996 9460
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 31760 8424 31812 8430
rect 31760 8366 31812 8372
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31772 6866 31800 8366
rect 31760 6860 31812 6866
rect 31760 6802 31812 6808
rect 31392 6792 31444 6798
rect 31392 6734 31444 6740
rect 31220 4440 31340 4468
rect 31220 4146 31248 4440
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31220 3913 31248 4082
rect 31206 3904 31262 3913
rect 31206 3839 31262 3848
rect 31208 3460 31260 3466
rect 31312 3448 31340 4082
rect 31404 3738 31432 6734
rect 31760 4208 31812 4214
rect 31864 4196 31892 8502
rect 31956 8498 31984 9454
rect 32140 8838 32168 9522
rect 32220 9512 32272 9518
rect 32324 9466 32352 17138
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 32272 9460 32352 9466
rect 32220 9454 32352 9460
rect 32232 9438 32352 9454
rect 32232 8906 32260 9438
rect 32220 8900 32272 8906
rect 32220 8842 32272 8848
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 32140 8498 32168 8774
rect 31944 8492 31996 8498
rect 31944 8434 31996 8440
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 31956 6662 31984 8434
rect 32416 7954 32444 15642
rect 32508 13258 32536 19314
rect 32600 18970 32628 19450
rect 32588 18964 32640 18970
rect 32588 18906 32640 18912
rect 32600 18766 32628 18906
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32692 18358 32720 26250
rect 32956 25356 33008 25362
rect 32956 25298 33008 25304
rect 32968 24206 32996 25298
rect 33048 24812 33100 24818
rect 33048 24754 33100 24760
rect 32956 24200 33008 24206
rect 32956 24142 33008 24148
rect 32968 22030 32996 24142
rect 33060 23594 33088 24754
rect 33140 24608 33192 24614
rect 33140 24550 33192 24556
rect 33152 24206 33180 24550
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33048 23588 33100 23594
rect 33048 23530 33100 23536
rect 33060 23322 33088 23530
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 32864 21684 32916 21690
rect 32864 21626 32916 21632
rect 32876 21350 32904 21626
rect 32864 21344 32916 21350
rect 32864 21286 32916 21292
rect 32772 19372 32824 19378
rect 32772 19314 32824 19320
rect 32680 18352 32732 18358
rect 32680 18294 32732 18300
rect 32692 17202 32720 18294
rect 32784 18290 32812 19314
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32876 18170 32904 21286
rect 32968 21010 32996 21966
rect 32956 21004 33008 21010
rect 32956 20946 33008 20952
rect 32784 18142 32904 18170
rect 32680 17196 32732 17202
rect 32680 17138 32732 17144
rect 32588 17060 32640 17066
rect 32588 17002 32640 17008
rect 32600 16794 32628 17002
rect 32588 16788 32640 16794
rect 32588 16730 32640 16736
rect 32496 13252 32548 13258
rect 32496 13194 32548 13200
rect 32496 12232 32548 12238
rect 32496 12174 32548 12180
rect 32508 10690 32536 12174
rect 32784 11150 32812 18142
rect 33140 16108 33192 16114
rect 33140 16050 33192 16056
rect 33048 15700 33100 15706
rect 33048 15642 33100 15648
rect 33060 15094 33088 15642
rect 33152 15502 33180 16050
rect 33140 15496 33192 15502
rect 33140 15438 33192 15444
rect 33048 15088 33100 15094
rect 33048 15030 33100 15036
rect 33152 13938 33180 15438
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 32864 13796 32916 13802
rect 32864 13738 32916 13744
rect 32876 11762 32904 13738
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 33152 12102 33180 12786
rect 33140 12096 33192 12102
rect 33140 12038 33192 12044
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32876 11150 32904 11698
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 32864 11144 32916 11150
rect 32864 11086 32916 11092
rect 32588 11076 32640 11082
rect 32588 11018 32640 11024
rect 32600 10810 32628 11018
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32508 10662 32628 10690
rect 32496 10600 32548 10606
rect 32496 10542 32548 10548
rect 32508 8430 32536 10542
rect 32496 8424 32548 8430
rect 32496 8366 32548 8372
rect 32404 7948 32456 7954
rect 32404 7890 32456 7896
rect 32404 7812 32456 7818
rect 32404 7754 32456 7760
rect 32416 7546 32444 7754
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32402 7440 32458 7449
rect 32402 7375 32404 7384
rect 32456 7375 32458 7384
rect 32404 7346 32456 7352
rect 32036 7200 32088 7206
rect 32036 7142 32088 7148
rect 32048 6798 32076 7142
rect 32508 6798 32536 8366
rect 32036 6792 32088 6798
rect 32496 6792 32548 6798
rect 32036 6734 32088 6740
rect 32310 6760 32366 6769
rect 32496 6734 32548 6740
rect 32310 6695 32312 6704
rect 32364 6695 32366 6704
rect 32312 6666 32364 6672
rect 31944 6656 31996 6662
rect 32600 6610 32628 10662
rect 32876 9110 32904 11086
rect 33244 11082 33272 35866
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 33784 27056 33836 27062
rect 33784 26998 33836 27004
rect 33508 26512 33560 26518
rect 33508 26454 33560 26460
rect 33520 25906 33548 26454
rect 33692 26308 33744 26314
rect 33692 26250 33744 26256
rect 33704 25906 33732 26250
rect 33508 25900 33560 25906
rect 33508 25842 33560 25848
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 33336 23118 33364 23598
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33324 21956 33376 21962
rect 33324 21898 33376 21904
rect 33336 21690 33364 21898
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 33520 21554 33548 24822
rect 33796 24682 33824 26998
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34152 26920 34204 26926
rect 34152 26862 34204 26868
rect 34164 26382 34192 26862
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34440 26382 34468 26726
rect 34152 26376 34204 26382
rect 34152 26318 34204 26324
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 34624 25498 34652 26930
rect 36360 26920 36412 26926
rect 36360 26862 36412 26868
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 34808 26466 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34808 26438 34928 26466
rect 34900 26330 34928 26438
rect 35256 26376 35308 26382
rect 34900 26314 35020 26330
rect 35256 26318 35308 26324
rect 34796 26308 34848 26314
rect 34796 26250 34848 26256
rect 34900 26308 35032 26314
rect 34900 26302 34980 26308
rect 34612 25492 34664 25498
rect 34612 25434 34664 25440
rect 34624 24886 34652 25434
rect 34612 24880 34664 24886
rect 34612 24822 34664 24828
rect 34428 24812 34480 24818
rect 34428 24754 34480 24760
rect 33784 24676 33836 24682
rect 33784 24618 33836 24624
rect 33600 21888 33652 21894
rect 33600 21830 33652 21836
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 33508 21548 33560 21554
rect 33508 21490 33560 21496
rect 33520 19922 33548 21490
rect 33612 20874 33640 21830
rect 34348 21690 34376 21830
rect 34336 21684 34388 21690
rect 34336 21626 34388 21632
rect 34440 21554 34468 24754
rect 34808 24138 34836 26250
rect 34900 26042 34928 26302
rect 34980 26250 35032 26256
rect 34888 26036 34940 26042
rect 34888 25978 34940 25984
rect 35268 25906 35296 26318
rect 35256 25900 35308 25906
rect 35256 25842 35308 25848
rect 35268 25770 35296 25842
rect 35256 25764 35308 25770
rect 35256 25706 35308 25712
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35716 24676 35768 24682
rect 35716 24618 35768 24624
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24132 34848 24138
rect 34796 24074 34848 24080
rect 34612 24064 34664 24070
rect 34612 24006 34664 24012
rect 34624 23730 34652 24006
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34532 21622 34560 22986
rect 34520 21616 34572 21622
rect 34520 21558 34572 21564
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33876 21548 33928 21554
rect 33876 21490 33928 21496
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 33600 20868 33652 20874
rect 33600 20810 33652 20816
rect 33796 20398 33824 21490
rect 33888 20602 33916 21490
rect 34336 21480 34388 21486
rect 34336 21422 34388 21428
rect 34348 20942 34376 21422
rect 34336 20936 34388 20942
rect 34336 20878 34388 20884
rect 33876 20596 33928 20602
rect 33876 20538 33928 20544
rect 34520 20528 34572 20534
rect 34520 20470 34572 20476
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 34428 20256 34480 20262
rect 34428 20198 34480 20204
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33520 19242 33548 19858
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 34348 19446 34376 19654
rect 34336 19440 34388 19446
rect 34440 19417 34468 20198
rect 34532 19854 34560 20470
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 34336 19382 34388 19388
rect 34426 19408 34482 19417
rect 34426 19343 34482 19352
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 33508 19236 33560 19242
rect 33508 19178 33560 19184
rect 33520 17202 33548 19178
rect 34152 18216 34204 18222
rect 34152 18158 34204 18164
rect 33876 17604 33928 17610
rect 33876 17546 33928 17552
rect 33888 17338 33916 17546
rect 34164 17338 34192 18158
rect 33692 17332 33744 17338
rect 33692 17274 33744 17280
rect 33876 17332 33928 17338
rect 33876 17274 33928 17280
rect 34152 17332 34204 17338
rect 34152 17274 34204 17280
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33324 16992 33376 16998
rect 33324 16934 33376 16940
rect 33336 16658 33364 16934
rect 33324 16652 33376 16658
rect 33324 16594 33376 16600
rect 33704 16250 33732 17274
rect 34152 16720 34204 16726
rect 34152 16662 34204 16668
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33784 16176 33836 16182
rect 33784 16118 33836 16124
rect 33796 15706 33824 16118
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 34060 16108 34112 16114
rect 34060 16050 34112 16056
rect 33888 15910 33916 16050
rect 33876 15904 33928 15910
rect 33876 15846 33928 15852
rect 33784 15700 33836 15706
rect 33784 15642 33836 15648
rect 33692 15496 33744 15502
rect 33612 15444 33692 15450
rect 33612 15438 33744 15444
rect 33416 15428 33468 15434
rect 33416 15370 33468 15376
rect 33612 15422 33732 15438
rect 33324 14816 33376 14822
rect 33324 14758 33376 14764
rect 33336 13938 33364 14758
rect 33428 14550 33456 15370
rect 33416 14544 33468 14550
rect 33416 14486 33468 14492
rect 33428 14006 33456 14486
rect 33416 14000 33468 14006
rect 33416 13942 33468 13948
rect 33612 13938 33640 15422
rect 34072 15366 34100 16050
rect 34164 15706 34192 16662
rect 34244 16108 34296 16114
rect 34244 16050 34296 16056
rect 34152 15700 34204 15706
rect 34152 15642 34204 15648
rect 34164 15502 34192 15642
rect 34152 15496 34204 15502
rect 34152 15438 34204 15444
rect 34060 15360 34112 15366
rect 34060 15302 34112 15308
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33796 14074 33824 14554
rect 34256 14278 34284 16050
rect 34244 14272 34296 14278
rect 34244 14214 34296 14220
rect 33784 14068 33836 14074
rect 33784 14010 33836 14016
rect 33324 13932 33376 13938
rect 33324 13874 33376 13880
rect 33508 13932 33560 13938
rect 33508 13874 33560 13880
rect 33600 13932 33652 13938
rect 33600 13874 33652 13880
rect 33324 11756 33376 11762
rect 33324 11698 33376 11704
rect 33232 11076 33284 11082
rect 33232 11018 33284 11024
rect 33048 10532 33100 10538
rect 33048 10474 33100 10480
rect 33060 9382 33088 10474
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 32968 9194 32996 9318
rect 32968 9166 33180 9194
rect 32864 9104 32916 9110
rect 32864 9046 32916 9052
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32876 8566 32904 8910
rect 32864 8560 32916 8566
rect 32864 8502 32916 8508
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 31944 6598 31996 6604
rect 31956 5710 31984 6598
rect 32508 6582 32628 6610
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 31812 4168 31892 4196
rect 31760 4150 31812 4156
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 31484 3664 31536 3670
rect 31484 3606 31536 3612
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 31260 3420 31340 3448
rect 31208 3402 31260 3408
rect 31206 3088 31262 3097
rect 31206 3023 31208 3032
rect 31260 3023 31262 3032
rect 31208 2994 31260 3000
rect 30944 2746 31064 2774
rect 30944 2446 30972 2746
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 30840 2372 30892 2378
rect 30840 2314 30892 2320
rect 30748 1896 30800 1902
rect 30748 1838 30800 1844
rect 30300 870 30420 898
rect 30392 800 30420 870
rect 30852 800 30880 2314
rect 31404 1766 31432 3470
rect 31496 2990 31524 3606
rect 31772 3398 31800 4150
rect 31956 3602 31984 5646
rect 31944 3596 31996 3602
rect 31944 3538 31996 3544
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 32036 3392 32088 3398
rect 32036 3334 32088 3340
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31392 1760 31444 1766
rect 31392 1702 31444 1708
rect 31772 800 31800 2994
rect 32048 2310 32076 3334
rect 32508 2774 32536 6582
rect 32692 6390 32720 7346
rect 32784 7206 32812 8366
rect 32864 7948 32916 7954
rect 32864 7890 32916 7896
rect 32876 7342 32904 7890
rect 33060 7886 33088 8502
rect 33152 7886 33180 9166
rect 33232 8900 33284 8906
rect 33232 8842 33284 8848
rect 33244 8022 33272 8842
rect 33336 8498 33364 11698
rect 33324 8492 33376 8498
rect 33324 8434 33376 8440
rect 33232 8016 33284 8022
rect 33232 7958 33284 7964
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 33140 7880 33192 7886
rect 33140 7822 33192 7828
rect 33232 7812 33284 7818
rect 33232 7754 33284 7760
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 32864 7336 32916 7342
rect 32864 7278 32916 7284
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 32772 7200 32824 7206
rect 32772 7142 32824 7148
rect 32956 7200 33008 7206
rect 32956 7142 33008 7148
rect 32968 7018 32996 7142
rect 32876 6990 32996 7018
rect 32876 6934 32904 6990
rect 32864 6928 32916 6934
rect 32864 6870 32916 6876
rect 32680 6384 32732 6390
rect 32680 6326 32732 6332
rect 32692 6186 32720 6326
rect 32680 6180 32732 6186
rect 32680 6122 32732 6128
rect 33060 5846 33088 7210
rect 33152 6798 33180 7686
rect 33244 7449 33272 7754
rect 33336 7546 33364 8434
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33324 7540 33376 7546
rect 33324 7482 33376 7488
rect 33230 7440 33286 7449
rect 33428 7410 33456 7686
rect 33230 7375 33286 7384
rect 33416 7404 33468 7410
rect 33244 7274 33272 7375
rect 33416 7346 33468 7352
rect 33232 7268 33284 7274
rect 33232 7210 33284 7216
rect 33428 7206 33456 7346
rect 33416 7200 33468 7206
rect 33416 7142 33468 7148
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 33140 6248 33192 6254
rect 33140 6190 33192 6196
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 33152 4078 33180 6190
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 33244 5302 33272 5510
rect 33232 5296 33284 5302
rect 33232 5238 33284 5244
rect 33140 4072 33192 4078
rect 32586 4040 32642 4049
rect 33140 4014 33192 4020
rect 32586 3975 32642 3984
rect 32600 3126 32628 3975
rect 33520 3126 33548 13874
rect 33612 12714 33640 13874
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 34072 12782 34100 12922
rect 34244 12844 34296 12850
rect 34244 12786 34296 12792
rect 34060 12776 34112 12782
rect 34060 12718 34112 12724
rect 33600 12708 33652 12714
rect 33600 12650 33652 12656
rect 33968 11280 34020 11286
rect 33968 11222 34020 11228
rect 33980 10674 34008 11222
rect 33968 10668 34020 10674
rect 33968 10610 34020 10616
rect 33968 10464 34020 10470
rect 33968 10406 34020 10412
rect 33980 9994 34008 10406
rect 33968 9988 34020 9994
rect 33968 9930 34020 9936
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 33876 9920 33928 9926
rect 33928 9868 34008 9874
rect 33876 9862 34008 9868
rect 33704 9586 33732 9862
rect 33888 9846 34008 9862
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33600 8016 33652 8022
rect 33600 7958 33652 7964
rect 33612 6254 33640 7958
rect 33704 7342 33732 9522
rect 33980 9518 34008 9846
rect 34072 9518 34100 12718
rect 34256 12646 34284 12786
rect 34244 12640 34296 12646
rect 34244 12582 34296 12588
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 34060 9512 34112 9518
rect 34060 9454 34112 9460
rect 33876 8288 33928 8294
rect 33876 8230 33928 8236
rect 33784 7812 33836 7818
rect 33784 7754 33836 7760
rect 33692 7336 33744 7342
rect 33692 7278 33744 7284
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 33612 5710 33640 6190
rect 33600 5704 33652 5710
rect 33600 5646 33652 5652
rect 33600 5364 33652 5370
rect 33600 5306 33652 5312
rect 32588 3120 32640 3126
rect 32588 3062 32640 3068
rect 33508 3120 33560 3126
rect 33508 3062 33560 3068
rect 33140 3052 33192 3058
rect 33140 2994 33192 3000
rect 32324 2746 32536 2774
rect 32324 2650 32352 2746
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32036 2304 32088 2310
rect 32036 2246 32088 2252
rect 32232 800 32260 2314
rect 33152 800 33180 2994
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33520 2514 33548 2586
rect 33612 2514 33640 5306
rect 33508 2508 33560 2514
rect 33508 2450 33560 2456
rect 33600 2508 33652 2514
rect 33600 2450 33652 2456
rect 33704 2446 33732 7278
rect 33796 7002 33824 7754
rect 33888 7410 33916 8230
rect 33876 7404 33928 7410
rect 33876 7346 33928 7352
rect 33784 6996 33836 7002
rect 33784 6938 33836 6944
rect 33980 5370 34008 9454
rect 34060 7880 34112 7886
rect 34060 7822 34112 7828
rect 33968 5364 34020 5370
rect 33968 5306 34020 5312
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 33888 3602 33916 5102
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 33888 3058 33916 3538
rect 33980 3058 34008 3878
rect 33876 3052 33928 3058
rect 33876 2994 33928 3000
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 34072 2378 34100 7822
rect 34152 6384 34204 6390
rect 34152 6326 34204 6332
rect 34164 6118 34192 6326
rect 34152 6112 34204 6118
rect 34152 6054 34204 6060
rect 34256 2650 34284 12582
rect 34348 7750 34376 19246
rect 34428 17536 34480 17542
rect 34428 17478 34480 17484
rect 34440 17270 34468 17478
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34532 16522 34560 19314
rect 34624 19242 34652 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34716 20788 34744 21626
rect 34808 21146 34836 21830
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21140 34848 21146
rect 34796 21082 34848 21088
rect 34808 20942 34836 21082
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 34980 20800 35032 20806
rect 34716 20760 34836 20788
rect 34808 20466 34836 20760
rect 34980 20742 35032 20748
rect 34992 20466 35020 20742
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 34980 20460 35032 20466
rect 34980 20402 35032 20408
rect 34716 20262 34744 20402
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34716 19378 34744 20198
rect 34808 19786 34836 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34796 19780 34848 19786
rect 34796 19722 34848 19728
rect 34888 19712 34940 19718
rect 34888 19654 34940 19660
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 34900 19292 34928 19654
rect 35452 19378 35480 23054
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 34808 19264 34928 19292
rect 34612 19236 34664 19242
rect 34612 19178 34664 19184
rect 34808 18698 34836 19264
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18692 34848 18698
rect 34796 18634 34848 18640
rect 34612 17536 34664 17542
rect 34612 17478 34664 17484
rect 34624 16590 34652 17478
rect 34808 17270 34836 18634
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35728 17898 35756 24618
rect 35820 22710 35848 26726
rect 36372 26314 36400 26862
rect 38016 26784 38068 26790
rect 38016 26726 38068 26732
rect 37832 26580 37884 26586
rect 37832 26522 37884 26528
rect 37844 26382 37872 26522
rect 38028 26382 38056 26726
rect 40316 26512 40368 26518
rect 39224 26450 39436 26466
rect 40316 26454 40368 26460
rect 38844 26444 38896 26450
rect 38844 26386 38896 26392
rect 39212 26444 39448 26450
rect 39264 26438 39396 26444
rect 39212 26386 39264 26392
rect 39396 26386 39448 26392
rect 37648 26376 37700 26382
rect 37648 26318 37700 26324
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 38016 26376 38068 26382
rect 38016 26318 38068 26324
rect 36360 26308 36412 26314
rect 36360 26250 36412 26256
rect 36176 25900 36228 25906
rect 36176 25842 36228 25848
rect 35900 25832 35952 25838
rect 35900 25774 35952 25780
rect 35912 23186 35940 25774
rect 36084 25696 36136 25702
rect 36084 25638 36136 25644
rect 36096 25362 36124 25638
rect 36084 25356 36136 25362
rect 36084 25298 36136 25304
rect 36188 24138 36216 25842
rect 36372 24818 36400 26250
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36556 26042 36584 26182
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 36556 25430 36584 25978
rect 37372 25968 37424 25974
rect 37372 25910 37424 25916
rect 36544 25424 36596 25430
rect 36544 25366 36596 25372
rect 36820 25356 36872 25362
rect 36820 25298 36872 25304
rect 36360 24812 36412 24818
rect 36360 24754 36412 24760
rect 36372 24410 36400 24754
rect 36360 24404 36412 24410
rect 36360 24346 36412 24352
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 36176 24132 36228 24138
rect 36176 24074 36228 24080
rect 35900 23180 35952 23186
rect 35900 23122 35952 23128
rect 36188 23118 36216 24074
rect 36268 23180 36320 23186
rect 36268 23122 36320 23128
rect 36176 23112 36228 23118
rect 36176 23054 36228 23060
rect 35808 22704 35860 22710
rect 35808 22646 35860 22652
rect 35820 22098 35848 22646
rect 35808 22092 35860 22098
rect 35808 22034 35860 22040
rect 36280 19378 36308 23122
rect 36556 22098 36584 24142
rect 36728 23792 36780 23798
rect 36728 23734 36780 23740
rect 36544 22092 36596 22098
rect 36544 22034 36596 22040
rect 36556 20466 36584 22034
rect 36636 20936 36688 20942
rect 36636 20878 36688 20884
rect 36544 20460 36596 20466
rect 36544 20402 36596 20408
rect 36360 19780 36412 19786
rect 36360 19722 36412 19728
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36176 19236 36228 19242
rect 36176 19178 36228 19184
rect 35728 17870 35848 17898
rect 35820 17678 35848 17870
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 35624 17672 35676 17678
rect 35808 17672 35860 17678
rect 35624 17614 35676 17620
rect 35806 17640 35808 17649
rect 35860 17640 35862 17649
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 35544 17134 35572 17614
rect 35532 17128 35584 17134
rect 35532 17070 35584 17076
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 34532 15706 34560 16050
rect 34520 15700 34572 15706
rect 34520 15642 34572 15648
rect 34520 14952 34572 14958
rect 34520 14894 34572 14900
rect 34532 14346 34560 14894
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 34532 10674 34560 14282
rect 34624 13462 34652 16526
rect 34796 16448 34848 16454
rect 34796 16390 34848 16396
rect 34704 15428 34756 15434
rect 34704 15370 34756 15376
rect 34612 13456 34664 13462
rect 34612 13398 34664 13404
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34532 10062 34560 10610
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34612 8832 34664 8838
rect 34612 8774 34664 8780
rect 34336 7744 34388 7750
rect 34336 7686 34388 7692
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34348 6322 34376 7346
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34532 6458 34560 6598
rect 34520 6452 34572 6458
rect 34520 6394 34572 6400
rect 34336 6316 34388 6322
rect 34336 6258 34388 6264
rect 34348 5642 34376 6258
rect 34336 5636 34388 5642
rect 34336 5578 34388 5584
rect 34520 4208 34572 4214
rect 34520 4150 34572 4156
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 33600 2372 33652 2378
rect 33600 2314 33652 2320
rect 34060 2372 34112 2378
rect 34060 2314 34112 2320
rect 33612 800 33640 2314
rect 34532 800 34560 4150
rect 34624 4010 34652 8774
rect 34716 4078 34744 15370
rect 34808 8838 34836 16390
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10130 35388 12718
rect 35544 12170 35572 17070
rect 35636 16998 35664 17614
rect 35806 17575 35862 17584
rect 36084 17536 36136 17542
rect 36084 17478 36136 17484
rect 35992 17264 36044 17270
rect 35992 17206 36044 17212
rect 35900 17196 35952 17202
rect 35900 17138 35952 17144
rect 35912 16998 35940 17138
rect 35624 16992 35676 16998
rect 35624 16934 35676 16940
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35636 14414 35664 16934
rect 35912 16794 35940 16934
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 36004 15434 36032 17206
rect 36096 17202 36124 17478
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36096 15910 36124 17138
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 35992 15428 36044 15434
rect 35992 15370 36044 15376
rect 35900 15360 35952 15366
rect 35900 15302 35952 15308
rect 35808 15020 35860 15026
rect 35912 15008 35940 15302
rect 35860 14980 35940 15008
rect 35808 14962 35860 14968
rect 35624 14408 35676 14414
rect 35624 14350 35676 14356
rect 35808 14272 35860 14278
rect 35808 14214 35860 14220
rect 35624 12844 35676 12850
rect 35624 12786 35676 12792
rect 35636 12442 35664 12786
rect 35624 12436 35676 12442
rect 35624 12378 35676 12384
rect 35532 12164 35584 12170
rect 35532 12106 35584 12112
rect 35544 11082 35572 12106
rect 35440 11076 35492 11082
rect 35440 11018 35492 11024
rect 35532 11076 35584 11082
rect 35532 11018 35584 11024
rect 35348 10124 35400 10130
rect 35348 10066 35400 10072
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 34808 7886 34836 8570
rect 35452 8498 35480 11018
rect 35544 10742 35572 11018
rect 35532 10736 35584 10742
rect 35532 10678 35584 10684
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35348 8288 35400 8294
rect 35348 8230 35400 8236
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 7954 35388 8230
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34808 5710 34836 7822
rect 35624 7744 35676 7750
rect 35624 7686 35676 7692
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35636 6798 35664 7686
rect 35728 6866 35756 8434
rect 35716 6860 35768 6866
rect 35716 6802 35768 6808
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35624 6792 35676 6798
rect 35820 6746 35848 14214
rect 35992 13728 36044 13734
rect 35992 13670 36044 13676
rect 36004 13326 36032 13670
rect 35992 13320 36044 13326
rect 35992 13262 36044 13268
rect 35900 13252 35952 13258
rect 35900 13194 35952 13200
rect 35912 12442 35940 13194
rect 35900 12436 35952 12442
rect 35900 12378 35952 12384
rect 35992 12368 36044 12374
rect 35992 12310 36044 12316
rect 36004 10742 36032 12310
rect 35992 10736 36044 10742
rect 35992 10678 36044 10684
rect 35992 10260 36044 10266
rect 35992 10202 36044 10208
rect 36004 8566 36032 10202
rect 36084 9512 36136 9518
rect 36084 9454 36136 9460
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 35992 8560 36044 8566
rect 35992 8502 36044 8508
rect 35912 8430 35940 8502
rect 35900 8424 35952 8430
rect 35900 8366 35952 8372
rect 35992 7880 36044 7886
rect 36096 7868 36124 9454
rect 36188 8430 36216 19178
rect 36372 18766 36400 19722
rect 36360 18760 36412 18766
rect 36648 18714 36676 20878
rect 36360 18702 36412 18708
rect 36556 18698 36676 18714
rect 36544 18692 36676 18698
rect 36596 18686 36676 18692
rect 36544 18634 36596 18640
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36360 17604 36412 17610
rect 36360 17546 36412 17552
rect 36372 17202 36400 17546
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36372 17082 36400 17138
rect 36280 17054 36400 17082
rect 36280 15978 36308 17054
rect 36360 16992 36412 16998
rect 36360 16934 36412 16940
rect 36268 15972 36320 15978
rect 36268 15914 36320 15920
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 36280 12238 36308 13126
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 36372 9602 36400 16934
rect 36464 14958 36492 18158
rect 36556 17746 36584 18634
rect 36544 17740 36596 17746
rect 36544 17682 36596 17688
rect 36556 17066 36584 17682
rect 36740 17218 36768 23734
rect 36832 23118 36860 25298
rect 37280 25152 37332 25158
rect 37280 25094 37332 25100
rect 37292 24206 37320 25094
rect 37280 24200 37332 24206
rect 37280 24142 37332 24148
rect 37384 23186 37412 25910
rect 37660 25838 37688 26318
rect 38752 26240 38804 26246
rect 38752 26182 38804 26188
rect 38764 25906 38792 26182
rect 38856 25974 38884 26386
rect 40040 26376 40092 26382
rect 39960 26324 40040 26330
rect 39960 26318 40092 26324
rect 40224 26376 40276 26382
rect 40224 26318 40276 26324
rect 39960 26302 40080 26318
rect 40132 26308 40184 26314
rect 38844 25968 38896 25974
rect 38844 25910 38896 25916
rect 38752 25900 38804 25906
rect 38752 25842 38804 25848
rect 39212 25900 39264 25906
rect 39212 25842 39264 25848
rect 37648 25832 37700 25838
rect 37648 25774 37700 25780
rect 37660 25294 37688 25774
rect 37648 25288 37700 25294
rect 37648 25230 37700 25236
rect 38752 25288 38804 25294
rect 38752 25230 38804 25236
rect 37660 24954 37688 25230
rect 37924 25152 37976 25158
rect 37924 25094 37976 25100
rect 37648 24948 37700 24954
rect 37648 24890 37700 24896
rect 37936 24818 37964 25094
rect 38384 24948 38436 24954
rect 38384 24890 38436 24896
rect 37924 24812 37976 24818
rect 37924 24754 37976 24760
rect 38396 24410 38424 24890
rect 38764 24818 38792 25230
rect 39224 24954 39252 25842
rect 39960 25498 39988 26302
rect 40132 26250 40184 26256
rect 40040 26240 40092 26246
rect 40040 26182 40092 26188
rect 40052 25906 40080 26182
rect 40144 26042 40172 26250
rect 40132 26036 40184 26042
rect 40132 25978 40184 25984
rect 40236 25974 40264 26318
rect 40224 25968 40276 25974
rect 40224 25910 40276 25916
rect 40328 25906 40356 26454
rect 40408 26376 40460 26382
rect 40408 26318 40460 26324
rect 40040 25900 40092 25906
rect 40040 25842 40092 25848
rect 40316 25900 40368 25906
rect 40316 25842 40368 25848
rect 39948 25492 40000 25498
rect 39948 25434 40000 25440
rect 39212 24948 39264 24954
rect 39212 24890 39264 24896
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 40052 24614 40080 25842
rect 40132 25696 40184 25702
rect 40132 25638 40184 25644
rect 39120 24608 39172 24614
rect 39120 24550 39172 24556
rect 40040 24608 40092 24614
rect 40040 24550 40092 24556
rect 38384 24404 38436 24410
rect 38384 24346 38436 24352
rect 39132 24206 39160 24550
rect 40144 24206 40172 25638
rect 40328 24818 40356 25842
rect 40420 25838 40448 26318
rect 40868 26308 40920 26314
rect 40868 26250 40920 26256
rect 40408 25832 40460 25838
rect 40408 25774 40460 25780
rect 40880 24818 40908 26250
rect 41052 25832 41104 25838
rect 41052 25774 41104 25780
rect 41064 25498 41092 25774
rect 41236 25696 41288 25702
rect 41236 25638 41288 25644
rect 41052 25492 41104 25498
rect 41052 25434 41104 25440
rect 40316 24812 40368 24818
rect 40316 24754 40368 24760
rect 40868 24812 40920 24818
rect 40868 24754 40920 24760
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40224 24200 40276 24206
rect 40224 24142 40276 24148
rect 38936 24064 38988 24070
rect 38936 24006 38988 24012
rect 39396 24064 39448 24070
rect 39396 24006 39448 24012
rect 38948 23882 38976 24006
rect 38856 23854 38976 23882
rect 37372 23180 37424 23186
rect 37372 23122 37424 23128
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36820 22976 36872 22982
rect 36820 22918 36872 22924
rect 36832 22098 36860 22918
rect 37384 22216 37412 23122
rect 38856 23050 38884 23854
rect 39408 23798 39436 24006
rect 39396 23792 39448 23798
rect 39396 23734 39448 23740
rect 40236 23662 40264 24142
rect 40328 23866 40356 24754
rect 40592 24744 40644 24750
rect 40592 24686 40644 24692
rect 40604 24206 40632 24686
rect 41248 24206 41276 25638
rect 40592 24200 40644 24206
rect 40592 24142 40644 24148
rect 41236 24200 41288 24206
rect 41236 24142 41288 24148
rect 40316 23860 40368 23866
rect 40316 23802 40368 23808
rect 40224 23656 40276 23662
rect 40224 23598 40276 23604
rect 40236 23118 40264 23598
rect 42168 23322 42196 39374
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 42616 25900 42668 25906
rect 42616 25842 42668 25848
rect 42628 24410 42656 25842
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 42616 24404 42668 24410
rect 42616 24346 42668 24352
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 42156 23316 42208 23322
rect 42156 23258 42208 23264
rect 40224 23112 40276 23118
rect 40224 23054 40276 23060
rect 38844 23044 38896 23050
rect 38844 22986 38896 22992
rect 37464 22228 37516 22234
rect 37384 22188 37464 22216
rect 36820 22092 36872 22098
rect 37384 22094 37412 22188
rect 37464 22170 37516 22176
rect 36820 22034 36872 22040
rect 37292 22066 37412 22094
rect 38856 22094 38884 22986
rect 38856 22066 38976 22094
rect 37096 20460 37148 20466
rect 37096 20402 37148 20408
rect 37108 19922 37136 20402
rect 37096 19916 37148 19922
rect 37096 19858 37148 19864
rect 37292 19378 37320 22066
rect 37556 21616 37608 21622
rect 37556 21558 37608 21564
rect 37372 21548 37424 21554
rect 37372 21490 37424 21496
rect 37384 19530 37412 21490
rect 37464 19984 37516 19990
rect 37464 19926 37516 19932
rect 37476 19854 37504 19926
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37384 19502 37504 19530
rect 37372 19440 37424 19446
rect 37372 19382 37424 19388
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37280 19236 37332 19242
rect 37280 19178 37332 19184
rect 37096 19168 37148 19174
rect 37096 19110 37148 19116
rect 36636 17196 36688 17202
rect 36740 17190 37044 17218
rect 36636 17138 36688 17144
rect 36648 17082 36676 17138
rect 36912 17128 36964 17134
rect 36544 17060 36596 17066
rect 36648 17054 36768 17082
rect 36912 17070 36964 17076
rect 36544 17002 36596 17008
rect 36740 16726 36768 17054
rect 36728 16720 36780 16726
rect 36728 16662 36780 16668
rect 36728 16516 36780 16522
rect 36728 16458 36780 16464
rect 36740 16114 36768 16458
rect 36728 16108 36780 16114
rect 36728 16050 36780 16056
rect 36740 15978 36768 16050
rect 36728 15972 36780 15978
rect 36728 15914 36780 15920
rect 36740 15638 36768 15914
rect 36820 15904 36872 15910
rect 36820 15846 36872 15852
rect 36832 15638 36860 15846
rect 36728 15632 36780 15638
rect 36728 15574 36780 15580
rect 36820 15632 36872 15638
rect 36820 15574 36872 15580
rect 36728 15496 36780 15502
rect 36726 15464 36728 15473
rect 36780 15464 36782 15473
rect 36636 15428 36688 15434
rect 36726 15399 36782 15408
rect 36636 15370 36688 15376
rect 36452 14952 36504 14958
rect 36452 14894 36504 14900
rect 36648 14618 36676 15370
rect 36740 15366 36768 15399
rect 36728 15360 36780 15366
rect 36728 15302 36780 15308
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 36728 14272 36780 14278
rect 36728 14214 36780 14220
rect 36740 13870 36768 14214
rect 36728 13864 36780 13870
rect 36728 13806 36780 13812
rect 36728 12640 36780 12646
rect 36728 12582 36780 12588
rect 36740 12238 36768 12582
rect 36728 12232 36780 12238
rect 36728 12174 36780 12180
rect 36728 11008 36780 11014
rect 36728 10950 36780 10956
rect 36740 10606 36768 10950
rect 36728 10600 36780 10606
rect 36728 10542 36780 10548
rect 36740 10266 36768 10542
rect 36728 10260 36780 10266
rect 36728 10202 36780 10208
rect 36280 9574 36400 9602
rect 36452 9648 36504 9654
rect 36452 9590 36504 9596
rect 36176 8424 36228 8430
rect 36176 8366 36228 8372
rect 36044 7840 36124 7868
rect 35992 7822 36044 7828
rect 35624 6734 35676 6740
rect 35544 6322 35572 6734
rect 35728 6718 35848 6746
rect 35624 6452 35676 6458
rect 35624 6394 35676 6400
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5704 34848 5710
rect 34796 5646 34848 5652
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34704 4072 34756 4078
rect 34704 4014 34756 4020
rect 34612 4004 34664 4010
rect 34612 3946 34664 3952
rect 34624 2446 34652 3946
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35544 3618 35572 6258
rect 35360 3590 35572 3618
rect 35360 3466 35388 3590
rect 35532 3528 35584 3534
rect 35532 3470 35584 3476
rect 35348 3460 35400 3466
rect 35348 3402 35400 3408
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34716 2394 34744 3334
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35544 2650 35572 3470
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 35636 2446 35664 6394
rect 35728 3194 35756 6718
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35820 5778 35848 6598
rect 36004 6254 36032 7822
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 35900 5704 35952 5710
rect 35900 5646 35952 5652
rect 35912 3602 35940 5646
rect 35992 5568 36044 5574
rect 35992 5510 36044 5516
rect 36004 5098 36032 5510
rect 35992 5092 36044 5098
rect 35992 5034 36044 5040
rect 36280 4554 36308 9574
rect 36464 8974 36492 9590
rect 36544 9444 36596 9450
rect 36544 9386 36596 9392
rect 36556 9178 36584 9386
rect 36544 9172 36596 9178
rect 36544 9114 36596 9120
rect 36636 9104 36688 9110
rect 36636 9046 36688 9052
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 36648 8498 36676 9046
rect 36636 8492 36688 8498
rect 36636 8434 36688 8440
rect 36728 8424 36780 8430
rect 36728 8366 36780 8372
rect 36740 6730 36768 8366
rect 36452 6724 36504 6730
rect 36452 6666 36504 6672
rect 36728 6724 36780 6730
rect 36728 6666 36780 6672
rect 36360 6248 36412 6254
rect 36360 6190 36412 6196
rect 36372 5710 36400 6190
rect 36360 5704 36412 5710
rect 36360 5646 36412 5652
rect 36464 5574 36492 6666
rect 36544 6656 36596 6662
rect 36544 6598 36596 6604
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 36556 5166 36584 6598
rect 36360 5160 36412 5166
rect 36360 5102 36412 5108
rect 36544 5160 36596 5166
rect 36544 5102 36596 5108
rect 36268 4548 36320 4554
rect 36268 4490 36320 4496
rect 36372 4078 36400 5102
rect 36556 4826 36584 5102
rect 36544 4820 36596 4826
rect 36544 4762 36596 4768
rect 36360 4072 36412 4078
rect 36360 4014 36412 4020
rect 36372 3890 36400 4014
rect 36372 3862 36492 3890
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 35716 3188 35768 3194
rect 35716 3130 35768 3136
rect 35900 3120 35952 3126
rect 35900 3062 35952 3068
rect 34980 2440 35032 2446
rect 34716 2388 34980 2394
rect 34716 2382 35032 2388
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 34716 2366 35020 2382
rect 35268 1902 35296 2382
rect 35256 1896 35308 1902
rect 35256 1838 35308 1844
rect 34980 944 35032 950
rect 34980 886 35032 892
rect 34992 800 35020 886
rect 35912 800 35940 3062
rect 36464 3058 36492 3862
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36360 2984 36412 2990
rect 36360 2926 36412 2932
rect 36268 2372 36320 2378
rect 36268 2314 36320 2320
rect 36280 950 36308 2314
rect 36268 944 36320 950
rect 36268 886 36320 892
rect 36372 800 36400 2926
rect 36924 2650 36952 17070
rect 37016 14618 37044 17190
rect 37004 14612 37056 14618
rect 37004 14554 37056 14560
rect 37016 14414 37044 14554
rect 37004 14408 37056 14414
rect 37004 14350 37056 14356
rect 37108 13326 37136 19110
rect 37292 18358 37320 19178
rect 37280 18352 37332 18358
rect 37280 18294 37332 18300
rect 37292 18170 37320 18294
rect 37200 18142 37320 18170
rect 37200 17542 37228 18142
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37292 17678 37320 18022
rect 37280 17672 37332 17678
rect 37280 17614 37332 17620
rect 37384 17610 37412 19382
rect 37476 19174 37504 19502
rect 37464 19168 37516 19174
rect 37464 19110 37516 19116
rect 37476 18766 37504 19110
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37372 17604 37424 17610
rect 37372 17546 37424 17552
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 37280 17536 37332 17542
rect 37280 17478 37332 17484
rect 37292 17270 37320 17478
rect 37476 17338 37504 18226
rect 37464 17332 37516 17338
rect 37464 17274 37516 17280
rect 37280 17264 37332 17270
rect 37280 17206 37332 17212
rect 37188 17060 37240 17066
rect 37188 17002 37240 17008
rect 37200 15026 37228 17002
rect 37292 16658 37320 17206
rect 37568 17202 37596 21558
rect 38660 20868 38712 20874
rect 38660 20810 38712 20816
rect 38016 20800 38068 20806
rect 38016 20742 38068 20748
rect 38028 20602 38056 20742
rect 37648 20596 37700 20602
rect 37648 20538 37700 20544
rect 38016 20596 38068 20602
rect 38016 20538 38068 20544
rect 37660 19378 37688 20538
rect 37740 20460 37792 20466
rect 37740 20402 37792 20408
rect 37752 20058 37780 20402
rect 38108 20256 38160 20262
rect 38108 20198 38160 20204
rect 37740 20052 37792 20058
rect 37740 19994 37792 20000
rect 38016 19848 38068 19854
rect 38016 19790 38068 19796
rect 38028 19689 38056 19790
rect 38014 19680 38070 19689
rect 38014 19615 38070 19624
rect 38120 19378 38148 20198
rect 38672 19922 38700 20810
rect 38844 20256 38896 20262
rect 38844 20198 38896 20204
rect 38856 19990 38884 20198
rect 38844 19984 38896 19990
rect 38844 19926 38896 19932
rect 38660 19916 38712 19922
rect 38660 19858 38712 19864
rect 38568 19712 38620 19718
rect 38566 19680 38568 19689
rect 38620 19680 38622 19689
rect 38566 19615 38622 19624
rect 38476 19440 38528 19446
rect 38476 19382 38528 19388
rect 37648 19372 37700 19378
rect 37648 19314 37700 19320
rect 38016 19372 38068 19378
rect 38016 19314 38068 19320
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 37648 18760 37700 18766
rect 37648 18702 37700 18708
rect 37660 18290 37688 18702
rect 37648 18284 37700 18290
rect 37648 18226 37700 18232
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 37738 17640 37794 17649
rect 37738 17575 37794 17584
rect 37556 17196 37608 17202
rect 37556 17138 37608 17144
rect 37280 16652 37332 16658
rect 37280 16594 37332 16600
rect 37280 16448 37332 16454
rect 37280 16390 37332 16396
rect 37464 16448 37516 16454
rect 37464 16390 37516 16396
rect 37292 16250 37320 16390
rect 37280 16244 37332 16250
rect 37280 16186 37332 16192
rect 37292 15638 37320 16186
rect 37476 16182 37504 16390
rect 37464 16176 37516 16182
rect 37464 16118 37516 16124
rect 37280 15632 37332 15638
rect 37280 15574 37332 15580
rect 37568 15366 37596 17138
rect 37648 16516 37700 16522
rect 37648 16458 37700 16464
rect 37660 16182 37688 16458
rect 37648 16176 37700 16182
rect 37648 16118 37700 16124
rect 37556 15360 37608 15366
rect 37556 15302 37608 15308
rect 37188 15020 37240 15026
rect 37188 14962 37240 14968
rect 37752 14006 37780 17575
rect 37936 17202 37964 17818
rect 38028 17814 38056 19314
rect 38108 18148 38160 18154
rect 38108 18090 38160 18096
rect 38016 17808 38068 17814
rect 38016 17750 38068 17756
rect 38028 17270 38056 17750
rect 38016 17264 38068 17270
rect 38016 17206 38068 17212
rect 37924 17196 37976 17202
rect 37924 17138 37976 17144
rect 37832 17060 37884 17066
rect 37832 17002 37884 17008
rect 37844 16794 37872 17002
rect 37832 16788 37884 16794
rect 37832 16730 37884 16736
rect 38120 16046 38148 18090
rect 38108 16040 38160 16046
rect 38108 15982 38160 15988
rect 38120 15586 38148 15982
rect 38028 15558 38148 15586
rect 37740 14000 37792 14006
rect 37740 13942 37792 13948
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37648 13932 37700 13938
rect 37648 13874 37700 13880
rect 37476 13462 37504 13874
rect 37464 13456 37516 13462
rect 37464 13398 37516 13404
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 37108 10470 37136 13262
rect 37292 12986 37320 13330
rect 37556 13252 37608 13258
rect 37556 13194 37608 13200
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37292 12782 37320 12922
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 37292 12434 37320 12718
rect 37200 12406 37320 12434
rect 37200 12306 37228 12406
rect 37188 12300 37240 12306
rect 37188 12242 37240 12248
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 37096 10464 37148 10470
rect 37096 10406 37148 10412
rect 37476 10062 37504 10950
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37200 9654 37228 9998
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 37200 9042 37228 9590
rect 37188 9036 37240 9042
rect 37188 8978 37240 8984
rect 37568 8974 37596 13194
rect 37660 12986 37688 13874
rect 37648 12980 37700 12986
rect 37648 12922 37700 12928
rect 37924 11552 37976 11558
rect 37924 11494 37976 11500
rect 37648 11144 37700 11150
rect 37648 11086 37700 11092
rect 37660 10810 37688 11086
rect 37936 11082 37964 11494
rect 38028 11218 38056 15558
rect 38108 14068 38160 14074
rect 38108 14010 38160 14016
rect 38120 12986 38148 14010
rect 38108 12980 38160 12986
rect 38108 12922 38160 12928
rect 38120 12374 38148 12922
rect 38292 12776 38344 12782
rect 38292 12718 38344 12724
rect 38304 12434 38332 12718
rect 38304 12406 38424 12434
rect 38108 12368 38160 12374
rect 38108 12310 38160 12316
rect 38016 11212 38068 11218
rect 38016 11154 38068 11160
rect 37924 11076 37976 11082
rect 37924 11018 37976 11024
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 37648 10804 37700 10810
rect 37648 10746 37700 10752
rect 38016 10668 38068 10674
rect 38016 10610 38068 10616
rect 38028 9926 38056 10610
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37556 8832 37608 8838
rect 37556 8774 37608 8780
rect 37568 8430 37596 8774
rect 37740 8560 37792 8566
rect 37740 8502 37792 8508
rect 37556 8424 37608 8430
rect 37608 8384 37688 8412
rect 37556 8366 37608 8372
rect 37660 6322 37688 8384
rect 37752 7546 37780 8502
rect 38016 8424 38068 8430
rect 38016 8366 38068 8372
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37844 7886 37872 8230
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37740 7540 37792 7546
rect 37740 7482 37792 7488
rect 38028 6322 38056 8366
rect 37648 6316 37700 6322
rect 37648 6258 37700 6264
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 38016 6316 38068 6322
rect 38016 6258 38068 6264
rect 37660 4758 37688 6258
rect 37844 5914 37872 6258
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 37832 5364 37884 5370
rect 37832 5306 37884 5312
rect 37648 4752 37700 4758
rect 37648 4694 37700 4700
rect 37280 3392 37332 3398
rect 37280 3334 37332 3340
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37292 2514 37320 3334
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37844 2446 37872 5306
rect 38016 4752 38068 4758
rect 38016 4694 38068 4700
rect 38028 4622 38056 4694
rect 38120 4622 38148 11018
rect 38396 10606 38424 12406
rect 38488 11082 38516 19382
rect 38660 18080 38712 18086
rect 38660 18022 38712 18028
rect 38672 17134 38700 18022
rect 38660 17128 38712 17134
rect 38660 17070 38712 17076
rect 38672 16658 38700 17070
rect 38660 16652 38712 16658
rect 38660 16594 38712 16600
rect 38844 16448 38896 16454
rect 38844 16390 38896 16396
rect 38856 15162 38884 16390
rect 38844 15156 38896 15162
rect 38844 15098 38896 15104
rect 38844 14408 38896 14414
rect 38844 14350 38896 14356
rect 38856 12322 38884 14350
rect 38948 13870 38976 22066
rect 40236 22030 40264 23054
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 40224 22024 40276 22030
rect 40224 21966 40276 21972
rect 40236 21010 40264 21966
rect 40592 21956 40644 21962
rect 40592 21898 40644 21904
rect 40604 21690 40632 21898
rect 40960 21888 41012 21894
rect 40960 21830 41012 21836
rect 40972 21690 41000 21830
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 40592 21684 40644 21690
rect 40592 21626 40644 21632
rect 40960 21684 41012 21690
rect 40960 21626 41012 21632
rect 40408 21480 40460 21486
rect 40408 21422 40460 21428
rect 40224 21004 40276 21010
rect 40224 20946 40276 20952
rect 40236 20534 40264 20946
rect 40224 20528 40276 20534
rect 40224 20470 40276 20476
rect 40420 19854 40448 21422
rect 40972 21146 41000 21626
rect 45192 21548 45244 21554
rect 45192 21490 45244 21496
rect 41236 21344 41288 21350
rect 41236 21286 41288 21292
rect 40960 21140 41012 21146
rect 40960 21082 41012 21088
rect 41248 20942 41276 21286
rect 45204 21146 45232 21490
rect 45836 21480 45888 21486
rect 45836 21422 45888 21428
rect 45192 21140 45244 21146
rect 45192 21082 45244 21088
rect 43444 21072 43496 21078
rect 43444 21014 43496 21020
rect 41236 20936 41288 20942
rect 41236 20878 41288 20884
rect 41420 20460 41472 20466
rect 41420 20402 41472 20408
rect 41432 20058 41460 20402
rect 42064 20256 42116 20262
rect 42064 20198 42116 20204
rect 41420 20052 41472 20058
rect 41420 19994 41472 20000
rect 42076 19854 42104 20198
rect 40408 19848 40460 19854
rect 40408 19790 40460 19796
rect 41604 19848 41656 19854
rect 41604 19790 41656 19796
rect 42064 19848 42116 19854
rect 42064 19790 42116 19796
rect 40316 18692 40368 18698
rect 40316 18634 40368 18640
rect 40224 18284 40276 18290
rect 40224 18226 40276 18232
rect 40040 18148 40092 18154
rect 40040 18090 40092 18096
rect 40052 17678 40080 18090
rect 40040 17672 40092 17678
rect 40040 17614 40092 17620
rect 40236 17542 40264 18226
rect 40224 17536 40276 17542
rect 40224 17478 40276 17484
rect 40236 17270 40264 17478
rect 40224 17264 40276 17270
rect 40224 17206 40276 17212
rect 40328 16658 40356 18634
rect 40316 16652 40368 16658
rect 40316 16594 40368 16600
rect 40040 16516 40092 16522
rect 40040 16458 40092 16464
rect 40052 16250 40080 16458
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 40224 16108 40276 16114
rect 40224 16050 40276 16056
rect 40236 15706 40264 16050
rect 40224 15700 40276 15706
rect 40224 15642 40276 15648
rect 40328 15570 40356 16594
rect 40420 16250 40448 19790
rect 41616 19378 41644 19790
rect 41604 19372 41656 19378
rect 41604 19314 41656 19320
rect 40960 19168 41012 19174
rect 40960 19110 41012 19116
rect 40972 18766 41000 19110
rect 41328 18828 41380 18834
rect 41328 18770 41380 18776
rect 40960 18760 41012 18766
rect 40960 18702 41012 18708
rect 40592 18624 40644 18630
rect 40592 18566 40644 18572
rect 40604 18426 40632 18566
rect 40500 18420 40552 18426
rect 40500 18362 40552 18368
rect 40592 18420 40644 18426
rect 40592 18362 40644 18368
rect 40512 17882 40540 18362
rect 41236 18352 41288 18358
rect 41236 18294 41288 18300
rect 40592 18284 40644 18290
rect 40592 18226 40644 18232
rect 40500 17876 40552 17882
rect 40500 17818 40552 17824
rect 40604 17814 40632 18226
rect 40592 17808 40644 17814
rect 40592 17750 40644 17756
rect 40604 17678 40632 17750
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40500 17536 40552 17542
rect 40500 17478 40552 17484
rect 40408 16244 40460 16250
rect 40408 16186 40460 16192
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 40316 14612 40368 14618
rect 40316 14554 40368 14560
rect 40224 14544 40276 14550
rect 40052 14492 40224 14498
rect 40052 14486 40276 14492
rect 40052 14470 40264 14486
rect 40052 14346 40080 14470
rect 40040 14340 40092 14346
rect 40040 14282 40092 14288
rect 40132 14340 40184 14346
rect 40132 14282 40184 14288
rect 38936 13864 38988 13870
rect 38988 13812 39252 13818
rect 38936 13806 39252 13812
rect 38948 13790 39252 13806
rect 38752 12300 38804 12306
rect 38752 12242 38804 12248
rect 38856 12294 39068 12322
rect 38660 12232 38712 12238
rect 38660 12174 38712 12180
rect 38568 11756 38620 11762
rect 38568 11698 38620 11704
rect 38580 11354 38608 11698
rect 38672 11558 38700 12174
rect 38660 11552 38712 11558
rect 38660 11494 38712 11500
rect 38568 11348 38620 11354
rect 38568 11290 38620 11296
rect 38764 11150 38792 12242
rect 38856 11762 38884 12294
rect 39040 12238 39068 12294
rect 39224 12238 39252 13790
rect 39856 13184 39908 13190
rect 39856 13126 39908 13132
rect 39868 12850 39896 13126
rect 40052 12986 40080 14282
rect 40040 12980 40092 12986
rect 40040 12922 40092 12928
rect 39856 12844 39908 12850
rect 39856 12786 39908 12792
rect 40040 12844 40092 12850
rect 40040 12786 40092 12792
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 39212 12232 39264 12238
rect 39212 12174 39264 12180
rect 38936 12164 38988 12170
rect 38936 12106 38988 12112
rect 38844 11756 38896 11762
rect 38844 11698 38896 11704
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38476 11076 38528 11082
rect 38476 11018 38528 11024
rect 38384 10600 38436 10606
rect 38384 10542 38436 10548
rect 38396 10130 38424 10542
rect 38384 10124 38436 10130
rect 38384 10066 38436 10072
rect 38396 7342 38424 10066
rect 38856 10062 38884 11698
rect 38948 11286 38976 12106
rect 39868 11830 39896 12786
rect 39028 11824 39080 11830
rect 39028 11766 39080 11772
rect 39856 11824 39908 11830
rect 39856 11766 39908 11772
rect 38936 11280 38988 11286
rect 38936 11222 38988 11228
rect 39040 11082 39068 11766
rect 39948 11756 40000 11762
rect 39948 11698 40000 11704
rect 39120 11688 39172 11694
rect 39120 11630 39172 11636
rect 39132 11150 39160 11630
rect 39960 11150 39988 11698
rect 40052 11626 40080 12786
rect 40144 11898 40172 14282
rect 40328 14278 40356 14554
rect 40316 14272 40368 14278
rect 40316 14214 40368 14220
rect 40224 12096 40276 12102
rect 40224 12038 40276 12044
rect 40408 12096 40460 12102
rect 40408 12038 40460 12044
rect 40132 11892 40184 11898
rect 40132 11834 40184 11840
rect 40040 11620 40092 11626
rect 40040 11562 40092 11568
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 39304 11144 39356 11150
rect 39304 11086 39356 11092
rect 39948 11144 40000 11150
rect 39948 11086 40000 11092
rect 38936 11076 38988 11082
rect 38936 11018 38988 11024
rect 39028 11076 39080 11082
rect 39028 11018 39080 11024
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 38660 9580 38712 9586
rect 38660 9522 38712 9528
rect 38672 7750 38700 9522
rect 38856 9110 38884 9998
rect 38844 9104 38896 9110
rect 38844 9046 38896 9052
rect 38856 8498 38884 9046
rect 38844 8492 38896 8498
rect 38844 8434 38896 8440
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 38672 7410 38700 7686
rect 38660 7404 38712 7410
rect 38660 7346 38712 7352
rect 38200 7336 38252 7342
rect 38200 7278 38252 7284
rect 38384 7336 38436 7342
rect 38384 7278 38436 7284
rect 38212 5370 38240 7278
rect 38396 6662 38424 7278
rect 38384 6656 38436 6662
rect 38384 6598 38436 6604
rect 38200 5364 38252 5370
rect 38200 5306 38252 5312
rect 38384 5364 38436 5370
rect 38384 5306 38436 5312
rect 38292 5024 38344 5030
rect 38292 4966 38344 4972
rect 38304 4622 38332 4966
rect 38396 4758 38424 5306
rect 38752 5024 38804 5030
rect 38752 4966 38804 4972
rect 38384 4752 38436 4758
rect 38384 4694 38436 4700
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38108 4616 38160 4622
rect 38108 4558 38160 4564
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38292 4480 38344 4486
rect 38292 4422 38344 4428
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 38212 3058 38240 3470
rect 38304 3058 38332 4422
rect 38660 4208 38712 4214
rect 38660 4150 38712 4156
rect 38200 3052 38252 3058
rect 38200 2994 38252 3000
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 37832 2440 37884 2446
rect 37832 2382 37884 2388
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37280 944 37332 950
rect 37280 886 37332 892
rect 37292 800 37320 886
rect 37752 800 37780 2314
rect 38672 800 38700 4150
rect 38764 3534 38792 4966
rect 38948 4146 38976 11018
rect 39040 10146 39068 11018
rect 39040 10118 39160 10146
rect 39028 9988 39080 9994
rect 39028 9930 39080 9936
rect 39040 9722 39068 9930
rect 39028 9716 39080 9722
rect 39028 9658 39080 9664
rect 39028 9580 39080 9586
rect 39132 9568 39160 10118
rect 39210 10024 39266 10033
rect 39210 9959 39212 9968
rect 39264 9959 39266 9968
rect 39212 9930 39264 9936
rect 39080 9540 39160 9568
rect 39212 9580 39264 9586
rect 39028 9522 39080 9528
rect 39316 9568 39344 11086
rect 40236 10266 40264 12038
rect 40420 10742 40448 12038
rect 40408 10736 40460 10742
rect 40408 10678 40460 10684
rect 40224 10260 40276 10266
rect 40224 10202 40276 10208
rect 39856 10192 39908 10198
rect 39856 10134 39908 10140
rect 39264 9540 39344 9568
rect 39486 9616 39542 9625
rect 39868 9586 39896 10134
rect 39486 9551 39542 9560
rect 39856 9580 39908 9586
rect 39212 9522 39264 9528
rect 39040 7274 39068 9522
rect 39224 8906 39252 9522
rect 39212 8900 39264 8906
rect 39212 8842 39264 8848
rect 39500 8634 39528 9551
rect 39856 9522 39908 9528
rect 40132 8968 40184 8974
rect 40132 8910 40184 8916
rect 39488 8628 39540 8634
rect 39488 8570 39540 8576
rect 40144 8430 40172 8910
rect 40316 8900 40368 8906
rect 40316 8842 40368 8848
rect 40040 8424 40092 8430
rect 40040 8366 40092 8372
rect 40132 8424 40184 8430
rect 40132 8366 40184 8372
rect 40052 7970 40080 8366
rect 40052 7942 40172 7970
rect 40328 7954 40356 8842
rect 40408 8560 40460 8566
rect 40408 8502 40460 8508
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 39212 7404 39264 7410
rect 39212 7346 39264 7352
rect 39028 7268 39080 7274
rect 39028 7210 39080 7216
rect 39120 4480 39172 4486
rect 39120 4422 39172 4428
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 39132 4078 39160 4422
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 38752 3528 38804 3534
rect 38752 3470 38804 3476
rect 39132 3194 39160 4014
rect 39120 3188 39172 3194
rect 39120 3130 39172 3136
rect 39224 2446 39252 7346
rect 40052 6118 40080 7822
rect 40144 7818 40172 7942
rect 40316 7948 40368 7954
rect 40316 7890 40368 7896
rect 40132 7812 40184 7818
rect 40132 7754 40184 7760
rect 40224 7812 40276 7818
rect 40224 7754 40276 7760
rect 40144 6322 40172 7754
rect 40236 7274 40264 7754
rect 40328 7426 40356 7890
rect 40420 7750 40448 8502
rect 40408 7744 40460 7750
rect 40408 7686 40460 7692
rect 40328 7398 40448 7426
rect 40224 7268 40276 7274
rect 40224 7210 40276 7216
rect 40132 6316 40184 6322
rect 40132 6258 40184 6264
rect 40040 6112 40092 6118
rect 40040 6054 40092 6060
rect 40236 5710 40264 7210
rect 40316 6112 40368 6118
rect 40316 6054 40368 6060
rect 40040 5704 40092 5710
rect 40040 5646 40092 5652
rect 40224 5704 40276 5710
rect 40224 5646 40276 5652
rect 40052 5098 40080 5646
rect 40328 5642 40356 6054
rect 40420 5710 40448 7398
rect 40408 5704 40460 5710
rect 40408 5646 40460 5652
rect 40316 5636 40368 5642
rect 40316 5578 40368 5584
rect 40040 5092 40092 5098
rect 40040 5034 40092 5040
rect 40052 3738 40080 5034
rect 40224 4480 40276 4486
rect 40224 4422 40276 4428
rect 40040 3732 40092 3738
rect 40040 3674 40092 3680
rect 40040 3460 40092 3466
rect 40040 3402 40092 3408
rect 39212 2440 39264 2446
rect 39212 2382 39264 2388
rect 38844 2372 38896 2378
rect 38844 2314 38896 2320
rect 38856 950 38884 2314
rect 38844 944 38896 950
rect 38844 886 38896 892
rect 39120 944 39172 950
rect 39120 886 39172 892
rect 39132 800 39160 886
rect 40052 800 40080 3402
rect 40236 2854 40264 4422
rect 40224 2848 40276 2854
rect 40224 2790 40276 2796
rect 40328 2650 40356 5578
rect 40512 3670 40540 17478
rect 40776 14000 40828 14006
rect 40776 13942 40828 13948
rect 40788 13326 40816 13942
rect 40776 13320 40828 13326
rect 40776 13262 40828 13268
rect 40776 12980 40828 12986
rect 40776 12922 40828 12928
rect 40788 12850 40816 12922
rect 40776 12844 40828 12850
rect 40776 12786 40828 12792
rect 40684 11144 40736 11150
rect 40684 11086 40736 11092
rect 40696 10606 40724 11086
rect 40684 10600 40736 10606
rect 40684 10542 40736 10548
rect 40696 9518 40724 10542
rect 40788 9586 40816 12786
rect 40776 9580 40828 9586
rect 40776 9522 40828 9528
rect 40684 9512 40736 9518
rect 40684 9454 40736 9460
rect 40788 8566 40816 9522
rect 40960 9376 41012 9382
rect 40960 9318 41012 9324
rect 40776 8560 40828 8566
rect 40776 8502 40828 8508
rect 40868 8492 40920 8498
rect 40868 8434 40920 8440
rect 40684 8356 40736 8362
rect 40880 8344 40908 8434
rect 40736 8316 40908 8344
rect 40684 8298 40736 8304
rect 40592 8288 40644 8294
rect 40592 8230 40644 8236
rect 40604 8090 40632 8230
rect 40592 8084 40644 8090
rect 40592 8026 40644 8032
rect 40500 3664 40552 3670
rect 40500 3606 40552 3612
rect 40316 2644 40368 2650
rect 40316 2586 40368 2592
rect 40972 2446 41000 9318
rect 41052 7880 41104 7886
rect 41052 7822 41104 7828
rect 41064 6798 41092 7822
rect 41052 6792 41104 6798
rect 41052 6734 41104 6740
rect 41064 5778 41092 6734
rect 41052 5772 41104 5778
rect 41052 5714 41104 5720
rect 41064 3534 41092 5714
rect 41144 5568 41196 5574
rect 41144 5510 41196 5516
rect 41156 5302 41184 5510
rect 41144 5296 41196 5302
rect 41144 5238 41196 5244
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 41064 3126 41092 3470
rect 41248 3194 41276 18294
rect 41340 18290 41368 18770
rect 41604 18624 41656 18630
rect 41604 18566 41656 18572
rect 41328 18284 41380 18290
rect 41328 18226 41380 18232
rect 41512 18284 41564 18290
rect 41512 18226 41564 18232
rect 41524 18086 41552 18226
rect 41616 18086 41644 18566
rect 42076 18222 42104 19790
rect 42892 19780 42944 19786
rect 42892 19722 42944 19728
rect 42432 19440 42484 19446
rect 42432 19382 42484 19388
rect 42444 18902 42472 19382
rect 42904 19310 42932 19722
rect 43352 19712 43404 19718
rect 43352 19654 43404 19660
rect 42982 19408 43038 19417
rect 43364 19378 43392 19654
rect 42982 19343 43038 19352
rect 43352 19372 43404 19378
rect 42892 19304 42944 19310
rect 42892 19246 42944 19252
rect 42800 19168 42852 19174
rect 42800 19110 42852 19116
rect 42812 18902 42840 19110
rect 42432 18896 42484 18902
rect 42432 18838 42484 18844
rect 42800 18896 42852 18902
rect 42800 18838 42852 18844
rect 42340 18760 42392 18766
rect 42340 18702 42392 18708
rect 42156 18692 42208 18698
rect 42156 18634 42208 18640
rect 42168 18426 42196 18634
rect 42156 18420 42208 18426
rect 42156 18362 42208 18368
rect 42064 18216 42116 18222
rect 42064 18158 42116 18164
rect 41512 18080 41564 18086
rect 41512 18022 41564 18028
rect 41604 18080 41656 18086
rect 41604 18022 41656 18028
rect 41616 17746 41644 18022
rect 41604 17740 41656 17746
rect 41604 17682 41656 17688
rect 41604 14272 41656 14278
rect 41604 14214 41656 14220
rect 41616 13326 41644 14214
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 41604 13320 41656 13326
rect 41604 13262 41656 13268
rect 41340 12238 41368 13262
rect 41420 12640 41472 12646
rect 41420 12582 41472 12588
rect 41432 12238 41460 12582
rect 42352 12434 42380 18702
rect 42996 15910 43024 19343
rect 43352 19314 43404 19320
rect 43456 18714 43484 21014
rect 45848 20942 45876 21422
rect 45836 20936 45888 20942
rect 45836 20878 45888 20884
rect 44456 20596 44508 20602
rect 44456 20538 44508 20544
rect 44468 19854 44496 20538
rect 45848 19854 45876 20878
rect 45928 20868 45980 20874
rect 45928 20810 45980 20816
rect 44180 19848 44232 19854
rect 44180 19790 44232 19796
rect 44456 19848 44508 19854
rect 44456 19790 44508 19796
rect 45560 19848 45612 19854
rect 45560 19790 45612 19796
rect 45652 19848 45704 19854
rect 45652 19790 45704 19796
rect 45836 19848 45888 19854
rect 45836 19790 45888 19796
rect 44192 19378 44220 19790
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 44180 19372 44232 19378
rect 44180 19314 44232 19320
rect 43916 19174 43944 19314
rect 43904 19168 43956 19174
rect 43904 19110 43956 19116
rect 43916 18902 43944 19110
rect 43904 18896 43956 18902
rect 43904 18838 43956 18844
rect 44192 18834 44220 19314
rect 44468 19310 44496 19790
rect 45572 19446 45600 19790
rect 45664 19514 45692 19790
rect 45652 19508 45704 19514
rect 45652 19450 45704 19456
rect 45560 19440 45612 19446
rect 45560 19382 45612 19388
rect 44456 19304 44508 19310
rect 44456 19246 44508 19252
rect 44468 18970 44496 19246
rect 44456 18964 44508 18970
rect 44456 18906 44508 18912
rect 44180 18828 44232 18834
rect 44180 18770 44232 18776
rect 43456 18686 43852 18714
rect 43076 18352 43128 18358
rect 43076 18294 43128 18300
rect 42984 15904 43036 15910
rect 42984 15846 43036 15852
rect 42616 15428 42668 15434
rect 42616 15370 42668 15376
rect 42628 15162 42656 15370
rect 42996 15162 43024 15846
rect 42616 15156 42668 15162
rect 42616 15098 42668 15104
rect 42984 15156 43036 15162
rect 42984 15098 43036 15104
rect 42260 12406 42380 12434
rect 41328 12232 41380 12238
rect 41328 12174 41380 12180
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 41340 11150 41368 12174
rect 41328 11144 41380 11150
rect 41328 11086 41380 11092
rect 42260 9178 42288 12406
rect 42340 12164 42392 12170
rect 42340 12106 42392 12112
rect 42352 10742 42380 12106
rect 42432 12096 42484 12102
rect 42432 12038 42484 12044
rect 42444 11694 42472 12038
rect 42432 11688 42484 11694
rect 42432 11630 42484 11636
rect 42340 10736 42392 10742
rect 42340 10678 42392 10684
rect 42248 9172 42300 9178
rect 42248 9114 42300 9120
rect 41512 8424 41564 8430
rect 41512 8366 41564 8372
rect 41524 7886 41552 8366
rect 41512 7880 41564 7886
rect 41512 7822 41564 7828
rect 41696 7336 41748 7342
rect 41696 7278 41748 7284
rect 41708 5370 41736 7278
rect 42156 6724 42208 6730
rect 42156 6666 42208 6672
rect 42168 6390 42196 6666
rect 42156 6384 42208 6390
rect 42156 6326 42208 6332
rect 42340 5568 42392 5574
rect 42340 5510 42392 5516
rect 41696 5364 41748 5370
rect 41696 5306 41748 5312
rect 41420 5228 41472 5234
rect 41420 5170 41472 5176
rect 41432 4826 41460 5170
rect 41708 5114 41736 5306
rect 42352 5302 42380 5510
rect 42340 5296 42392 5302
rect 41786 5264 41842 5273
rect 42340 5238 42392 5244
rect 41786 5199 41788 5208
rect 41840 5199 41842 5208
rect 41788 5170 41840 5176
rect 41708 5086 41828 5114
rect 41420 4820 41472 4826
rect 41420 4762 41472 4768
rect 41696 4820 41748 4826
rect 41696 4762 41748 4768
rect 41708 4622 41736 4762
rect 41800 4622 41828 5086
rect 41696 4616 41748 4622
rect 41696 4558 41748 4564
rect 41788 4616 41840 4622
rect 41788 4558 41840 4564
rect 42064 4616 42116 4622
rect 42064 4558 42116 4564
rect 41420 4480 41472 4486
rect 41420 4422 41472 4428
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 41052 3120 41104 3126
rect 41052 3062 41104 3068
rect 41432 3058 41460 4422
rect 41800 4214 41828 4558
rect 42076 4282 42104 4558
rect 42064 4276 42116 4282
rect 42064 4218 42116 4224
rect 41788 4208 41840 4214
rect 41788 4150 41840 4156
rect 41512 3120 41564 3126
rect 41512 3062 41564 3068
rect 41420 3052 41472 3058
rect 41420 2994 41472 3000
rect 40960 2440 41012 2446
rect 40960 2382 41012 2388
rect 40316 2372 40368 2378
rect 40316 2314 40368 2320
rect 40500 2372 40552 2378
rect 40500 2314 40552 2320
rect 40328 950 40356 2314
rect 40316 944 40368 950
rect 40316 886 40368 892
rect 40512 800 40540 2314
rect 41524 1578 41552 3062
rect 42444 2514 42472 11630
rect 42984 11076 43036 11082
rect 42984 11018 43036 11024
rect 42996 10810 43024 11018
rect 42984 10804 43036 10810
rect 42984 10746 43036 10752
rect 42524 10464 42576 10470
rect 42524 10406 42576 10412
rect 42536 9926 42564 10406
rect 42524 9920 42576 9926
rect 42524 9862 42576 9868
rect 42432 2508 42484 2514
rect 42432 2450 42484 2456
rect 42536 2446 42564 9862
rect 43088 7698 43116 18294
rect 43456 18290 43484 18686
rect 43824 18630 43852 18686
rect 44180 18692 44232 18698
rect 44180 18634 44232 18640
rect 44272 18692 44324 18698
rect 44272 18634 44324 18640
rect 43720 18624 43772 18630
rect 43720 18566 43772 18572
rect 43812 18624 43864 18630
rect 43812 18566 43864 18572
rect 43732 18290 43760 18566
rect 43260 18284 43312 18290
rect 43260 18226 43312 18232
rect 43444 18284 43496 18290
rect 43444 18226 43496 18232
rect 43536 18284 43588 18290
rect 43536 18226 43588 18232
rect 43720 18284 43772 18290
rect 43720 18226 43772 18232
rect 43272 18154 43300 18226
rect 43260 18148 43312 18154
rect 43260 18090 43312 18096
rect 43548 17338 43576 18226
rect 44192 18154 44220 18634
rect 44284 18222 44312 18634
rect 44468 18426 44496 18906
rect 45572 18698 45600 19382
rect 45940 19242 45968 20810
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 45928 19236 45980 19242
rect 45928 19178 45980 19184
rect 45940 18834 45968 19178
rect 45928 18828 45980 18834
rect 45928 18770 45980 18776
rect 45560 18692 45612 18698
rect 45560 18634 45612 18640
rect 44456 18420 44508 18426
rect 44456 18362 44508 18368
rect 45572 18358 45600 18634
rect 45744 18624 45796 18630
rect 45744 18566 45796 18572
rect 45560 18352 45612 18358
rect 45560 18294 45612 18300
rect 44272 18216 44324 18222
rect 44272 18158 44324 18164
rect 44180 18148 44232 18154
rect 44180 18090 44232 18096
rect 45756 17338 45784 18566
rect 45940 17338 45968 18770
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 43536 17332 43588 17338
rect 43536 17274 43588 17280
rect 45744 17332 45796 17338
rect 45744 17274 45796 17280
rect 45928 17332 45980 17338
rect 45928 17274 45980 17280
rect 46388 17332 46440 17338
rect 46388 17274 46440 17280
rect 43904 17264 43956 17270
rect 43904 17206 43956 17212
rect 44456 17264 44508 17270
rect 44456 17206 44508 17212
rect 43536 17196 43588 17202
rect 43536 17138 43588 17144
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 43548 16114 43576 17138
rect 43824 16794 43852 17138
rect 43812 16788 43864 16794
rect 43812 16730 43864 16736
rect 43720 16720 43772 16726
rect 43720 16662 43772 16668
rect 43628 16448 43680 16454
rect 43628 16390 43680 16396
rect 43640 16114 43668 16390
rect 43732 16182 43760 16662
rect 43824 16590 43852 16730
rect 43812 16584 43864 16590
rect 43812 16526 43864 16532
rect 43916 16402 43944 17206
rect 44180 17196 44232 17202
rect 44180 17138 44232 17144
rect 44192 16538 44220 17138
rect 43824 16374 43944 16402
rect 44100 16510 44220 16538
rect 43720 16176 43772 16182
rect 43720 16118 43772 16124
rect 43824 16114 43852 16374
rect 43536 16108 43588 16114
rect 43536 16050 43588 16056
rect 43628 16108 43680 16114
rect 43628 16050 43680 16056
rect 43812 16108 43864 16114
rect 43812 16050 43864 16056
rect 43996 16108 44048 16114
rect 43996 16050 44048 16056
rect 43548 15314 43576 16050
rect 43824 15450 43852 16050
rect 44008 15858 44036 16050
rect 44100 15858 44128 16510
rect 44178 16008 44234 16017
rect 44178 15943 44180 15952
rect 44232 15943 44234 15952
rect 44180 15914 44232 15920
rect 44008 15830 44220 15858
rect 43824 15422 43944 15450
rect 43812 15360 43864 15366
rect 43548 15286 43760 15314
rect 43812 15302 43864 15308
rect 43732 15026 43760 15286
rect 43824 15162 43852 15302
rect 43812 15156 43864 15162
rect 43812 15098 43864 15104
rect 43824 15026 43852 15098
rect 43916 15094 43944 15422
rect 43904 15088 43956 15094
rect 43904 15030 43956 15036
rect 44192 15026 44220 15830
rect 43720 15020 43772 15026
rect 43720 14962 43772 14968
rect 43812 15020 43864 15026
rect 43812 14962 43864 14968
rect 44088 15020 44140 15026
rect 44088 14962 44140 14968
rect 44180 15020 44232 15026
rect 44180 14962 44232 14968
rect 43732 12918 43760 14962
rect 43812 13184 43864 13190
rect 43812 13126 43864 13132
rect 43720 12912 43772 12918
rect 43720 12854 43772 12860
rect 43260 11552 43312 11558
rect 43260 11494 43312 11500
rect 43168 11008 43220 11014
rect 43168 10950 43220 10956
rect 43180 10674 43208 10950
rect 43272 10674 43300 11494
rect 43352 11144 43404 11150
rect 43352 11086 43404 11092
rect 43168 10668 43220 10674
rect 43168 10610 43220 10616
rect 43260 10668 43312 10674
rect 43260 10610 43312 10616
rect 43272 9722 43300 10610
rect 43260 9716 43312 9722
rect 43260 9658 43312 9664
rect 43260 7744 43312 7750
rect 43088 7670 43208 7698
rect 43260 7686 43312 7692
rect 42616 7472 42668 7478
rect 42616 7414 42668 7420
rect 42628 4026 42656 7414
rect 42800 7404 42852 7410
rect 42800 7346 42852 7352
rect 42812 6458 42840 7346
rect 42984 7200 43036 7206
rect 42984 7142 43036 7148
rect 42996 6798 43024 7142
rect 42984 6792 43036 6798
rect 42984 6734 43036 6740
rect 42892 6656 42944 6662
rect 42892 6598 42944 6604
rect 43076 6656 43128 6662
rect 43076 6598 43128 6604
rect 42904 6458 42932 6598
rect 42800 6452 42852 6458
rect 42800 6394 42852 6400
rect 42892 6452 42944 6458
rect 42892 6394 42944 6400
rect 43088 6322 43116 6598
rect 43076 6316 43128 6322
rect 43076 6258 43128 6264
rect 43076 6180 43128 6186
rect 43076 6122 43128 6128
rect 42892 5704 42944 5710
rect 42892 5646 42944 5652
rect 42800 5568 42852 5574
rect 42800 5510 42852 5516
rect 42812 5370 42840 5510
rect 42904 5409 42932 5646
rect 42890 5400 42946 5409
rect 42800 5364 42852 5370
rect 42890 5335 42946 5344
rect 42800 5306 42852 5312
rect 42892 4820 42944 4826
rect 42892 4762 42944 4768
rect 42904 4146 42932 4762
rect 43088 4758 43116 6122
rect 43076 4752 43128 4758
rect 43076 4694 43128 4700
rect 43088 4214 43116 4694
rect 43076 4208 43128 4214
rect 43076 4150 43128 4156
rect 42892 4140 42944 4146
rect 42892 4082 42944 4088
rect 42984 4072 43036 4078
rect 42628 4020 42984 4026
rect 42628 4014 43036 4020
rect 42628 3998 43024 4014
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 42628 3534 42656 3878
rect 42616 3528 42668 3534
rect 42616 3470 42668 3476
rect 43180 3194 43208 7670
rect 43272 3942 43300 7686
rect 43364 4978 43392 11086
rect 43536 11076 43588 11082
rect 43536 11018 43588 11024
rect 43444 10668 43496 10674
rect 43444 10610 43496 10616
rect 43456 8634 43484 10610
rect 43548 9926 43576 11018
rect 43536 9920 43588 9926
rect 43536 9862 43588 9868
rect 43628 9920 43680 9926
rect 43628 9862 43680 9868
rect 43640 9450 43668 9862
rect 43628 9444 43680 9450
rect 43628 9386 43680 9392
rect 43444 8628 43496 8634
rect 43444 8570 43496 8576
rect 43456 5710 43484 8570
rect 43628 6112 43680 6118
rect 43628 6054 43680 6060
rect 43640 5778 43668 6054
rect 43628 5772 43680 5778
rect 43628 5714 43680 5720
rect 43444 5704 43496 5710
rect 43444 5646 43496 5652
rect 43456 5166 43484 5646
rect 43628 5636 43680 5642
rect 43628 5578 43680 5584
rect 43444 5160 43496 5166
rect 43444 5102 43496 5108
rect 43364 4950 43484 4978
rect 43352 4072 43404 4078
rect 43352 4014 43404 4020
rect 43260 3936 43312 3942
rect 43260 3878 43312 3884
rect 43364 3738 43392 4014
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 43168 3188 43220 3194
rect 43168 3130 43220 3136
rect 42800 3052 42852 3058
rect 42800 2994 42852 3000
rect 42524 2440 42576 2446
rect 42524 2382 42576 2388
rect 41432 1550 41552 1578
rect 41432 800 41460 1550
rect 41880 944 41932 950
rect 41880 886 41932 892
rect 41892 800 41920 886
rect 42812 800 42840 2994
rect 43456 2446 43484 4950
rect 43640 4282 43668 5578
rect 43628 4276 43680 4282
rect 43628 4218 43680 4224
rect 43824 2514 43852 13126
rect 44100 12374 44128 14962
rect 44192 14346 44220 14962
rect 44180 14340 44232 14346
rect 44180 14282 44232 14288
rect 44088 12368 44140 12374
rect 44088 12310 44140 12316
rect 44272 11212 44324 11218
rect 44272 11154 44324 11160
rect 44284 10810 44312 11154
rect 44272 10804 44324 10810
rect 44272 10746 44324 10752
rect 43996 9716 44048 9722
rect 43996 9658 44048 9664
rect 44008 6662 44036 9658
rect 44284 6882 44312 10746
rect 44100 6854 44312 6882
rect 43996 6656 44048 6662
rect 43996 6598 44048 6604
rect 44008 5574 44036 6598
rect 44100 6458 44128 6854
rect 44272 6792 44324 6798
rect 44272 6734 44324 6740
rect 44284 6458 44312 6734
rect 44364 6656 44416 6662
rect 44364 6598 44416 6604
rect 44088 6452 44140 6458
rect 44088 6394 44140 6400
rect 44272 6452 44324 6458
rect 44272 6394 44324 6400
rect 43996 5568 44048 5574
rect 43996 5510 44048 5516
rect 44008 4826 44036 5510
rect 44100 5386 44128 6394
rect 44376 6338 44404 6598
rect 44284 6310 44404 6338
rect 44284 5914 44312 6310
rect 44272 5908 44324 5914
rect 44272 5850 44324 5856
rect 44100 5358 44220 5386
rect 44192 5166 44220 5358
rect 44180 5160 44232 5166
rect 44180 5102 44232 5108
rect 43996 4820 44048 4826
rect 43996 4762 44048 4768
rect 43996 4684 44048 4690
rect 43996 4626 44048 4632
rect 44008 4282 44036 4626
rect 43996 4276 44048 4282
rect 43996 4218 44048 4224
rect 44180 3052 44232 3058
rect 44180 2994 44232 3000
rect 43812 2508 43864 2514
rect 43812 2450 43864 2456
rect 43444 2440 43496 2446
rect 43444 2382 43496 2388
rect 42892 2372 42944 2378
rect 42892 2314 42944 2320
rect 43260 2372 43312 2378
rect 43260 2314 43312 2320
rect 42904 950 42932 2314
rect 42892 944 42944 950
rect 42892 886 42944 892
rect 43272 800 43300 2314
rect 44192 800 44220 2994
rect 44284 2310 44312 5850
rect 44364 4208 44416 4214
rect 44364 4150 44416 4156
rect 44376 3534 44404 4150
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 44376 2922 44404 3470
rect 44468 3194 44496 17206
rect 45652 17196 45704 17202
rect 45652 17138 45704 17144
rect 45468 17060 45520 17066
rect 45468 17002 45520 17008
rect 45284 16992 45336 16998
rect 45284 16934 45336 16940
rect 44916 16244 44968 16250
rect 44916 16186 44968 16192
rect 44822 5400 44878 5409
rect 44822 5335 44878 5344
rect 44640 5160 44692 5166
rect 44640 5102 44692 5108
rect 44652 4078 44680 5102
rect 44836 5030 44864 5335
rect 44824 5024 44876 5030
rect 44824 4966 44876 4972
rect 44640 4072 44692 4078
rect 44640 4014 44692 4020
rect 44928 3194 44956 16186
rect 45296 14958 45324 16934
rect 45480 16454 45508 17002
rect 45664 16590 45692 17138
rect 45756 17134 45784 17274
rect 45744 17128 45796 17134
rect 45744 17070 45796 17076
rect 46112 17128 46164 17134
rect 46112 17070 46164 17076
rect 45836 17060 45888 17066
rect 45836 17002 45888 17008
rect 45744 16652 45796 16658
rect 45744 16594 45796 16600
rect 45652 16584 45704 16590
rect 45652 16526 45704 16532
rect 45560 16516 45612 16522
rect 45560 16458 45612 16464
rect 45468 16448 45520 16454
rect 45468 16390 45520 16396
rect 45572 16250 45600 16458
rect 45560 16244 45612 16250
rect 45560 16186 45612 16192
rect 45756 16046 45784 16594
rect 45848 16046 45876 17002
rect 46124 16590 46152 17070
rect 46400 16590 46428 17274
rect 46112 16584 46164 16590
rect 46112 16526 46164 16532
rect 46388 16584 46440 16590
rect 46388 16526 46440 16532
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 45744 16040 45796 16046
rect 45744 15982 45796 15988
rect 45836 16040 45888 16046
rect 45836 15982 45888 15988
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 45284 14952 45336 14958
rect 45284 14894 45336 14900
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 53104 13524 53156 13530
rect 53104 13466 53156 13472
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 47952 12368 48004 12374
rect 47952 12310 48004 12316
rect 45284 6316 45336 6322
rect 45284 6258 45336 6264
rect 45296 5166 45324 6258
rect 45284 5160 45336 5166
rect 45284 5102 45336 5108
rect 44456 3188 44508 3194
rect 44456 3130 44508 3136
rect 44916 3188 44968 3194
rect 44916 3130 44968 3136
rect 45296 3126 45324 5102
rect 46848 4208 46900 4214
rect 46848 4150 46900 4156
rect 45284 3120 45336 3126
rect 45284 3062 45336 3068
rect 45560 3052 45612 3058
rect 45560 2994 45612 3000
rect 44364 2916 44416 2922
rect 44364 2858 44416 2864
rect 44640 2372 44692 2378
rect 44640 2314 44692 2320
rect 44272 2304 44324 2310
rect 44272 2246 44324 2252
rect 44652 800 44680 2314
rect 45572 800 45600 2994
rect 46020 2372 46072 2378
rect 46020 2314 46072 2320
rect 46032 800 46060 2314
rect 46860 1970 46888 4150
rect 47964 3194 47992 12310
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 49700 5364 49752 5370
rect 49700 5306 49752 5312
rect 47952 3188 48004 3194
rect 47952 3130 48004 3136
rect 49712 3058 49740 5306
rect 51632 5024 51684 5030
rect 51632 4966 51684 4972
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 51644 3058 51672 4966
rect 46940 3052 46992 3058
rect 46940 2994 46992 3000
rect 49700 3052 49752 3058
rect 49700 2994 49752 3000
rect 51632 3052 51684 3058
rect 51632 2994 51684 3000
rect 46848 1964 46900 1970
rect 46848 1906 46900 1912
rect 46952 800 46980 2994
rect 48780 2984 48832 2990
rect 48780 2926 48832 2932
rect 50160 2984 50212 2990
rect 50160 2926 50212 2932
rect 51540 2984 51592 2990
rect 51540 2926 51592 2932
rect 47400 2372 47452 2378
rect 47400 2314 47452 2320
rect 48320 2372 48372 2378
rect 48320 2314 48372 2320
rect 47412 800 47440 2314
rect 48332 800 48360 2314
rect 48792 800 48820 2926
rect 49700 2372 49752 2378
rect 49700 2314 49752 2320
rect 48872 2304 48924 2310
rect 48872 2246 48924 2252
rect 48884 2038 48912 2246
rect 48872 2032 48924 2038
rect 48872 1974 48924 1980
rect 49712 800 49740 2314
rect 50172 800 50200 2926
rect 51080 2372 51132 2378
rect 51080 2314 51132 2320
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 51092 800 51120 2314
rect 51448 2304 51500 2310
rect 51448 2246 51500 2252
rect 51460 1834 51488 2246
rect 51448 1828 51500 1834
rect 51448 1770 51500 1776
rect 51552 800 51580 2926
rect 53116 2650 53144 13466
rect 55956 11824 56008 11830
rect 55956 11766 56008 11772
rect 54116 8288 54168 8294
rect 54116 8230 54168 8236
rect 54128 3194 54156 8230
rect 54852 4140 54904 4146
rect 54852 4082 54904 4088
rect 54116 3188 54168 3194
rect 54116 3130 54168 3136
rect 54864 3058 54892 4082
rect 55968 3194 55996 11766
rect 56968 5296 57020 5302
rect 56968 5238 57020 5244
rect 55956 3188 56008 3194
rect 55956 3130 56008 3136
rect 56980 3126 57008 5238
rect 57060 3460 57112 3466
rect 57060 3402 57112 3408
rect 56968 3120 57020 3126
rect 56968 3062 57020 3068
rect 53840 3052 53892 3058
rect 53840 2994 53892 3000
rect 54852 3052 54904 3058
rect 54852 2994 54904 3000
rect 56600 3052 56652 3058
rect 56600 2994 56652 3000
rect 53104 2644 53156 2650
rect 53104 2586 53156 2592
rect 52460 2372 52512 2378
rect 52460 2314 52512 2320
rect 52472 800 52500 2314
rect 52920 944 52972 950
rect 52920 886 52972 892
rect 52932 800 52960 886
rect 53852 800 53880 2994
rect 54300 2984 54352 2990
rect 54300 2926 54352 2932
rect 54116 2372 54168 2378
rect 54116 2314 54168 2320
rect 54128 950 54156 2314
rect 54116 944 54168 950
rect 54116 886 54168 892
rect 54312 800 54340 2926
rect 55220 2440 55272 2446
rect 55220 2382 55272 2388
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 55232 800 55260 2382
rect 55772 2372 55824 2378
rect 55772 2314 55824 2320
rect 55784 1698 55812 2314
rect 56428 1970 56456 2382
rect 56416 1964 56468 1970
rect 56416 1906 56468 1912
rect 55772 1692 55824 1698
rect 55772 1634 55824 1640
rect 55680 944 55732 950
rect 55680 886 55732 892
rect 55692 800 55720 886
rect 56612 800 56640 2994
rect 56692 2372 56744 2378
rect 56692 2314 56744 2320
rect 56704 950 56732 2314
rect 56692 944 56744 950
rect 56692 886 56744 892
rect 57072 800 57100 3402
rect 57980 2984 58032 2990
rect 57980 2926 58032 2932
rect 57992 800 58020 2926
rect 9784 734 10088 762
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57978 0 58034 800
<< via2 >>
rect 1122 41112 1178 41168
rect 1030 40296 1086 40352
rect 938 39500 994 39536
rect 938 39480 940 39500
rect 940 39480 992 39500
rect 992 39480 994 39500
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 938 38664 994 38720
rect 938 37848 994 37904
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 938 37032 994 37088
rect 938 36216 994 36272
rect 938 35400 994 35456
rect 938 34584 994 34640
rect 938 34176 994 34232
rect 1030 33768 1086 33824
rect 938 33396 940 33416
rect 940 33396 992 33416
rect 992 33396 994 33416
rect 938 33360 994 33396
rect 1122 32952 1178 33008
rect 938 32544 994 32600
rect 938 32136 994 32192
rect 1030 31728 1086 31784
rect 938 31320 994 31376
rect 938 30912 994 30968
rect 938 30504 994 30560
rect 1030 30116 1086 30152
rect 1030 30096 1032 30116
rect 1032 30096 1084 30116
rect 1084 30096 1086 30116
rect 938 29688 994 29744
rect 938 29280 994 29336
rect 938 28872 994 28928
rect 1030 28464 1086 28520
rect 938 28056 994 28112
rect 938 27648 994 27704
rect 1030 27240 1086 27296
rect 938 26832 994 26888
rect 1030 26424 1086 26480
rect 1122 26016 1178 26072
rect 938 25608 994 25664
rect 1122 25200 1178 25256
rect 1030 24792 1086 24848
rect 938 24384 994 24440
rect 1030 23976 1086 24032
rect 1030 23568 1086 23624
rect 938 23160 994 23216
rect 938 22752 994 22808
rect 1030 22344 1086 22400
rect 938 21956 994 21992
rect 938 21936 940 21956
rect 940 21936 992 21956
rect 992 21936 994 21956
rect 938 21528 994 21584
rect 938 21120 994 21176
rect 1030 20712 1086 20768
rect 938 20340 940 20360
rect 940 20340 992 20360
rect 992 20340 994 20360
rect 938 20304 994 20340
rect 938 19916 994 19952
rect 938 19896 940 19916
rect 940 19896 992 19916
rect 992 19896 994 19916
rect 938 19488 994 19544
rect 938 19080 994 19136
rect 938 18672 994 18728
rect 1122 18264 1178 18320
rect 1030 17856 1086 17912
rect 938 17448 994 17504
rect 938 17040 994 17096
rect 938 16632 994 16688
rect 938 16224 994 16280
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1950 16088 2006 16144
rect 1122 15816 1178 15872
rect 1030 15408 1086 15464
rect 938 15000 994 15056
rect 938 14592 994 14648
rect 1030 14184 1086 14240
rect 938 13776 994 13832
rect 938 13368 994 13424
rect 938 12980 994 13016
rect 938 12960 940 12980
rect 940 12960 992 12980
rect 992 12960 994 12980
rect 938 12552 994 12608
rect 938 12180 940 12200
rect 940 12180 992 12200
rect 992 12180 994 12200
rect 938 12144 994 12180
rect 1030 11736 1086 11792
rect 938 11328 994 11384
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1122 10920 1178 10976
rect 938 10548 940 10568
rect 940 10548 992 10568
rect 992 10548 994 10568
rect 938 10512 994 10548
rect 938 9696 994 9752
rect 1030 9288 1086 9344
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 938 8064 994 8120
rect 1122 8472 1178 8528
rect 1030 7656 1086 7712
rect 938 7248 994 7304
rect 938 6840 994 6896
rect 938 6432 994 6488
rect 1030 6024 1086 6080
rect 938 5244 940 5264
rect 940 5244 992 5264
rect 992 5244 994 5264
rect 938 5208 994 5244
rect 938 4800 994 4856
rect 938 4392 994 4448
rect 938 3612 940 3632
rect 940 3612 992 3632
rect 992 3612 994 3632
rect 938 3576 994 3612
rect 938 2760 994 2816
rect 1030 2352 1086 2408
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4618 11736 4674 11792
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3790 6316 3846 6352
rect 3790 6296 3792 6316
rect 3792 6296 3844 6316
rect 3844 6296 3846 6316
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2870 1536 2926 1592
rect 3422 1944 3478 2000
rect 3330 1128 3386 1184
rect 4066 3168 4122 3224
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5814 2916 5870 2952
rect 5814 2896 5816 2916
rect 5816 2896 5868 2916
rect 5868 2896 5870 2916
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 10046 8336 10102 8392
rect 10506 5344 10562 5400
rect 1122 720 1178 776
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 13082 18808 13138 18864
rect 12898 16632 12954 16688
rect 11150 5652 11152 5672
rect 11152 5652 11204 5672
rect 11204 5652 11206 5672
rect 11150 5616 11206 5652
rect 11334 4664 11390 4720
rect 12806 2488 12862 2544
rect 15290 16532 15292 16552
rect 15292 16532 15344 16552
rect 15344 16532 15346 16552
rect 15290 16496 15346 16532
rect 15198 9580 15254 9616
rect 15198 9560 15200 9580
rect 15200 9560 15252 9580
rect 15252 9560 15254 9580
rect 15290 9424 15346 9480
rect 14646 5636 14702 5672
rect 14646 5616 14648 5636
rect 14648 5616 14700 5636
rect 14700 5616 14702 5636
rect 14830 5344 14886 5400
rect 14002 3440 14058 3496
rect 15198 3032 15254 3088
rect 15474 9580 15530 9616
rect 15474 9560 15476 9580
rect 15476 9560 15528 9580
rect 15528 9560 15530 9580
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 17038 16652 17094 16688
rect 17038 16632 17040 16652
rect 17040 16632 17092 16652
rect 17092 16632 17094 16652
rect 16486 9288 16542 9344
rect 17406 16496 17462 16552
rect 17406 9424 17462 9480
rect 16854 8336 16910 8392
rect 16762 3576 16818 3632
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 17866 9288 17922 9344
rect 17866 3576 17922 3632
rect 17406 2488 17462 2544
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19338 5208 19394 5264
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 21730 16632 21786 16688
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20626 3596 20682 3632
rect 20626 3576 20628 3596
rect 20628 3576 20680 3596
rect 20680 3576 20682 3596
rect 20350 3440 20406 3496
rect 21086 3032 21142 3088
rect 22190 11756 22246 11792
rect 22190 11736 22192 11756
rect 22192 11736 22244 11756
rect 22244 11736 22246 11756
rect 23754 15952 23810 16008
rect 23386 11736 23442 11792
rect 25318 16652 25374 16688
rect 25318 16632 25320 16652
rect 25320 16632 25372 16652
rect 25372 16632 25374 16652
rect 24674 16108 24730 16144
rect 26422 18844 26424 18864
rect 26424 18844 26476 18864
rect 26476 18844 26478 18864
rect 26422 18808 26478 18844
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 25870 16632 25926 16688
rect 24674 16088 24676 16108
rect 24676 16088 24728 16108
rect 24728 16088 24730 16108
rect 23478 11600 23534 11656
rect 23386 9968 23442 10024
rect 22282 6296 22338 6352
rect 22374 6196 22376 6216
rect 22376 6196 22428 6216
rect 22428 6196 22430 6216
rect 22374 6160 22430 6196
rect 23294 5344 23350 5400
rect 25042 6160 25098 6216
rect 24950 2896 25006 2952
rect 27158 11636 27160 11656
rect 27160 11636 27212 11656
rect 27212 11636 27214 11656
rect 27158 11600 27214 11636
rect 27526 6160 27582 6216
rect 27434 4120 27490 4176
rect 27894 5364 27950 5400
rect 27894 5344 27896 5364
rect 27896 5344 27948 5364
rect 27948 5344 27950 5364
rect 29458 15408 29514 15464
rect 30102 6740 30104 6760
rect 30104 6740 30156 6760
rect 30156 6740 30158 6760
rect 30102 6704 30158 6740
rect 29918 4684 29974 4720
rect 29918 4664 29920 4684
rect 29920 4664 29972 4684
rect 29972 4664 29974 4684
rect 29918 3848 29974 3904
rect 30010 3032 30066 3088
rect 32494 19624 32550 19680
rect 31206 3848 31262 3904
rect 32402 7404 32458 7440
rect 32402 7384 32404 7404
rect 32404 7384 32456 7404
rect 32456 7384 32458 7404
rect 32310 6724 32366 6760
rect 32310 6704 32312 6724
rect 32312 6704 32364 6724
rect 32364 6704 32366 6724
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34426 19352 34482 19408
rect 31206 3052 31262 3088
rect 31206 3032 31208 3052
rect 31208 3032 31260 3052
rect 31260 3032 31262 3052
rect 33230 7384 33286 7440
rect 32586 3984 32642 4040
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35806 17620 35808 17640
rect 35808 17620 35860 17640
rect 35860 17620 35862 17640
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35806 17584 35862 17620
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 36726 15444 36728 15464
rect 36728 15444 36780 15464
rect 36780 15444 36782 15464
rect 36726 15408 36782 15444
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38014 19624 38070 19680
rect 38566 19660 38568 19680
rect 38568 19660 38620 19680
rect 38620 19660 38622 19680
rect 38566 19624 38622 19660
rect 37738 17584 37794 17640
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 39210 9988 39266 10024
rect 39210 9968 39212 9988
rect 39212 9968 39264 9988
rect 39264 9968 39266 9988
rect 39486 9560 39542 9616
rect 42982 19352 43038 19408
rect 41786 5228 41842 5264
rect 41786 5208 41788 5228
rect 41788 5208 41840 5228
rect 41840 5208 41842 5228
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 44178 15972 44234 16008
rect 44178 15952 44180 15972
rect 44180 15952 44232 15972
rect 44232 15952 44234 15972
rect 42890 5344 42946 5400
rect 44822 5344 44878 5400
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 0 41170 800 41200
rect 1117 41170 1183 41173
rect 0 41168 1183 41170
rect 0 41112 1122 41168
rect 1178 41112 1183 41168
rect 0 41110 1183 41112
rect 0 41080 800 41110
rect 1117 41107 1183 41110
rect 0 40672 800 40792
rect 0 40354 800 40384
rect 1025 40354 1091 40357
rect 0 40352 1091 40354
rect 0 40296 1030 40352
rect 1086 40296 1091 40352
rect 0 40294 1091 40296
rect 0 40264 800 40294
rect 1025 40291 1091 40294
rect 0 39856 800 39976
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39538 800 39568
rect 933 39538 999 39541
rect 0 39536 999 39538
rect 0 39480 938 39536
rect 994 39480 999 39536
rect 0 39478 999 39480
rect 0 39448 800 39478
rect 933 39475 999 39478
rect 19570 39200 19886 39201
rect 0 39040 800 39160
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 0 38722 800 38752
rect 933 38722 999 38725
rect 0 38720 999 38722
rect 0 38664 938 38720
rect 994 38664 999 38720
rect 0 38662 999 38664
rect 0 38632 800 38662
rect 933 38659 999 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38224 800 38344
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 0 37906 800 37936
rect 933 37906 999 37909
rect 0 37904 999 37906
rect 0 37848 938 37904
rect 994 37848 999 37904
rect 0 37846 999 37848
rect 0 37816 800 37846
rect 933 37843 999 37846
rect 4210 37568 4526 37569
rect 0 37408 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 0 37090 800 37120
rect 933 37090 999 37093
rect 0 37088 999 37090
rect 0 37032 938 37088
rect 994 37032 999 37088
rect 0 37030 999 37032
rect 0 37000 800 37030
rect 933 37027 999 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36592 800 36712
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36274 800 36304
rect 933 36274 999 36277
rect 0 36272 999 36274
rect 0 36216 938 36272
rect 994 36216 999 36272
rect 0 36214 999 36216
rect 0 36184 800 36214
rect 933 36211 999 36214
rect 19570 35936 19886 35937
rect 0 35776 800 35896
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 0 35458 800 35488
rect 933 35458 999 35461
rect 0 35456 999 35458
rect 0 35400 938 35456
rect 994 35400 999 35456
rect 0 35398 999 35400
rect 0 35368 800 35398
rect 933 35395 999 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 34960 800 35080
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 0 34642 800 34672
rect 933 34642 999 34645
rect 0 34640 999 34642
rect 0 34584 938 34640
rect 994 34584 999 34640
rect 0 34582 999 34584
rect 0 34552 800 34582
rect 933 34579 999 34582
rect 4210 34304 4526 34305
rect 0 34234 800 34264
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 933 34234 999 34237
rect 0 34232 999 34234
rect 0 34176 938 34232
rect 994 34176 999 34232
rect 0 34174 999 34176
rect 0 34144 800 34174
rect 933 34171 999 34174
rect 0 33826 800 33856
rect 1025 33826 1091 33829
rect 0 33824 1091 33826
rect 0 33768 1030 33824
rect 1086 33768 1091 33824
rect 0 33766 1091 33768
rect 0 33736 800 33766
rect 1025 33763 1091 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 0 33418 800 33448
rect 933 33418 999 33421
rect 0 33416 999 33418
rect 0 33360 938 33416
rect 994 33360 999 33416
rect 0 33358 999 33360
rect 0 33328 800 33358
rect 933 33355 999 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 33010 800 33040
rect 1117 33010 1183 33013
rect 0 33008 1183 33010
rect 0 32952 1122 33008
rect 1178 32952 1183 33008
rect 0 32950 1183 32952
rect 0 32920 800 32950
rect 1117 32947 1183 32950
rect 19570 32672 19886 32673
rect 0 32602 800 32632
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 933 32602 999 32605
rect 0 32600 999 32602
rect 0 32544 938 32600
rect 994 32544 999 32600
rect 0 32542 999 32544
rect 0 32512 800 32542
rect 933 32539 999 32542
rect 0 32194 800 32224
rect 933 32194 999 32197
rect 0 32192 999 32194
rect 0 32136 938 32192
rect 994 32136 999 32192
rect 0 32134 999 32136
rect 0 32104 800 32134
rect 933 32131 999 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 0 31786 800 31816
rect 1025 31786 1091 31789
rect 0 31784 1091 31786
rect 0 31728 1030 31784
rect 1086 31728 1091 31784
rect 0 31726 1091 31728
rect 0 31696 800 31726
rect 1025 31723 1091 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 0 31378 800 31408
rect 933 31378 999 31381
rect 0 31376 999 31378
rect 0 31320 938 31376
rect 994 31320 999 31376
rect 0 31318 999 31320
rect 0 31288 800 31318
rect 933 31315 999 31318
rect 4210 31040 4526 31041
rect 0 30970 800 31000
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 933 30970 999 30973
rect 0 30968 999 30970
rect 0 30912 938 30968
rect 994 30912 999 30968
rect 0 30910 999 30912
rect 0 30880 800 30910
rect 933 30907 999 30910
rect 0 30562 800 30592
rect 933 30562 999 30565
rect 0 30560 999 30562
rect 0 30504 938 30560
rect 994 30504 999 30560
rect 0 30502 999 30504
rect 0 30472 800 30502
rect 933 30499 999 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 0 30154 800 30184
rect 1025 30154 1091 30157
rect 0 30152 1091 30154
rect 0 30096 1030 30152
rect 1086 30096 1091 30152
rect 0 30094 1091 30096
rect 0 30064 800 30094
rect 1025 30091 1091 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29746 800 29776
rect 933 29746 999 29749
rect 0 29744 999 29746
rect 0 29688 938 29744
rect 994 29688 999 29744
rect 0 29686 999 29688
rect 0 29656 800 29686
rect 933 29683 999 29686
rect 19570 29408 19886 29409
rect 0 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 933 29338 999 29341
rect 0 29336 999 29338
rect 0 29280 938 29336
rect 994 29280 999 29336
rect 0 29278 999 29280
rect 0 29248 800 29278
rect 933 29275 999 29278
rect 0 28930 800 28960
rect 933 28930 999 28933
rect 0 28928 999 28930
rect 0 28872 938 28928
rect 994 28872 999 28928
rect 0 28870 999 28872
rect 0 28840 800 28870
rect 933 28867 999 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28522 800 28552
rect 1025 28522 1091 28525
rect 0 28520 1091 28522
rect 0 28464 1030 28520
rect 1086 28464 1091 28520
rect 0 28462 1091 28464
rect 0 28432 800 28462
rect 1025 28459 1091 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 28114 800 28144
rect 933 28114 999 28117
rect 0 28112 999 28114
rect 0 28056 938 28112
rect 994 28056 999 28112
rect 0 28054 999 28056
rect 0 28024 800 28054
rect 933 28051 999 28054
rect 4210 27776 4526 27777
rect 0 27706 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 933 27706 999 27709
rect 0 27704 999 27706
rect 0 27648 938 27704
rect 994 27648 999 27704
rect 0 27646 999 27648
rect 0 27616 800 27646
rect 933 27643 999 27646
rect 0 27298 800 27328
rect 1025 27298 1091 27301
rect 0 27296 1091 27298
rect 0 27240 1030 27296
rect 1086 27240 1091 27296
rect 0 27238 1091 27240
rect 0 27208 800 27238
rect 1025 27235 1091 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 0 26890 800 26920
rect 933 26890 999 26893
rect 0 26888 999 26890
rect 0 26832 938 26888
rect 994 26832 999 26888
rect 0 26830 999 26832
rect 0 26800 800 26830
rect 933 26827 999 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 0 26482 800 26512
rect 1025 26482 1091 26485
rect 0 26480 1091 26482
rect 0 26424 1030 26480
rect 1086 26424 1091 26480
rect 0 26422 1091 26424
rect 0 26392 800 26422
rect 1025 26419 1091 26422
rect 19570 26144 19886 26145
rect 0 26074 800 26104
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 1117 26074 1183 26077
rect 0 26072 1183 26074
rect 0 26016 1122 26072
rect 1178 26016 1183 26072
rect 0 26014 1183 26016
rect 0 25984 800 26014
rect 1117 26011 1183 26014
rect 0 25666 800 25696
rect 933 25666 999 25669
rect 0 25664 999 25666
rect 0 25608 938 25664
rect 994 25608 999 25664
rect 0 25606 999 25608
rect 0 25576 800 25606
rect 933 25603 999 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 1117 25258 1183 25261
rect 0 25256 1183 25258
rect 0 25200 1122 25256
rect 1178 25200 1183 25256
rect 0 25198 1183 25200
rect 0 25168 800 25198
rect 1117 25195 1183 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24850 800 24880
rect 1025 24850 1091 24853
rect 0 24848 1091 24850
rect 0 24792 1030 24848
rect 1086 24792 1091 24848
rect 0 24790 1091 24792
rect 0 24760 800 24790
rect 1025 24787 1091 24790
rect 4210 24512 4526 24513
rect 0 24442 800 24472
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 933 24442 999 24445
rect 0 24440 999 24442
rect 0 24384 938 24440
rect 994 24384 999 24440
rect 0 24382 999 24384
rect 0 24352 800 24382
rect 933 24379 999 24382
rect 0 24034 800 24064
rect 1025 24034 1091 24037
rect 0 24032 1091 24034
rect 0 23976 1030 24032
rect 1086 23976 1091 24032
rect 0 23974 1091 23976
rect 0 23944 800 23974
rect 1025 23971 1091 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 0 23626 800 23656
rect 1025 23626 1091 23629
rect 0 23624 1091 23626
rect 0 23568 1030 23624
rect 1086 23568 1091 23624
rect 0 23566 1091 23568
rect 0 23536 800 23566
rect 1025 23563 1091 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23218 800 23248
rect 933 23218 999 23221
rect 0 23216 999 23218
rect 0 23160 938 23216
rect 994 23160 999 23216
rect 0 23158 999 23160
rect 0 23128 800 23158
rect 933 23155 999 23158
rect 19570 22880 19886 22881
rect 0 22810 800 22840
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 933 22810 999 22813
rect 0 22808 999 22810
rect 0 22752 938 22808
rect 994 22752 999 22808
rect 0 22750 999 22752
rect 0 22720 800 22750
rect 933 22747 999 22750
rect 0 22402 800 22432
rect 1025 22402 1091 22405
rect 0 22400 1091 22402
rect 0 22344 1030 22400
rect 1086 22344 1091 22400
rect 0 22342 1091 22344
rect 0 22312 800 22342
rect 1025 22339 1091 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21994 800 22024
rect 933 21994 999 21997
rect 0 21992 999 21994
rect 0 21936 938 21992
rect 994 21936 999 21992
rect 0 21934 999 21936
rect 0 21904 800 21934
rect 933 21931 999 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 0 20770 800 20800
rect 1025 20770 1091 20773
rect 0 20768 1091 20770
rect 0 20712 1030 20768
rect 1086 20712 1091 20768
rect 0 20710 1091 20712
rect 0 20680 800 20710
rect 1025 20707 1091 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 0 20362 800 20392
rect 933 20362 999 20365
rect 0 20360 999 20362
rect 0 20304 938 20360
rect 994 20304 999 20360
rect 0 20302 999 20304
rect 0 20272 800 20302
rect 933 20299 999 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19954 800 19984
rect 933 19954 999 19957
rect 0 19952 999 19954
rect 0 19896 938 19952
rect 994 19896 999 19952
rect 0 19894 999 19896
rect 0 19864 800 19894
rect 933 19891 999 19894
rect 32489 19682 32555 19685
rect 38009 19682 38075 19685
rect 38561 19682 38627 19685
rect 32489 19680 38627 19682
rect 32489 19624 32494 19680
rect 32550 19624 38014 19680
rect 38070 19624 38566 19680
rect 38622 19624 38627 19680
rect 32489 19622 38627 19624
rect 32489 19619 32555 19622
rect 38009 19619 38075 19622
rect 38561 19619 38627 19622
rect 19570 19616 19886 19617
rect 0 19546 800 19576
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 933 19546 999 19549
rect 0 19544 999 19546
rect 0 19488 938 19544
rect 994 19488 999 19544
rect 0 19486 999 19488
rect 0 19456 800 19486
rect 933 19483 999 19486
rect 34421 19410 34487 19413
rect 42977 19410 43043 19413
rect 34421 19408 43043 19410
rect 34421 19352 34426 19408
rect 34482 19352 42982 19408
rect 43038 19352 43043 19408
rect 34421 19350 43043 19352
rect 34421 19347 34487 19350
rect 42977 19347 43043 19350
rect 0 19138 800 19168
rect 933 19138 999 19141
rect 0 19136 999 19138
rect 0 19080 938 19136
rect 994 19080 999 19136
rect 0 19078 999 19080
rect 0 19048 800 19078
rect 933 19075 999 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 13077 18866 13143 18869
rect 26417 18866 26483 18869
rect 13077 18864 26483 18866
rect 13077 18808 13082 18864
rect 13138 18808 26422 18864
rect 26478 18808 26483 18864
rect 13077 18806 26483 18808
rect 13077 18803 13143 18806
rect 26417 18803 26483 18806
rect 0 18730 800 18760
rect 933 18730 999 18733
rect 0 18728 999 18730
rect 0 18672 938 18728
rect 994 18672 999 18728
rect 0 18670 999 18672
rect 0 18640 800 18670
rect 933 18667 999 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 0 18322 800 18352
rect 1117 18322 1183 18325
rect 0 18320 1183 18322
rect 0 18264 1122 18320
rect 1178 18264 1183 18320
rect 0 18262 1183 18264
rect 0 18232 800 18262
rect 1117 18259 1183 18262
rect 4210 17984 4526 17985
rect 0 17914 800 17944
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 1025 17914 1091 17917
rect 0 17912 1091 17914
rect 0 17856 1030 17912
rect 1086 17856 1091 17912
rect 0 17854 1091 17856
rect 0 17824 800 17854
rect 1025 17851 1091 17854
rect 35801 17642 35867 17645
rect 37733 17642 37799 17645
rect 35801 17640 37799 17642
rect 35801 17584 35806 17640
rect 35862 17584 37738 17640
rect 37794 17584 37799 17640
rect 35801 17582 37799 17584
rect 35801 17579 35867 17582
rect 37733 17579 37799 17582
rect 0 17506 800 17536
rect 933 17506 999 17509
rect 0 17504 999 17506
rect 0 17448 938 17504
rect 994 17448 999 17504
rect 0 17446 999 17448
rect 0 17416 800 17446
rect 933 17443 999 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16690 800 16720
rect 933 16690 999 16693
rect 0 16688 999 16690
rect 0 16632 938 16688
rect 994 16632 999 16688
rect 0 16630 999 16632
rect 0 16600 800 16630
rect 933 16627 999 16630
rect 12893 16690 12959 16693
rect 17033 16690 17099 16693
rect 12893 16688 17099 16690
rect 12893 16632 12898 16688
rect 12954 16632 17038 16688
rect 17094 16632 17099 16688
rect 12893 16630 17099 16632
rect 12893 16627 12959 16630
rect 17033 16627 17099 16630
rect 21725 16690 21791 16693
rect 25313 16690 25379 16693
rect 25865 16690 25931 16693
rect 21725 16688 25931 16690
rect 21725 16632 21730 16688
rect 21786 16632 25318 16688
rect 25374 16632 25870 16688
rect 25926 16632 25931 16688
rect 21725 16630 25931 16632
rect 21725 16627 21791 16630
rect 25313 16627 25379 16630
rect 25865 16627 25931 16630
rect 15285 16554 15351 16557
rect 17401 16554 17467 16557
rect 15285 16552 17467 16554
rect 15285 16496 15290 16552
rect 15346 16496 17406 16552
rect 17462 16496 17467 16552
rect 15285 16494 17467 16496
rect 15285 16491 15351 16494
rect 17401 16491 17467 16494
rect 19570 16352 19886 16353
rect 0 16282 800 16312
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 933 16282 999 16285
rect 0 16280 999 16282
rect 0 16224 938 16280
rect 994 16224 999 16280
rect 0 16222 999 16224
rect 0 16192 800 16222
rect 933 16219 999 16222
rect 1945 16146 2011 16149
rect 24669 16146 24735 16149
rect 1945 16144 24735 16146
rect 1945 16088 1950 16144
rect 2006 16088 24674 16144
rect 24730 16088 24735 16144
rect 1945 16086 24735 16088
rect 1945 16083 2011 16086
rect 24669 16083 24735 16086
rect 23749 16010 23815 16013
rect 44173 16010 44239 16013
rect 23749 16008 44239 16010
rect 23749 15952 23754 16008
rect 23810 15952 44178 16008
rect 44234 15952 44239 16008
rect 23749 15950 44239 15952
rect 23749 15947 23815 15950
rect 44173 15947 44239 15950
rect 0 15874 800 15904
rect 1117 15874 1183 15877
rect 0 15872 1183 15874
rect 0 15816 1122 15872
rect 1178 15816 1183 15872
rect 0 15814 1183 15816
rect 0 15784 800 15814
rect 1117 15811 1183 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 0 15466 800 15496
rect 1025 15466 1091 15469
rect 0 15464 1091 15466
rect 0 15408 1030 15464
rect 1086 15408 1091 15464
rect 0 15406 1091 15408
rect 0 15376 800 15406
rect 1025 15403 1091 15406
rect 29453 15466 29519 15469
rect 36721 15466 36787 15469
rect 29453 15464 36787 15466
rect 29453 15408 29458 15464
rect 29514 15408 36726 15464
rect 36782 15408 36787 15464
rect 29453 15406 36787 15408
rect 29453 15403 29519 15406
rect 36721 15403 36787 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 4210 14720 4526 14721
rect 0 14650 800 14680
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 933 14650 999 14653
rect 0 14648 999 14650
rect 0 14592 938 14648
rect 994 14592 999 14648
rect 0 14590 999 14592
rect 0 14560 800 14590
rect 933 14587 999 14590
rect 0 14242 800 14272
rect 1025 14242 1091 14245
rect 0 14240 1091 14242
rect 0 14184 1030 14240
rect 1086 14184 1091 14240
rect 0 14182 1091 14184
rect 0 14152 800 14182
rect 1025 14179 1091 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 0 13834 800 13864
rect 933 13834 999 13837
rect 0 13832 999 13834
rect 0 13776 938 13832
rect 994 13776 999 13832
rect 0 13774 999 13776
rect 0 13744 800 13774
rect 933 13771 999 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 0 13426 800 13456
rect 933 13426 999 13429
rect 0 13424 999 13426
rect 0 13368 938 13424
rect 994 13368 999 13424
rect 0 13366 999 13368
rect 0 13336 800 13366
rect 933 13363 999 13366
rect 19570 13088 19886 13089
rect 0 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 0 12610 800 12640
rect 933 12610 999 12613
rect 0 12608 999 12610
rect 0 12552 938 12608
rect 994 12552 999 12608
rect 0 12550 999 12552
rect 0 12520 800 12550
rect 933 12547 999 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12202 800 12232
rect 933 12202 999 12205
rect 0 12200 999 12202
rect 0 12144 938 12200
rect 994 12144 999 12200
rect 0 12142 999 12144
rect 0 12112 800 12142
rect 933 12139 999 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11794 800 11824
rect 1025 11794 1091 11797
rect 0 11792 1091 11794
rect 0 11736 1030 11792
rect 1086 11736 1091 11792
rect 0 11734 1091 11736
rect 0 11704 800 11734
rect 1025 11731 1091 11734
rect 4613 11794 4679 11797
rect 22185 11794 22251 11797
rect 23381 11794 23447 11797
rect 4613 11792 23447 11794
rect 4613 11736 4618 11792
rect 4674 11736 22190 11792
rect 22246 11736 23386 11792
rect 23442 11736 23447 11792
rect 4613 11734 23447 11736
rect 4613 11731 4679 11734
rect 22185 11731 22251 11734
rect 23381 11731 23447 11734
rect 23473 11658 23539 11661
rect 27153 11658 27219 11661
rect 23473 11656 27219 11658
rect 23473 11600 23478 11656
rect 23534 11600 27158 11656
rect 27214 11600 27219 11656
rect 23473 11598 27219 11600
rect 23473 11595 23539 11598
rect 27153 11595 27219 11598
rect 4210 11456 4526 11457
rect 0 11386 800 11416
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 933 11386 999 11389
rect 0 11384 999 11386
rect 0 11328 938 11384
rect 994 11328 999 11384
rect 0 11326 999 11328
rect 0 11296 800 11326
rect 933 11323 999 11326
rect 0 10978 800 11008
rect 1117 10978 1183 10981
rect 0 10976 1183 10978
rect 0 10920 1122 10976
rect 1178 10920 1183 10976
rect 0 10918 1183 10920
rect 0 10888 800 10918
rect 1117 10915 1183 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 0 10570 800 10600
rect 933 10570 999 10573
rect 0 10568 999 10570
rect 0 10512 938 10568
rect 994 10512 999 10568
rect 0 10510 999 10512
rect 0 10480 800 10510
rect 933 10507 999 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 0 10072 800 10192
rect 23381 10026 23447 10029
rect 39205 10026 39271 10029
rect 23381 10024 39271 10026
rect 23381 9968 23386 10024
rect 23442 9968 39210 10024
rect 39266 9968 39271 10024
rect 23381 9966 39271 9968
rect 23381 9963 23447 9966
rect 39205 9963 39271 9966
rect 19570 9824 19886 9825
rect 0 9754 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 933 9754 999 9757
rect 0 9752 999 9754
rect 0 9696 938 9752
rect 994 9696 999 9752
rect 0 9694 999 9696
rect 0 9664 800 9694
rect 933 9691 999 9694
rect 15193 9618 15259 9621
rect 15469 9618 15535 9621
rect 39481 9618 39547 9621
rect 15193 9616 39547 9618
rect 15193 9560 15198 9616
rect 15254 9560 15474 9616
rect 15530 9560 39486 9616
rect 39542 9560 39547 9616
rect 15193 9558 39547 9560
rect 15193 9555 15259 9558
rect 15469 9555 15535 9558
rect 39481 9555 39547 9558
rect 15285 9482 15351 9485
rect 17401 9482 17467 9485
rect 15285 9480 17467 9482
rect 15285 9424 15290 9480
rect 15346 9424 17406 9480
rect 17462 9424 17467 9480
rect 15285 9422 17467 9424
rect 15285 9419 15351 9422
rect 17401 9419 17467 9422
rect 0 9346 800 9376
rect 1025 9346 1091 9349
rect 0 9344 1091 9346
rect 0 9288 1030 9344
rect 1086 9288 1091 9344
rect 0 9286 1091 9288
rect 0 9256 800 9286
rect 1025 9283 1091 9286
rect 16481 9346 16547 9349
rect 17861 9346 17927 9349
rect 16481 9344 17927 9346
rect 16481 9288 16486 9344
rect 16542 9288 17866 9344
rect 17922 9288 17927 9344
rect 16481 9286 17927 9288
rect 16481 9283 16547 9286
rect 17861 9283 17927 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 0 8530 800 8560
rect 1117 8530 1183 8533
rect 0 8528 1183 8530
rect 0 8472 1122 8528
rect 1178 8472 1183 8528
rect 0 8470 1183 8472
rect 0 8440 800 8470
rect 1117 8467 1183 8470
rect 10041 8394 10107 8397
rect 16849 8394 16915 8397
rect 10041 8392 16915 8394
rect 10041 8336 10046 8392
rect 10102 8336 16854 8392
rect 16910 8336 16915 8392
rect 10041 8334 16915 8336
rect 10041 8331 10107 8334
rect 16849 8331 16915 8334
rect 4210 8192 4526 8193
rect 0 8122 800 8152
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 933 8122 999 8125
rect 0 8120 999 8122
rect 0 8064 938 8120
rect 994 8064 999 8120
rect 0 8062 999 8064
rect 0 8032 800 8062
rect 933 8059 999 8062
rect 0 7714 800 7744
rect 1025 7714 1091 7717
rect 0 7712 1091 7714
rect 0 7656 1030 7712
rect 1086 7656 1091 7712
rect 0 7654 1091 7656
rect 0 7624 800 7654
rect 1025 7651 1091 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 32397 7442 32463 7445
rect 33225 7442 33291 7445
rect 32397 7440 33291 7442
rect 32397 7384 32402 7440
rect 32458 7384 33230 7440
rect 33286 7384 33291 7440
rect 32397 7382 33291 7384
rect 32397 7379 32463 7382
rect 33225 7379 33291 7382
rect 0 7306 800 7336
rect 933 7306 999 7309
rect 0 7304 999 7306
rect 0 7248 938 7304
rect 994 7248 999 7304
rect 0 7246 999 7248
rect 0 7216 800 7246
rect 933 7243 999 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 30097 6762 30163 6765
rect 32305 6762 32371 6765
rect 30097 6760 32371 6762
rect 30097 6704 30102 6760
rect 30158 6704 32310 6760
rect 32366 6704 32371 6760
rect 30097 6702 32371 6704
rect 30097 6699 30163 6702
rect 32305 6699 32371 6702
rect 19570 6560 19886 6561
rect 0 6490 800 6520
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 933 6490 999 6493
rect 0 6488 999 6490
rect 0 6432 938 6488
rect 994 6432 999 6488
rect 0 6430 999 6432
rect 0 6400 800 6430
rect 933 6427 999 6430
rect 3785 6354 3851 6357
rect 22277 6354 22343 6357
rect 3785 6352 22343 6354
rect 3785 6296 3790 6352
rect 3846 6296 22282 6352
rect 22338 6296 22343 6352
rect 3785 6294 22343 6296
rect 3785 6291 3851 6294
rect 22277 6291 22343 6294
rect 22369 6218 22435 6221
rect 25037 6218 25103 6221
rect 27521 6218 27587 6221
rect 22369 6216 27587 6218
rect 22369 6160 22374 6216
rect 22430 6160 25042 6216
rect 25098 6160 27526 6216
rect 27582 6160 27587 6216
rect 22369 6158 27587 6160
rect 22369 6155 22435 6158
rect 25037 6155 25103 6158
rect 27521 6155 27587 6158
rect 0 6082 800 6112
rect 1025 6082 1091 6085
rect 0 6080 1091 6082
rect 0 6024 1030 6080
rect 1086 6024 1091 6080
rect 0 6022 1091 6024
rect 0 5992 800 6022
rect 1025 6019 1091 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5584 800 5704
rect 11145 5674 11211 5677
rect 14641 5674 14707 5677
rect 11145 5672 14707 5674
rect 11145 5616 11150 5672
rect 11206 5616 14646 5672
rect 14702 5616 14707 5672
rect 11145 5614 14707 5616
rect 11145 5611 11211 5614
rect 14641 5611 14707 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 10501 5402 10567 5405
rect 14825 5402 14891 5405
rect 10501 5400 14891 5402
rect 10501 5344 10506 5400
rect 10562 5344 14830 5400
rect 14886 5344 14891 5400
rect 10501 5342 14891 5344
rect 10501 5339 10567 5342
rect 14825 5339 14891 5342
rect 23289 5402 23355 5405
rect 27889 5402 27955 5405
rect 23289 5400 27955 5402
rect 23289 5344 23294 5400
rect 23350 5344 27894 5400
rect 27950 5344 27955 5400
rect 23289 5342 27955 5344
rect 23289 5339 23355 5342
rect 27889 5339 27955 5342
rect 42885 5402 42951 5405
rect 44817 5402 44883 5405
rect 42885 5400 44883 5402
rect 42885 5344 42890 5400
rect 42946 5344 44822 5400
rect 44878 5344 44883 5400
rect 42885 5342 44883 5344
rect 42885 5339 42951 5342
rect 44817 5339 44883 5342
rect 0 5266 800 5296
rect 933 5266 999 5269
rect 0 5264 999 5266
rect 0 5208 938 5264
rect 994 5208 999 5264
rect 0 5206 999 5208
rect 0 5176 800 5206
rect 933 5203 999 5206
rect 19333 5266 19399 5269
rect 41781 5266 41847 5269
rect 19333 5264 41847 5266
rect 19333 5208 19338 5264
rect 19394 5208 41786 5264
rect 41842 5208 41847 5264
rect 19333 5206 41847 5208
rect 19333 5203 19399 5206
rect 41781 5203 41847 5206
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 11329 4722 11395 4725
rect 29913 4722 29979 4725
rect 11329 4720 29979 4722
rect 11329 4664 11334 4720
rect 11390 4664 29918 4720
rect 29974 4664 29979 4720
rect 11329 4662 29979 4664
rect 11329 4659 11395 4662
rect 29913 4659 29979 4662
rect 0 4450 800 4480
rect 933 4450 999 4453
rect 0 4448 999 4450
rect 0 4392 938 4448
rect 994 4392 999 4448
rect 0 4390 999 4392
rect 0 4360 800 4390
rect 933 4387 999 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 27429 4178 27495 4181
rect 27429 4176 27538 4178
rect 27429 4120 27434 4176
rect 27490 4120 27538 4176
rect 27429 4115 27538 4120
rect 0 3952 800 4072
rect 27478 4042 27538 4115
rect 32581 4042 32647 4045
rect 27478 4040 32647 4042
rect 27478 3984 32586 4040
rect 32642 3984 32647 4040
rect 27478 3982 32647 3984
rect 32581 3979 32647 3982
rect 29913 3906 29979 3909
rect 31201 3906 31267 3909
rect 29913 3904 31267 3906
rect 29913 3848 29918 3904
rect 29974 3848 31206 3904
rect 31262 3848 31267 3904
rect 29913 3846 31267 3848
rect 29913 3843 29979 3846
rect 31201 3843 31267 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 16757 3634 16823 3637
rect 17861 3634 17927 3637
rect 20621 3634 20687 3637
rect 16757 3632 20687 3634
rect 16757 3576 16762 3632
rect 16818 3576 17866 3632
rect 17922 3576 20626 3632
rect 20682 3576 20687 3632
rect 16757 3574 20687 3576
rect 16757 3571 16823 3574
rect 17861 3571 17927 3574
rect 20621 3571 20687 3574
rect 13997 3498 14063 3501
rect 20345 3498 20411 3501
rect 13997 3496 20411 3498
rect 13997 3440 14002 3496
rect 14058 3440 20350 3496
rect 20406 3440 20411 3496
rect 13997 3438 20411 3440
rect 13997 3435 14063 3438
rect 20345 3435 20411 3438
rect 19570 3296 19886 3297
rect 0 3226 800 3256
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4061 3226 4127 3229
rect 0 3224 4127 3226
rect 0 3168 4066 3224
rect 4122 3168 4127 3224
rect 0 3166 4127 3168
rect 0 3136 800 3166
rect 4061 3163 4127 3166
rect 15193 3090 15259 3093
rect 21081 3090 21147 3093
rect 15193 3088 21147 3090
rect 15193 3032 15198 3088
rect 15254 3032 21086 3088
rect 21142 3032 21147 3088
rect 15193 3030 21147 3032
rect 15193 3027 15259 3030
rect 21081 3027 21147 3030
rect 30005 3090 30071 3093
rect 31201 3090 31267 3093
rect 30005 3088 31267 3090
rect 30005 3032 30010 3088
rect 30066 3032 31206 3088
rect 31262 3032 31267 3088
rect 30005 3030 31267 3032
rect 30005 3027 30071 3030
rect 31201 3027 31267 3030
rect 5809 2954 5875 2957
rect 24945 2954 25011 2957
rect 5809 2952 25011 2954
rect 5809 2896 5814 2952
rect 5870 2896 24950 2952
rect 25006 2896 25011 2952
rect 5809 2894 25011 2896
rect 5809 2891 5875 2894
rect 24945 2891 25011 2894
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 12801 2546 12867 2549
rect 17401 2546 17467 2549
rect 12801 2544 17467 2546
rect 12801 2488 12806 2544
rect 12862 2488 17406 2544
rect 17462 2488 17467 2544
rect 12801 2486 17467 2488
rect 12801 2483 12867 2486
rect 17401 2483 17467 2486
rect 0 2410 800 2440
rect 1025 2410 1091 2413
rect 0 2408 1091 2410
rect 0 2352 1030 2408
rect 1086 2352 1091 2408
rect 0 2350 1091 2352
rect 0 2320 800 2350
rect 1025 2347 1091 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 0 2002 800 2032
rect 3417 2002 3483 2005
rect 0 2000 3483 2002
rect 0 1944 3422 2000
rect 3478 1944 3483 2000
rect 0 1942 3483 1944
rect 0 1912 800 1942
rect 3417 1939 3483 1942
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
rect 0 1186 800 1216
rect 3325 1186 3391 1189
rect 0 1184 3391 1186
rect 0 1128 3330 1184
rect 3386 1128 3391 1184
rect 0 1126 3391 1128
rect 0 1096 800 1126
rect 3325 1123 3391 1126
rect 0 778 800 808
rect 1117 778 1183 781
rect 0 776 1183 778
rect 0 720 1122 776
rect 1178 720 1183 776
rect 0 718 1183 720
rect 0 688 800 718
rect 1117 715 1183 718
<< via3 >>
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 39744 4528 39760
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 39200 19888 39760
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 39744 35248 39760
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 39200 50608 39760
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 27600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 27876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1676037725
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1676037725
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1676037725
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1676037725
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1676037725
transform 1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_263
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1676037725
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1676037725
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_317
timestamp 1676037725
transform 1 0 30268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_323
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_353
timestamp 1676037725
transform 1 0 33580 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1676037725
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1676037725
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1676037725
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_413
timestamp 1676037725
transform 1 0 39100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1676037725
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_495
timestamp 1676037725
transform 1 0 46644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1676037725
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1676037725
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_541
timestamp 1676037725
transform 1 0 50876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_551
timestamp 1676037725
transform 1 0 51796 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1676037725
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_569
timestamp 1676037725
transform 1 0 53452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_579
timestamp 1676037725
transform 1 0 54372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1676037725
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_597
timestamp 1676037725
transform 1 0 56028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_607
timestamp 1676037725
transform 1 0 56948 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1676037725
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1676037725
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1676037725
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_70
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_76
timestamp 1676037725
transform 1 0 8096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1676037725
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 1676037725
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1676037725
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1676037725
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1676037725
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1676037725
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1676037725
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_250
timestamp 1676037725
transform 1 0 24104 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_258
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_265 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_288
timestamp 1676037725
transform 1 0 27600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1676037725
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_316
timestamp 1676037725
transform 1 0 30176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1676037725
transform 1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_347
timestamp 1676037725
transform 1 0 33028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_352
timestamp 1676037725
transform 1 0 33488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_381
timestamp 1676037725
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1676037725
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_399
timestamp 1676037725
transform 1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_419
timestamp 1676037725
transform 1 0 39652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_427
timestamp 1676037725
transform 1 0 40388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1676037725
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_455
timestamp 1676037725
transform 1 0 42964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_463
timestamp 1676037725
transform 1 0 43700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_481
timestamp 1676037725
transform 1 0 45356 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_488
timestamp 1676037725
transform 1 0 46000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1676037725
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_511
timestamp 1676037725
transform 1 0 48116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_533
timestamp 1676037725
transform 1 0 50140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_540
timestamp 1676037725
transform 1 0 50784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_548
timestamp 1676037725
transform 1 0 51520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1676037725
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_573
timestamp 1676037725
transform 1 0 53820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_580
timestamp 1676037725
transform 1 0 54464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_590
timestamp 1676037725
transform 1 0 55384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_600
timestamp 1676037725
transform 1 0 56304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_610
timestamp 1676037725
transform 1 0 57224 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 1676037725
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1676037725
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1676037725
transform 1 0 5336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1676037725
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1676037725
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_126
timestamp 1676037725
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_148
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1676037725
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1676037725
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_184
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_203
timestamp 1676037725
transform 1 0 19780 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_218
timestamp 1676037725
transform 1 0 21160 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_228
timestamp 1676037725
transform 1 0 22080 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_284
timestamp 1676037725
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1676037725
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_297
timestamp 1676037725
transform 1 0 28428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1676037725
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_318
timestamp 1676037725
transform 1 0 30360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1676037725
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_352
timestamp 1676037725
transform 1 0 33488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_374
timestamp 1676037725
transform 1 0 35512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_395
timestamp 1676037725
transform 1 0 37444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1676037725
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_428
timestamp 1676037725
transform 1 0 40480 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_450
timestamp 1676037725
transform 1 0 42504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_462
timestamp 1676037725
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1676037725
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1676037725
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1676037725
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1676037725
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1676037725
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_601
timestamp 1676037725
transform 1 0 56396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_615
timestamp 1676037725
transform 1 0 57684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_623
timestamp 1676037725
transform 1 0 58420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1676037725
transform 1 0 4968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1676037725
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_82
timestamp 1676037725
transform 1 0 8648 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_94
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1676037725
transform 1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_150
timestamp 1676037725
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1676037725
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1676037725
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_199
timestamp 1676037725
transform 1 0 19412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1676037725
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1676037725
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1676037725
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_315
timestamp 1676037725
transform 1 0 30084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_323
timestamp 1676037725
transform 1 0 30820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1676037725
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_350
timestamp 1676037725
transform 1 0 33304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_362
timestamp 1676037725
transform 1 0 34408 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_368
timestamp 1676037725
transform 1 0 34960 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_380
timestamp 1676037725
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_413
timestamp 1676037725
transform 1 0 39100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_425
timestamp 1676037725
transform 1 0 40204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_437
timestamp 1676037725
transform 1 0 41308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_445
timestamp 1676037725
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_459
timestamp 1676037725
transform 1 0 43332 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_465
timestamp 1676037725
transform 1 0 43884 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_475
timestamp 1676037725
transform 1 0 44804 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_488
timestamp 1676037725
transform 1 0 46000 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1676037725
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1676037725
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_35
timestamp 1676037725
transform 1 0 4324 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1676037725
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_59
timestamp 1676037725
transform 1 0 6532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_115
timestamp 1676037725
transform 1 0 11684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_127
timestamp 1676037725
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_161
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1676037725
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_182
timestamp 1676037725
transform 1 0 17848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1676037725
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1676037725
transform 1 0 20056 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_213
timestamp 1676037725
transform 1 0 20700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_225
timestamp 1676037725
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_231
timestamp 1676037725
transform 1 0 22356 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_239
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_271
timestamp 1676037725
transform 1 0 26036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_318
timestamp 1676037725
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_330
timestamp 1676037725
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_342
timestamp 1676037725
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp 1676037725
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1676037725
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_405
timestamp 1676037725
transform 1 0 38364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1676037725
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_437
timestamp 1676037725
transform 1 0 41308 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_446
timestamp 1676037725
transform 1 0 42136 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_458
timestamp 1676037725
transform 1 0 43240 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_470
timestamp 1676037725
transform 1 0 44344 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_19
timestamp 1676037725
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_44
timestamp 1676037725
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp 1676037725
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_80
timestamp 1676037725
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_92
timestamp 1676037725
transform 1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1676037725
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1676037725
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_148
timestamp 1676037725
transform 1 0 14720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_156
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1676037725
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_176
timestamp 1676037725
transform 1 0 17296 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1676037725
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_245
timestamp 1676037725
transform 1 0 23644 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_255
timestamp 1676037725
transform 1 0 24564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_267
timestamp 1676037725
transform 1 0 25668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_291
timestamp 1676037725
transform 1 0 27876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_303
timestamp 1676037725
transform 1 0 28980 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1676037725
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1676037725
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_377
timestamp 1676037725
transform 1 0 35788 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1676037725
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1676037725
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_471
timestamp 1676037725
transform 1 0 44436 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_484
timestamp 1676037725
transform 1 0 45632 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_496
timestamp 1676037725
transform 1 0 46736 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1676037725
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_35
timestamp 1676037725
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1676037725
transform 1 0 5060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1676037725
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1676037725
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1676037725
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1676037725
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_125
timestamp 1676037725
transform 1 0 12604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1676037725
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_149
timestamp 1676037725
transform 1 0 14812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_161
timestamp 1676037725
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_185
timestamp 1676037725
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1676037725
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_216
timestamp 1676037725
transform 1 0 20976 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_228
timestamp 1676037725
transform 1 0 22080 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_239
timestamp 1676037725
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_269
timestamp 1676037725
transform 1 0 25852 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_287
timestamp 1676037725
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1676037725
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_334
timestamp 1676037725
transform 1 0 31832 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_346
timestamp 1676037725
transform 1 0 32936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_399
timestamp 1676037725
transform 1 0 37812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_411
timestamp 1676037725
transform 1 0 38916 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_430
timestamp 1676037725
transform 1 0 40664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_434
timestamp 1676037725
transform 1 0 41032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_451
timestamp 1676037725
transform 1 0 42596 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_463
timestamp 1676037725
transform 1 0 43700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1676037725
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1676037725
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1676037725
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_72
timestamp 1676037725
transform 1 0 7728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1676037725
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1676037725
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1676037725
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1676037725
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_122
timestamp 1676037725
transform 1 0 12328 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1676037725
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1676037725
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_144
timestamp 1676037725
transform 1 0 14352 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_156
timestamp 1676037725
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_200
timestamp 1676037725
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1676037725
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_236
timestamp 1676037725
transform 1 0 22816 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_248
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_260
timestamp 1676037725
transform 1 0 25024 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1676037725
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_312
timestamp 1676037725
transform 1 0 29808 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_324
timestamp 1676037725
transform 1 0 30912 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_355
timestamp 1676037725
transform 1 0 33764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_404
timestamp 1676037725
transform 1 0 38272 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_425
timestamp 1676037725
transform 1 0 40204 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_437
timestamp 1676037725
transform 1 0 41308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_445
timestamp 1676037725
transform 1 0 42044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_458
timestamp 1676037725
transform 1 0 43240 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_464
timestamp 1676037725
transform 1 0 43792 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_470
timestamp 1676037725
transform 1 0 44344 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_482
timestamp 1676037725
transform 1 0 45448 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_494
timestamp 1676037725
transform 1 0 46552 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_502
timestamp 1676037725
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_35
timestamp 1676037725
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_59
timestamp 1676037725
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_71
timestamp 1676037725
transform 1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp 1676037725
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1676037725
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1676037725
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1676037725
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_258
timestamp 1676037725
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_270
timestamp 1676037725
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_282
timestamp 1676037725
transform 1 0 27048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1676037725
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1676037725
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_320
timestamp 1676037725
transform 1 0 30544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1676037725
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_340
timestamp 1676037725
transform 1 0 32384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_344
timestamp 1676037725
transform 1 0 32752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1676037725
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_378
timestamp 1676037725
transform 1 0 35880 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_387
timestamp 1676037725
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_399
timestamp 1676037725
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_411
timestamp 1676037725
transform 1 0 38916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_453
timestamp 1676037725
transform 1 0 42780 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_461
timestamp 1676037725
transform 1 0 43516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_471
timestamp 1676037725
transform 1 0 44436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_18
timestamp 1676037725
transform 1 0 2760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_26
timestamp 1676037725
transform 1 0 3496 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp 1676037725
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_43
timestamp 1676037725
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1676037725
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1676037725
transform 1 0 9752 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1676037725
transform 1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_120
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_132
timestamp 1676037725
transform 1 0 13248 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_148
timestamp 1676037725
transform 1 0 14720 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_202
timestamp 1676037725
transform 1 0 19688 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1676037725
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1676037725
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_242
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_254
timestamp 1676037725
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_347
timestamp 1676037725
transform 1 0 33028 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_354
timestamp 1676037725
transform 1 0 33672 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_366
timestamp 1676037725
transform 1 0 34776 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_378
timestamp 1676037725
transform 1 0 35880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_397
timestamp 1676037725
transform 1 0 37628 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_407
timestamp 1676037725
transform 1 0 38548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_419
timestamp 1676037725
transform 1 0 39652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_431
timestamp 1676037725
transform 1 0 40756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_443
timestamp 1676037725
transform 1 0 41860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_456
timestamp 1676037725
transform 1 0 43056 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_468
timestamp 1676037725
transform 1 0 44160 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_480
timestamp 1676037725
transform 1 0 45264 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_492
timestamp 1676037725
transform 1 0 46368 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1676037725
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1676037725
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1676037725
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1676037725
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_47
timestamp 1676037725
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_59
timestamp 1676037725
transform 1 0 6532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1676037725
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1676037725
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_112
timestamp 1676037725
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_130
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_164
timestamp 1676037725
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_176
timestamp 1676037725
transform 1 0 17296 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_184
timestamp 1676037725
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1676037725
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_225
timestamp 1676037725
transform 1 0 21804 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_237
timestamp 1676037725
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1676037725
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_285
timestamp 1676037725
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_297
timestamp 1676037725
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1676037725
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_329
timestamp 1676037725
transform 1 0 31372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_335
timestamp 1676037725
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_346
timestamp 1676037725
transform 1 0 32936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_356
timestamp 1676037725
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_374
timestamp 1676037725
transform 1 0 35512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_378
timestamp 1676037725
transform 1 0 35880 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_395
timestamp 1676037725
transform 1 0 37444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_407
timestamp 1676037725
transform 1 0 38548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_430
timestamp 1676037725
transform 1 0 40664 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_453
timestamp 1676037725
transform 1 0 42780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_465
timestamp 1676037725
transform 1 0 43884 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_473
timestamp 1676037725
transform 1 0 44620 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1676037725
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1676037725
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1676037725
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_65
timestamp 1676037725
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_76
timestamp 1676037725
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_88
timestamp 1676037725
transform 1 0 9200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_96
timestamp 1676037725
transform 1 0 9936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1676037725
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_127
timestamp 1676037725
transform 1 0 12788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1676037725
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_155
timestamp 1676037725
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1676037725
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp 1676037725
transform 1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_211
timestamp 1676037725
transform 1 0 20516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_233
timestamp 1676037725
transform 1 0 22540 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_250
timestamp 1676037725
transform 1 0 24104 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_258
timestamp 1676037725
transform 1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1676037725
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_346
timestamp 1676037725
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_356
timestamp 1676037725
transform 1 0 33856 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_368
timestamp 1676037725
transform 1 0 34960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1676037725
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1676037725
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_400
timestamp 1676037725
transform 1 0 37904 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_412
timestamp 1676037725
transform 1 0 39008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_419
timestamp 1676037725
transform 1 0 39652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_428
timestamp 1676037725
transform 1 0 40480 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_435
timestamp 1676037725
transform 1 0 41124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1676037725
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1676037725
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1676037725
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1676037725
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1676037725
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1676037725
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_104
timestamp 1676037725
transform 1 0 10672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1676037725
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_184
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_205
timestamp 1676037725
transform 1 0 19964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1676037725
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1676037725
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_295
timestamp 1676037725
transform 1 0 28244 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1676037725
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_327
timestamp 1676037725
transform 1 0 31188 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_336
timestamp 1676037725
transform 1 0 32016 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_348
timestamp 1676037725
transform 1 0 33120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1676037725
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_373
timestamp 1676037725
transform 1 0 35420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_380
timestamp 1676037725
transform 1 0 36064 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_395
timestamp 1676037725
transform 1 0 37444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_407
timestamp 1676037725
transform 1 0 38548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_429
timestamp 1676037725
transform 1 0 40572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_441
timestamp 1676037725
transform 1 0 41676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_453
timestamp 1676037725
transform 1 0 42780 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_465
timestamp 1676037725
transform 1 0 43884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_473
timestamp 1676037725
transform 1 0 44620 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1676037725
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1676037725
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1676037725
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1676037725
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_68
timestamp 1676037725
transform 1 0 7360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1676037725
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1676037725
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1676037725
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_127
timestamp 1676037725
transform 1 0 12788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_139
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_151
timestamp 1676037725
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 1676037725
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_199
timestamp 1676037725
transform 1 0 19412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_211
timestamp 1676037725
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_234
timestamp 1676037725
transform 1 0 22632 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_246
timestamp 1676037725
transform 1 0 23736 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_258
timestamp 1676037725
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1676037725
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_285
timestamp 1676037725
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_294
timestamp 1676037725
transform 1 0 28152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_326
timestamp 1676037725
transform 1 0 31096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_333
timestamp 1676037725
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_342
timestamp 1676037725
transform 1 0 32568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_350
timestamp 1676037725
transform 1 0 33304 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_360
timestamp 1676037725
transform 1 0 34224 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_372
timestamp 1676037725
transform 1 0 35328 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_378
timestamp 1676037725
transform 1 0 35880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_409
timestamp 1676037725
transform 1 0 38732 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_424
timestamp 1676037725
transform 1 0 40112 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_446
timestamp 1676037725
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1676037725
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1676037725
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1676037725
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1676037725
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_49
timestamp 1676037725
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1676037725
transform 1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1676037725
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_110
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_149
timestamp 1676037725
transform 1 0 14812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_161
timestamp 1676037725
transform 1 0 15916 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1676037725
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_187
timestamp 1676037725
transform 1 0 18308 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1676037725
transform 1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_213
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1676037725
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_276
timestamp 1676037725
transform 1 0 26496 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_282
timestamp 1676037725
transform 1 0 27048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1676037725
transform 1 0 27416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_290
timestamp 1676037725
transform 1 0 27784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_293
timestamp 1676037725
transform 1 0 28060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1676037725
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_326
timestamp 1676037725
transform 1 0 31096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_334
timestamp 1676037725
transform 1 0 31832 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_352
timestamp 1676037725
transform 1 0 33488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_371
timestamp 1676037725
transform 1 0 35236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_388
timestamp 1676037725
transform 1 0 36800 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_408
timestamp 1676037725
transform 1 0 38640 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1676037725
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_466
timestamp 1676037725
transform 1 0 43976 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1676037725
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1676037725
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1676037725
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1676037725
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1676037725
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1676037725
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1676037725
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1676037725
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1676037725
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1676037725
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1676037725
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_18
timestamp 1676037725
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_26
timestamp 1676037725
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_38
timestamp 1676037725
transform 1 0 4600 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1676037725
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1676037725
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1676037725
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1676037725
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1676037725
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_127
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1676037725
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_202
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1676037725
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_263
timestamp 1676037725
transform 1 0 25300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1676037725
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_320
timestamp 1676037725
transform 1 0 30544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_345
timestamp 1676037725
transform 1 0 32844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_360
timestamp 1676037725
transform 1 0 34224 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_372
timestamp 1676037725
transform 1 0 35328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1676037725
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_397
timestamp 1676037725
transform 1 0 37628 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_407
timestamp 1676037725
transform 1 0 38548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_419
timestamp 1676037725
transform 1 0 39652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_427
timestamp 1676037725
transform 1 0 40388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1676037725
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_463
timestamp 1676037725
transform 1 0 43700 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1676037725
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1676037725
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1676037725
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1676037725
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1676037725
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1676037725
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1676037725
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1676037725
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1676037725
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1676037725
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_46
timestamp 1676037725
transform 1 0 5336 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1676037725
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1676037725
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_66
timestamp 1676037725
transform 1 0 7176 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1676037725
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1676037725
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_113
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_156
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_167
timestamp 1676037725
transform 1 0 16468 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1676037725
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_234
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1676037725
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_263
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_287
timestamp 1676037725
transform 1 0 27508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1676037725
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_319
timestamp 1676037725
transform 1 0 30452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_331
timestamp 1676037725
transform 1 0 31556 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_339
timestamp 1676037725
transform 1 0 32292 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1676037725
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_403
timestamp 1676037725
transform 1 0 38180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_409
timestamp 1676037725
transform 1 0 38732 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_417
timestamp 1676037725
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_453
timestamp 1676037725
transform 1 0 42780 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_461
timestamp 1676037725
transform 1 0 43516 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_472
timestamp 1676037725
transform 1 0 44528 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1676037725
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1676037725
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1676037725
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1676037725
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1676037725
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1676037725
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1676037725
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1676037725
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1676037725
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1676037725
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_19
timestamp 1676037725
transform 1 0 2852 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_34
timestamp 1676037725
transform 1 0 4232 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_40
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 1676037725
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 1676037725
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_79
timestamp 1676037725
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_100
timestamp 1676037725
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1676037725
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_183
timestamp 1676037725
transform 1 0 17940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_195
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1676037725
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1676037725
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_230
timestamp 1676037725
transform 1 0 22264 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_242
timestamp 1676037725
transform 1 0 23368 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_254
timestamp 1676037725
transform 1 0 24472 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_262
timestamp 1676037725
transform 1 0 25208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1676037725
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_299
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_315
timestamp 1676037725
transform 1 0 30084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_327
timestamp 1676037725
transform 1 0 31188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1676037725
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_411
timestamp 1676037725
transform 1 0 38916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_425
timestamp 1676037725
transform 1 0 40204 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_437
timestamp 1676037725
transform 1 0 41308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1676037725
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1676037725
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1676037725
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1676037725
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1676037725
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1676037725
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1676037725
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1676037725
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1676037725
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1676037725
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1676037725
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1676037725
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_47
timestamp 1676037725
transform 1 0 5428 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1676037725
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1676037725
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_114
timestamp 1676037725
transform 1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_123
timestamp 1676037725
transform 1 0 12420 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1676037725
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_161
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_173
timestamp 1676037725
transform 1 0 17020 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_180
timestamp 1676037725
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1676037725
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_205
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1676037725
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_216
timestamp 1676037725
transform 1 0 20976 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_261
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_267
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1676037725
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_283
timestamp 1676037725
transform 1 0 27140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1676037725
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1676037725
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_349
timestamp 1676037725
transform 1 0 33212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1676037725
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_378
timestamp 1676037725
transform 1 0 35880 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_384
timestamp 1676037725
transform 1 0 36432 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1676037725
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_406
timestamp 1676037725
transform 1 0 38456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_415
timestamp 1676037725
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_428
timestamp 1676037725
transform 1 0 40480 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_436
timestamp 1676037725
transform 1 0 41216 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_453
timestamp 1676037725
transform 1 0 42780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_465
timestamp 1676037725
transform 1 0 43884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1676037725
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1676037725
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1676037725
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1676037725
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1676037725
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1676037725
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1676037725
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1676037725
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1676037725
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1676037725
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1676037725
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_11
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_19
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_31
timestamp 1676037725
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_43
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_92
timestamp 1676037725
transform 1 0 9568 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1676037725
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1676037725
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_174
timestamp 1676037725
transform 1 0 17112 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_186
timestamp 1676037725
transform 1 0 18216 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_195
timestamp 1676037725
transform 1 0 19044 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_207
timestamp 1676037725
transform 1 0 20148 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1676037725
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_235
timestamp 1676037725
transform 1 0 22724 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_259
timestamp 1676037725
transform 1 0 24932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1676037725
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_286
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_290
timestamp 1676037725
transform 1 0 27784 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_298
timestamp 1676037725
transform 1 0 28520 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_308
timestamp 1676037725
transform 1 0 29440 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_320
timestamp 1676037725
transform 1 0 30544 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_328
timestamp 1676037725
transform 1 0 31280 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_343
timestamp 1676037725
transform 1 0 32660 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_353
timestamp 1676037725
transform 1 0 33580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_365
timestamp 1676037725
transform 1 0 34684 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_371
timestamp 1676037725
transform 1 0 35236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1676037725
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_404
timestamp 1676037725
transform 1 0 38272 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_416
timestamp 1676037725
transform 1 0 39376 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_428
timestamp 1676037725
transform 1 0 40480 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_433
timestamp 1676037725
transform 1 0 40940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_445
timestamp 1676037725
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1676037725
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1676037725
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1676037725
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1676037725
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1676037725
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1676037725
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1676037725
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1676037725
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1676037725
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1676037725
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1676037725
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1676037725
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_35
timestamp 1676037725
transform 1 0 4324 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_43
timestamp 1676037725
transform 1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_49
timestamp 1676037725
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_69
timestamp 1676037725
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_96
timestamp 1676037725
transform 1 0 9936 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_108
timestamp 1676037725
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_125
timestamp 1676037725
transform 1 0 12604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1676037725
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1676037725
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_277
timestamp 1676037725
transform 1 0 26588 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1676037725
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1676037725
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_319
timestamp 1676037725
transform 1 0 30452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_326
timestamp 1676037725
transform 1 0 31096 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_339
timestamp 1676037725
transform 1 0 32292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_351
timestamp 1676037725
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_373
timestamp 1676037725
transform 1 0 35420 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_383
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_399
timestamp 1676037725
transform 1 0 37812 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_411
timestamp 1676037725
transform 1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_456
timestamp 1676037725
transform 1 0 43056 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_468
timestamp 1676037725
transform 1 0 44160 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1676037725
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1676037725
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1676037725
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1676037725
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1676037725
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1676037725
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1676037725
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1676037725
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1676037725
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1676037725
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_22
timestamp 1676037725
transform 1 0 3128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1676037725
transform 1 0 3864 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_91
timestamp 1676037725
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1676037725
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1676037725
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1676037725
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1676037725
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_233
timestamp 1676037725
transform 1 0 22540 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_252
timestamp 1676037725
transform 1 0 24288 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1676037725
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_323
timestamp 1676037725
transform 1 0 30820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_345
timestamp 1676037725
transform 1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_357
timestamp 1676037725
transform 1 0 33948 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_369
timestamp 1676037725
transform 1 0 35052 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_381
timestamp 1676037725
transform 1 0 36156 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_389
timestamp 1676037725
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_402
timestamp 1676037725
transform 1 0 38088 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_413
timestamp 1676037725
transform 1 0 39100 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_436
timestamp 1676037725
transform 1 0 41216 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1676037725
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1676037725
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1676037725
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1676037725
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1676037725
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1676037725
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1676037725
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1676037725
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1676037725
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1676037725
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1676037725
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1676037725
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_50
timestamp 1676037725
transform 1 0 5704 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_62
timestamp 1676037725
transform 1 0 6808 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1676037725
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_117
timestamp 1676037725
transform 1 0 11868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_161
timestamp 1676037725
transform 1 0 15916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1676037725
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1676037725
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_273
timestamp 1676037725
transform 1 0 26220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_281
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_296
timestamp 1676037725
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_317
timestamp 1676037725
transform 1 0 30268 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_329
timestamp 1676037725
transform 1 0 31372 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_341
timestamp 1676037725
transform 1 0 32476 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1676037725
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1676037725
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_388
timestamp 1676037725
transform 1 0 36800 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_400
timestamp 1676037725
transform 1 0 37904 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_412
timestamp 1676037725
transform 1 0 39008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_428
timestamp 1676037725
transform 1 0 40480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_434
timestamp 1676037725
transform 1 0 41032 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_438
timestamp 1676037725
transform 1 0 41400 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_450
timestamp 1676037725
transform 1 0 42504 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_462
timestamp 1676037725
transform 1 0 43608 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1676037725
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1676037725
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1676037725
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1676037725
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1676037725
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1676037725
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1676037725
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1676037725
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1676037725
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1676037725
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1676037725
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_9
timestamp 1676037725
transform 1 0 1932 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1676037725
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1676037725
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1676037725
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_90
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_206
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1676037725
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_294
timestamp 1676037725
transform 1 0 28152 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_306
timestamp 1676037725
transform 1 0 29256 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_318
timestamp 1676037725
transform 1 0 30360 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_324
timestamp 1676037725
transform 1 0 30912 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1676037725
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_355
timestamp 1676037725
transform 1 0 33764 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_367
timestamp 1676037725
transform 1 0 34868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_375
timestamp 1676037725
transform 1 0 35604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1676037725
transform 1 0 36064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1676037725
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_411
timestamp 1676037725
transform 1 0 38916 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_423
timestamp 1676037725
transform 1 0 40020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1676037725
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_457
timestamp 1676037725
transform 1 0 43148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_472
timestamp 1676037725
transform 1 0 44528 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_483
timestamp 1676037725
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_495
timestamp 1676037725
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1676037725
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1676037725
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1676037725
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1676037725
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1676037725
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1676037725
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1676037725
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1676037725
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1676037725
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1676037725
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1676037725
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_11
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1676037725
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_151
timestamp 1676037725
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_163
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_175
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_211
timestamp 1676037725
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_236
timestamp 1676037725
transform 1 0 22816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1676037725
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_273
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_285
timestamp 1676037725
transform 1 0 27324 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_290
timestamp 1676037725
transform 1 0 27784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1676037725
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_318
timestamp 1676037725
transform 1 0 30360 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_330
timestamp 1676037725
transform 1 0 31464 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_342
timestamp 1676037725
transform 1 0 32568 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_348
timestamp 1676037725
transform 1 0 33120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_392
timestamp 1676037725
transform 1 0 37168 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_404
timestamp 1676037725
transform 1 0 38272 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1676037725
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_451
timestamp 1676037725
transform 1 0 42596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_463
timestamp 1676037725
transform 1 0 43700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1676037725
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1676037725
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1676037725
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1676037725
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1676037725
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1676037725
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1676037725
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1676037725
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1676037725
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1676037725
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1676037725
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_29
timestamp 1676037725
transform 1 0 3772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_41
timestamp 1676037725
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_65
timestamp 1676037725
transform 1 0 7084 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_87
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_99
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_183
timestamp 1676037725
transform 1 0 17940 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_257
timestamp 1676037725
transform 1 0 24748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_323
timestamp 1676037725
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_355
timestamp 1676037725
transform 1 0 33764 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_364
timestamp 1676037725
transform 1 0 34592 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_376
timestamp 1676037725
transform 1 0 35696 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_384
timestamp 1676037725
transform 1 0 36432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_400
timestamp 1676037725
transform 1 0 37904 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_412
timestamp 1676037725
transform 1 0 39008 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_420
timestamp 1676037725
transform 1 0 39744 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_470
timestamp 1676037725
transform 1 0 44344 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_482
timestamp 1676037725
transform 1 0 45448 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_490
timestamp 1676037725
transform 1 0 46184 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_502
timestamp 1676037725
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1676037725
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1676037725
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1676037725
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1676037725
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1676037725
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1676037725
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1676037725
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1676037725
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1676037725
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1676037725
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1676037725
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_35
timestamp 1676037725
transform 1 0 4324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 1676037725
transform 1 0 6348 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1676037725
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_99
timestamp 1676037725
transform 1 0 10212 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_111
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_123
timestamp 1676037725
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1676037725
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_181
timestamp 1676037725
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1676037725
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1676037725
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_293
timestamp 1676037725
transform 1 0 28060 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1676037725
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_328
timestamp 1676037725
transform 1 0 31280 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_340
timestamp 1676037725
transform 1 0 32384 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_352
timestamp 1676037725
transform 1 0 33488 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_372
timestamp 1676037725
transform 1 0 35328 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_384
timestamp 1676037725
transform 1 0 36432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_402
timestamp 1676037725
transform 1 0 38088 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_414
timestamp 1676037725
transform 1 0 39192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_425
timestamp 1676037725
transform 1 0 40204 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_442
timestamp 1676037725
transform 1 0 41768 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_462
timestamp 1676037725
transform 1 0 43608 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1676037725
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_485
timestamp 1676037725
transform 1 0 45724 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_495
timestamp 1676037725
transform 1 0 46644 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_510
timestamp 1676037725
transform 1 0 48024 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_522
timestamp 1676037725
transform 1 0 49128 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_530
timestamp 1676037725
transform 1 0 49864 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1676037725
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1676037725
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1676037725
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1676037725
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1676037725
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1676037725
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1676037725
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1676037725
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1676037725
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_18
timestamp 1676037725
transform 1 0 2760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_34
timestamp 1676037725
transform 1 0 4232 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_43
timestamp 1676037725
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_91
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1676037725
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_121
timestamp 1676037725
transform 1 0 12236 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_157
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_200
timestamp 1676037725
transform 1 0 19504 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_212
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_251
timestamp 1676037725
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_262
timestamp 1676037725
transform 1 0 25208 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1676037725
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_299
timestamp 1676037725
transform 1 0 28612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_305
timestamp 1676037725
transform 1 0 29164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1676037725
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_321
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1676037725
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_352
timestamp 1676037725
transform 1 0 33488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_364
timestamp 1676037725
transform 1 0 34592 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_374
timestamp 1676037725
transform 1 0 35512 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1676037725
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_402
timestamp 1676037725
transform 1 0 38088 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_414
timestamp 1676037725
transform 1 0 39192 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_426
timestamp 1676037725
transform 1 0 40296 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_438
timestamp 1676037725
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1676037725
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_472
timestamp 1676037725
transform 1 0 44528 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_480
timestamp 1676037725
transform 1 0 45264 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_489
timestamp 1676037725
transform 1 0 46092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_499
timestamp 1676037725
transform 1 0 47012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1676037725
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1676037725
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1676037725
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1676037725
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1676037725
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1676037725
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1676037725
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1676037725
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1676037725
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1676037725
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1676037725
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_11
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_48
timestamp 1676037725
transform 1 0 5520 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_60
timestamp 1676037725
transform 1 0 6624 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_149
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_205
timestamp 1676037725
transform 1 0 19964 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_217
timestamp 1676037725
transform 1 0 21068 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_229
timestamp 1676037725
transform 1 0 22172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1676037725
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1676037725
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1676037725
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_329
timestamp 1676037725
transform 1 0 31372 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1676037725
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_371
timestamp 1676037725
transform 1 0 35236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_378
timestamp 1676037725
transform 1 0 35880 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_384
timestamp 1676037725
transform 1 0 36432 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_432
timestamp 1676037725
transform 1 0 40848 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_444
timestamp 1676037725
transform 1 0 41952 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_456
timestamp 1676037725
transform 1 0 43056 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_468
timestamp 1676037725
transform 1 0 44160 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1676037725
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1676037725
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1676037725
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1676037725
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1676037725
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1676037725
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1676037725
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1676037725
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1676037725
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1676037725
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1676037725
transform 1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_19
timestamp 1676037725
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1676037725
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_177
timestamp 1676037725
transform 1 0 17388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1676037725
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_203
timestamp 1676037725
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1676037725
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_252
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1676037725
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1676037725
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_317
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_343
timestamp 1676037725
transform 1 0 32660 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_355
timestamp 1676037725
transform 1 0 33764 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_367
timestamp 1676037725
transform 1 0 34868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_379
timestamp 1676037725
transform 1 0 35972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_398
timestamp 1676037725
transform 1 0 37720 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_410
timestamp 1676037725
transform 1 0 38824 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_431
timestamp 1676037725
transform 1 0 40756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_443
timestamp 1676037725
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_457
timestamp 1676037725
transform 1 0 43148 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_467
timestamp 1676037725
transform 1 0 44068 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_475
timestamp 1676037725
transform 1 0 44804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_487
timestamp 1676037725
transform 1 0 45908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_499
timestamp 1676037725
transform 1 0 47012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1676037725
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1676037725
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1676037725
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1676037725
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1676037725
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1676037725
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1676037725
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1676037725
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1676037725
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1676037725
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1676037725
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1676037725
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1676037725
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_61
timestamp 1676037725
transform 1 0 6716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_73
timestamp 1676037725
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1676037725
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_99
timestamp 1676037725
transform 1 0 10212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_111
timestamp 1676037725
transform 1 0 11316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1676037725
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_206
timestamp 1676037725
transform 1 0 20056 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_214
timestamp 1676037725
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_225
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_240
timestamp 1676037725
transform 1 0 23184 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_273
timestamp 1676037725
transform 1 0 26220 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_282
timestamp 1676037725
transform 1 0 27048 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_294
timestamp 1676037725
transform 1 0 28152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1676037725
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_325
timestamp 1676037725
transform 1 0 31004 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_337
timestamp 1676037725
transform 1 0 32108 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_349
timestamp 1676037725
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1676037725
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_394
timestamp 1676037725
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_406
timestamp 1676037725
transform 1 0 38456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1676037725
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_441
timestamp 1676037725
transform 1 0 41676 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_456
timestamp 1676037725
transform 1 0 43056 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_468
timestamp 1676037725
transform 1 0 44160 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1676037725
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_488
timestamp 1676037725
transform 1 0 46000 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_500
timestamp 1676037725
transform 1 0 47104 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_512
timestamp 1676037725
transform 1 0 48208 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_524
timestamp 1676037725
transform 1 0 49312 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1676037725
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1676037725
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1676037725
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1676037725
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1676037725
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1676037725
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1676037725
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1676037725
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1676037725
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_11
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_67
timestamp 1676037725
transform 1 0 7268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1676037725
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1676037725
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_290
timestamp 1676037725
transform 1 0 27784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_302
timestamp 1676037725
transform 1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_308
timestamp 1676037725
transform 1 0 29440 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1676037725
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_343
timestamp 1676037725
transform 1 0 32660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_355
timestamp 1676037725
transform 1 0 33764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_372
timestamp 1676037725
transform 1 0 35328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1676037725
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_403
timestamp 1676037725
transform 1 0 38180 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_415
timestamp 1676037725
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_427
timestamp 1676037725
transform 1 0 40388 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_436
timestamp 1676037725
transform 1 0 41216 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_453
timestamp 1676037725
transform 1 0 42780 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_468
timestamp 1676037725
transform 1 0 44160 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_477
timestamp 1676037725
transform 1 0 44988 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_489
timestamp 1676037725
transform 1 0 46092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_501
timestamp 1676037725
transform 1 0 47196 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1676037725
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1676037725
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1676037725
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1676037725
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1676037725
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1676037725
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1676037725
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1676037725
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1676037725
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1676037725
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1676037725
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_37
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_43
timestamp 1676037725
transform 1 0 5060 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_66
timestamp 1676037725
transform 1 0 7176 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_98
timestamp 1676037725
transform 1 0 10120 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_111
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_123
timestamp 1676037725
transform 1 0 12420 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_149
timestamp 1676037725
transform 1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1676037725
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_202
timestamp 1676037725
transform 1 0 19688 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_223
timestamp 1676037725
transform 1 0 21620 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_235
timestamp 1676037725
transform 1 0 22724 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1676037725
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_262
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_297
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_315
timestamp 1676037725
transform 1 0 30084 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_327
timestamp 1676037725
transform 1 0 31188 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_339
timestamp 1676037725
transform 1 0 32292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_351
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_394
timestamp 1676037725
transform 1 0 37352 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_406
timestamp 1676037725
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1676037725
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_437
timestamp 1676037725
transform 1 0 41308 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_441
timestamp 1676037725
transform 1 0 41676 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_453
timestamp 1676037725
transform 1 0 42780 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_465
timestamp 1676037725
transform 1 0 43884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_473
timestamp 1676037725
transform 1 0 44620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_487
timestamp 1676037725
transform 1 0 45908 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_499
timestamp 1676037725
transform 1 0 47012 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_511
timestamp 1676037725
transform 1 0 48116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_523
timestamp 1676037725
transform 1 0 49220 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1676037725
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1676037725
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1676037725
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1676037725
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1676037725
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1676037725
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1676037725
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1676037725
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1676037725
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1676037725
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_25
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_33
timestamp 1676037725
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_77
timestamp 1676037725
transform 1 0 8188 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_94
timestamp 1676037725
transform 1 0 9752 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_211
timestamp 1676037725
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1676037725
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1676037725
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_290
timestamp 1676037725
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_298
timestamp 1676037725
transform 1 0 28520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_326
timestamp 1676037725
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_353
timestamp 1676037725
transform 1 0 33580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_363
timestamp 1676037725
transform 1 0 34500 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_372
timestamp 1676037725
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1676037725
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_411
timestamp 1676037725
transform 1 0 38916 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_423
timestamp 1676037725
transform 1 0 40020 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1676037725
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1676037725
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1676037725
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1676037725
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1676037725
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1676037725
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1676037725
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1676037725
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1676037725
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1676037725
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1676037725
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1676037725
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_18
timestamp 1676037725
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_73
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1676037725
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1676037725
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_102
timestamp 1676037725
transform 1 0 10488 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1676037725
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_164
timestamp 1676037725
transform 1 0 16192 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_176
timestamp 1676037725
transform 1 0 17296 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_215
timestamp 1676037725
transform 1 0 20884 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_225
timestamp 1676037725
transform 1 0 21804 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_235
timestamp 1676037725
transform 1 0 22724 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_275
timestamp 1676037725
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_286
timestamp 1676037725
transform 1 0 27416 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_298
timestamp 1676037725
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1676037725
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_315
timestamp 1676037725
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_322
timestamp 1676037725
transform 1 0 30728 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_331
timestamp 1676037725
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_343
timestamp 1676037725
transform 1 0 32660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_370
timestamp 1676037725
transform 1 0 35144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_382
timestamp 1676037725
transform 1 0 36248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1676037725
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_412
timestamp 1676037725
transform 1 0 39008 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_450
timestamp 1676037725
transform 1 0 42504 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_462
timestamp 1676037725
transform 1 0 43608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_470
timestamp 1676037725
transform 1 0 44344 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1676037725
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_487
timestamp 1676037725
transform 1 0 45908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_499
timestamp 1676037725
transform 1 0 47012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_511
timestamp 1676037725
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_523
timestamp 1676037725
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1676037725
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1676037725
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1676037725
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1676037725
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1676037725
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1676037725
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1676037725
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1676037725
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1676037725
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1676037725
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_11
timestamp 1676037725
transform 1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_33
timestamp 1676037725
transform 1 0 4140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1676037725
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_67
timestamp 1676037725
transform 1 0 7268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_79
timestamp 1676037725
transform 1 0 8372 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_144
timestamp 1676037725
transform 1 0 14352 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_156
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_182
timestamp 1676037725
transform 1 0 17848 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_201
timestamp 1676037725
transform 1 0 19596 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_213
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_233
timestamp 1676037725
transform 1 0 22540 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_245
timestamp 1676037725
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_257
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_290
timestamp 1676037725
transform 1 0 27784 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1676037725
transform 1 0 28520 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_315
timestamp 1676037725
transform 1 0 30084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1676037725
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_356
timestamp 1676037725
transform 1 0 33856 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_363
timestamp 1676037725
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_375
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1676037725
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_400
timestamp 1676037725
transform 1 0 37904 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_404
timestamp 1676037725
transform 1 0 38272 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_416
timestamp 1676037725
transform 1 0 39376 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_428
timestamp 1676037725
transform 1 0 40480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_435
timestamp 1676037725
transform 1 0 41124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1676037725
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1676037725
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1676037725
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1676037725
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1676037725
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1676037725
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1676037725
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1676037725
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1676037725
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1676037725
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1676037725
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1676037725
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1676037725
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_35
timestamp 1676037725
transform 1 0 4324 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_59
timestamp 1676037725
transform 1 0 6532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_71
timestamp 1676037725
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1676037725
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_101
timestamp 1676037725
transform 1 0 10396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1676037725
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_149
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_161
timestamp 1676037725
transform 1 0 15916 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_185
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_208
timestamp 1676037725
transform 1 0 20240 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_220
timestamp 1676037725
transform 1 0 21344 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_238
timestamp 1676037725
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1676037725
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_267
timestamp 1676037725
transform 1 0 25668 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_279
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_291
timestamp 1676037725
transform 1 0 27876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1676037725
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_317
timestamp 1676037725
transform 1 0 30268 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1676037725
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_338
timestamp 1676037725
transform 1 0 32200 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_373
timestamp 1676037725
transform 1 0 35420 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_404
timestamp 1676037725
transform 1 0 38272 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1676037725
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_441
timestamp 1676037725
transform 1 0 41676 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_453
timestamp 1676037725
transform 1 0 42780 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_465
timestamp 1676037725
transform 1 0 43884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_473
timestamp 1676037725
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1676037725
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1676037725
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1676037725
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1676037725
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1676037725
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1676037725
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1676037725
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1676037725
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1676037725
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1676037725
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_18
timestamp 1676037725
transform 1 0 2760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_26
timestamp 1676037725
transform 1 0 3496 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1676037725
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_80
timestamp 1676037725
transform 1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1676037725
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1676037725
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_133
timestamp 1676037725
transform 1 0 13340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1676037725
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_177
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_189
timestamp 1676037725
transform 1 0 18492 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_194
timestamp 1676037725
transform 1 0 18952 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_206
timestamp 1676037725
transform 1 0 20056 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1676037725
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_256
timestamp 1676037725
transform 1 0 24656 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1676037725
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_310
timestamp 1676037725
transform 1 0 29624 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_322
timestamp 1676037725
transform 1 0 30728 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1676037725
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1676037725
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1676037725
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1676037725
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1676037725
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1676037725
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1676037725
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1676037725
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1676037725
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1676037725
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1676037725
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1676037725
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1676037725
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1676037725
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1676037725
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_19
timestamp 1676037725
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_45
timestamp 1676037725
transform 1 0 5244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1676037725
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_117
timestamp 1676037725
transform 1 0 11868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1676037725
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_175
timestamp 1676037725
transform 1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_179
timestamp 1676037725
transform 1 0 17572 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_184
timestamp 1676037725
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_217
timestamp 1676037725
transform 1 0 21068 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_274
timestamp 1676037725
transform 1 0 26312 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_286
timestamp 1676037725
transform 1 0 27416 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_292
timestamp 1676037725
transform 1 0 27968 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_318
timestamp 1676037725
transform 1 0 30360 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_330
timestamp 1676037725
transform 1 0 31464 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_342
timestamp 1676037725
transform 1 0 32568 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_348
timestamp 1676037725
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1676037725
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_412
timestamp 1676037725
transform 1 0 39008 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_429
timestamp 1676037725
transform 1 0 40572 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_448
timestamp 1676037725
transform 1 0 42320 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_460
timestamp 1676037725
transform 1 0 43424 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1676037725
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1676037725
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1676037725
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1676037725
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1676037725
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1676037725
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1676037725
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1676037725
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1676037725
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1676037725
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1676037725
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1676037725
transform 1 0 2116 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_24
timestamp 1676037725
transform 1 0 3312 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_36
timestamp 1676037725
transform 1 0 4416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_40
timestamp 1676037725
transform 1 0 4784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1676037725
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_75
timestamp 1676037725
transform 1 0 8004 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_87
timestamp 1676037725
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_99
timestamp 1676037725
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_177
timestamp 1676037725
transform 1 0 17388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_189
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_201
timestamp 1676037725
transform 1 0 19596 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_269
timestamp 1676037725
transform 1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1676037725
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_318
timestamp 1676037725
transform 1 0 30360 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_326
timestamp 1676037725
transform 1 0 31096 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_342
timestamp 1676037725
transform 1 0 32568 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_355
timestamp 1676037725
transform 1 0 33764 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_367
timestamp 1676037725
transform 1 0 34868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_379
timestamp 1676037725
transform 1 0 35972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_425
timestamp 1676037725
transform 1 0 40204 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1676037725
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1676037725
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1676037725
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1676037725
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1676037725
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1676037725
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1676037725
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1676037725
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1676037725
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1676037725
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1676037725
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_115
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_127
timestamp 1676037725
transform 1 0 12788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_164
timestamp 1676037725
transform 1 0 16192 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_176
timestamp 1676037725
transform 1 0 17296 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1676037725
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_206
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_218
timestamp 1676037725
transform 1 0 21160 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_236
timestamp 1676037725
transform 1 0 22816 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_263
timestamp 1676037725
transform 1 0 25300 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_271
timestamp 1676037725
transform 1 0 26036 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_341
timestamp 1676037725
transform 1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_384
timestamp 1676037725
transform 1 0 36432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_406
timestamp 1676037725
transform 1 0 38456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1676037725
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_461
timestamp 1676037725
transform 1 0 43516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 1676037725
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1676037725
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1676037725
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1676037725
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1676037725
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1676037725
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1676037725
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1676037725
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1676037725
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1676037725
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1676037725
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1676037725
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_19
timestamp 1676037725
transform 1 0 2852 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1676037725
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1676037725
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_191
timestamp 1676037725
transform 1 0 18676 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_208
timestamp 1676037725
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1676037725
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_268
timestamp 1676037725
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_304
timestamp 1676037725
transform 1 0 29072 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_310
timestamp 1676037725
transform 1 0 29624 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_319
timestamp 1676037725
transform 1 0 30452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1676037725
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_343
timestamp 1676037725
transform 1 0 32660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_355
timestamp 1676037725
transform 1 0 33764 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_359
timestamp 1676037725
transform 1 0 34132 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_365
timestamp 1676037725
transform 1 0 34684 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_377
timestamp 1676037725
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1676037725
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_401
timestamp 1676037725
transform 1 0 37996 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_410
timestamp 1676037725
transform 1 0 38824 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_422
timestamp 1676037725
transform 1 0 39928 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_428
timestamp 1676037725
transform 1 0 40480 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1676037725
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1676037725
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1676037725
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1676037725
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1676037725
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1676037725
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1676037725
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1676037725
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1676037725
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1676037725
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1676037725
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1676037725
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1676037725
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_9
timestamp 1676037725
transform 1 0 1932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_45
timestamp 1676037725
transform 1 0 5244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_62
timestamp 1676037725
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1676037725
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_159
timestamp 1676037725
transform 1 0 15732 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_171
timestamp 1676037725
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_183
timestamp 1676037725
transform 1 0 17940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_202
timestamp 1676037725
transform 1 0 19688 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_214
timestamp 1676037725
transform 1 0 20792 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_231
timestamp 1676037725
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1676037725
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_272
timestamp 1676037725
transform 1 0 26128 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_284
timestamp 1676037725
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_296
timestamp 1676037725
transform 1 0 28336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_330
timestamp 1676037725
transform 1 0 31464 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_342
timestamp 1676037725
transform 1 0 32568 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1676037725
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1676037725
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1676037725
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_402
timestamp 1676037725
transform 1 0 38088 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_414
timestamp 1676037725
transform 1 0 39192 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1676037725
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1676037725
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1676037725
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1676037725
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1676037725
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1676037725
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1676037725
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1676037725
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1676037725
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1676037725
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1676037725
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1676037725
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1676037725
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_11
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_19
timestamp 1676037725
transform 1 0 2852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_38
timestamp 1676037725
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1676037725
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_79
timestamp 1676037725
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_91
timestamp 1676037725
transform 1 0 9476 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1676037725
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_153
timestamp 1676037725
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_188
timestamp 1676037725
transform 1 0 18400 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_200
timestamp 1676037725
transform 1 0 19504 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_212
timestamp 1676037725
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_305
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_309
timestamp 1676037725
transform 1 0 29532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_344
timestamp 1676037725
transform 1 0 32752 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_352
timestamp 1676037725
transform 1 0 33488 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_359
timestamp 1676037725
transform 1 0 34132 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_367
timestamp 1676037725
transform 1 0 34868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_371
timestamp 1676037725
transform 1 0 35236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1676037725
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1676037725
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_417
timestamp 1676037725
transform 1 0 39468 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_425
timestamp 1676037725
transform 1 0 40204 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_433
timestamp 1676037725
transform 1 0 40940 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_440
timestamp 1676037725
transform 1 0 41584 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_454
timestamp 1676037725
transform 1 0 42872 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_466
timestamp 1676037725
transform 1 0 43976 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_478
timestamp 1676037725
transform 1 0 45080 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_490
timestamp 1676037725
transform 1 0 46184 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_502
timestamp 1676037725
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1676037725
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1676037725
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1676037725
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1676037725
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1676037725
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1676037725
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1676037725
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1676037725
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1676037725
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1676037725
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1676037725
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1676037725
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1676037725
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_62
timestamp 1676037725
transform 1 0 6808 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_68
timestamp 1676037725
transform 1 0 7360 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp 1676037725
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1676037725
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1676037725
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_163
timestamp 1676037725
transform 1 0 16100 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1676037725
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_205
timestamp 1676037725
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_214
timestamp 1676037725
transform 1 0 20792 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_223
timestamp 1676037725
transform 1 0 21620 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_231
timestamp 1676037725
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_259
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_271
timestamp 1676037725
transform 1 0 26036 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_283
timestamp 1676037725
transform 1 0 27140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_295
timestamp 1676037725
transform 1 0 28244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_327
timestamp 1676037725
transform 1 0 31188 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_344
timestamp 1676037725
transform 1 0 32752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_354
timestamp 1676037725
transform 1 0 33672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_358
timestamp 1676037725
transform 1 0 34040 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1676037725
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_373
timestamp 1676037725
transform 1 0 35420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_386
timestamp 1676037725
transform 1 0 36616 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_402
timestamp 1676037725
transform 1 0 38088 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1676037725
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_432
timestamp 1676037725
transform 1 0 40848 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_444
timestamp 1676037725
transform 1 0 41952 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_456
timestamp 1676037725
transform 1 0 43056 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_468
timestamp 1676037725
transform 1 0 44160 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1676037725
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1676037725
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1676037725
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1676037725
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1676037725
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1676037725
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1676037725
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1676037725
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1676037725
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1676037725
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1676037725
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1676037725
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_19
timestamp 1676037725
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_31
timestamp 1676037725
transform 1 0 3956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_43
timestamp 1676037725
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_145
timestamp 1676037725
transform 1 0 14444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1676037725
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_158
timestamp 1676037725
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1676037725
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_199
timestamp 1676037725
transform 1 0 19412 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_204
timestamp 1676037725
transform 1 0 19872 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1676037725
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1676037725
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_256
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_268
timestamp 1676037725
transform 1 0 25760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_368
timestamp 1676037725
transform 1 0 34960 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_380
timestamp 1676037725
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1676037725
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1676037725
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1676037725
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1676037725
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1676037725
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1676037725
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1676037725
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1676037725
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1676037725
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1676037725
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1676037725
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_11
timestamp 1676037725
transform 1 0 2116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1676037725
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_206
timestamp 1676037725
transform 1 0 20056 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_218
timestamp 1676037725
transform 1 0 21160 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_230
timestamp 1676037725
transform 1 0 22264 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1676037725
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1676037725
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1676037725
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1676037725
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1676037725
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1676037725
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1676037725
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1676037725
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1676037725
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1676037725
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1676037725
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1676037725
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_11
timestamp 1676037725
transform 1 0 2116 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_19
timestamp 1676037725
transform 1 0 2852 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_31
timestamp 1676037725
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1676037725
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1676037725
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1676037725
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1676037725
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1676037725
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1676037725
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1676037725
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1676037725
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1676037725
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1676037725
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1676037725
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1676037725
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1676037725
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1676037725
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_11
timestamp 1676037725
transform 1 0 2116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1676037725
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1676037725
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1676037725
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1676037725
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1676037725
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1676037725
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1676037725
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1676037725
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1676037725
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1676037725
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1676037725
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1676037725
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1676037725
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1676037725
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1676037725
transform 1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_19
timestamp 1676037725
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_31
timestamp 1676037725
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_43
timestamp 1676037725
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1676037725
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1676037725
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1676037725
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1676037725
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1676037725
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1676037725
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1676037725
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1676037725
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1676037725
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1676037725
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1676037725
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1676037725
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_11
timestamp 1676037725
transform 1 0 2116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1676037725
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1676037725
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1676037725
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1676037725
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1676037725
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1676037725
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1676037725
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1676037725
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1676037725
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1676037725
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1676037725
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1676037725
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1676037725
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1676037725
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1676037725
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1676037725
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_11
timestamp 1676037725
transform 1 0 2116 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1676037725
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1676037725
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1676037725
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1676037725
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1676037725
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1676037725
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1676037725
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1676037725
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1676037725
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1676037725
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1676037725
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1676037725
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1676037725
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1676037725
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1676037725
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1676037725
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1676037725
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1676037725
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_11
timestamp 1676037725
transform 1 0 2116 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1676037725
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1676037725
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1676037725
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1676037725
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1676037725
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1676037725
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1676037725
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1676037725
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1676037725
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1676037725
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1676037725
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1676037725
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_11
timestamp 1676037725
transform 1 0 2116 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_23
timestamp 1676037725
transform 1 0 3220 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_35
timestamp 1676037725
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_47
timestamp 1676037725
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1676037725
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1676037725
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1676037725
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1676037725
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1676037725
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1676037725
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1676037725
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1676037725
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1676037725
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1676037725
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1676037725
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1676037725
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1676037725
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1676037725
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1676037725
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1676037725
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_9
timestamp 1676037725
transform 1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_17
timestamp 1676037725
transform 1 0 2668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 1676037725
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1676037725
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1676037725
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1676037725
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1676037725
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1676037725
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1676037725
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1676037725
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1676037725
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1676037725
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1676037725
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1676037725
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1676037725
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_11
timestamp 1676037725
transform 1 0 2116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_23
timestamp 1676037725
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1676037725
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1676037725
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1676037725
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1676037725
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1676037725
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1676037725
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1676037725
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1676037725
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1676037725
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1676037725
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1676037725
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1676037725
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1676037725
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1676037725
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1676037725
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1676037725
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1676037725
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1676037725
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1676037725
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1676037725
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1676037725
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1676037725
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1676037725
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1676037725
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1676037725
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1676037725
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1676037725
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1676037725
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_11
timestamp 1676037725
transform 1 0 2116 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_23
timestamp 1676037725
transform 1 0 3220 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_35
timestamp 1676037725
transform 1 0 4324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1676037725
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1676037725
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1676037725
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1676037725
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1676037725
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1676037725
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1676037725
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1676037725
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1676037725
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1676037725
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1676037725
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1676037725
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1676037725
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1676037725
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1676037725
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1676037725
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1676037725
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1676037725
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1676037725
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1676037725
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1676037725
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1676037725
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1676037725
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1676037725
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1676037725
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1676037725
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1676037725
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1676037725
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1676037725
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1676037725
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1676037725
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1676037725
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1676037725
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1676037725
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1676037725
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1676037725
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_17
timestamp 1676037725
transform 1 0 2668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_29
timestamp 1676037725
transform 1 0 3772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_41
timestamp 1676037725
transform 1 0 4876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1676037725
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1676037725
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1676037725
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1676037725
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1676037725
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1676037725
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1676037725
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1676037725
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1676037725
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1676037725
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1676037725
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1676037725
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1676037725
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_11
timestamp 1676037725
transform 1 0 2116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1676037725
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1676037725
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1676037725
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1676037725
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1676037725
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1676037725
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1676037725
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1676037725
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1676037725
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1676037725
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1676037725
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1676037725
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1676037725
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1676037725
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1676037725
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1676037725
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1676037725
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1676037725
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1676037725
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1676037725
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_11
timestamp 1676037725
transform 1 0 2116 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_23
timestamp 1676037725
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_35
timestamp 1676037725
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1676037725
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1676037725
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1676037725
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1676037725
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1676037725
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1676037725
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1676037725
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1676037725
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1676037725
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1676037725
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1676037725
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1676037725
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1676037725
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1676037725
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1676037725
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1676037725
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1676037725
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1676037725
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1676037725
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1676037725
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1676037725
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1676037725
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1676037725
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1676037725
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1676037725
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1676037725
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1676037725
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1676037725
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1676037725
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1676037725
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1676037725
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1676037725
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1676037725
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1676037725
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1676037725
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1676037725
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_11
timestamp 1676037725
transform 1 0 2116 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_23
timestamp 1676037725
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1676037725
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1676037725
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1676037725
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1676037725
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1676037725
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1676037725
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1676037725
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1676037725
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1676037725
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1676037725
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1676037725
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1676037725
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1676037725
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1676037725
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1676037725
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1676037725
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_11
timestamp 1676037725
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1676037725
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1676037725
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1676037725
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1676037725
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1676037725
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1676037725
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1676037725
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1676037725
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1676037725
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1676037725
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1676037725
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1676037725
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1676037725
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1676037725
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1676037725
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1676037725
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1676037725
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1676037725
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1676037725
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1676037725
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1676037725
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1676037725
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1676037725
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1676037725
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1676037725
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1676037725
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_11
timestamp 1676037725
transform 1 0 2116 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_23
timestamp 1676037725
transform 1 0 3220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1676037725
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1676037725
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1676037725
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1676037725
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1676037725
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1676037725
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1676037725
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1676037725
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1676037725
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1676037725
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_11
timestamp 1676037725
transform 1 0 2116 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1676037725
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1676037725
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1676037725
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1676037725
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1676037725
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1676037725
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1676037725
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1676037725
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1676037725
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1676037725
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1676037725
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1676037725
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1676037725
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1676037725
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1676037725
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1676037725
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1676037725
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1676037725
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1676037725
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1676037725
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_11
timestamp 1676037725
transform 1 0 2116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_37
timestamp 1676037725
transform 1 0 4508 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_49
timestamp 1676037725
transform 1 0 5612 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_55
timestamp 1676037725
transform 1 0 6164 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_57
timestamp 1676037725
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_69
timestamp 1676037725
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1676037725
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_113
timestamp 1676037725
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_125
timestamp 1676037725
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1676037725
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_169
timestamp 1676037725
transform 1 0 16652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_181
timestamp 1676037725
transform 1 0 17756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1676037725
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_202
timestamp 1676037725
transform 1 0 19688 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_214
timestamp 1676037725
transform 1 0 20792 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_222
timestamp 1676037725
transform 1 0 21528 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_225
timestamp 1676037725
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_237
timestamp 1676037725
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1676037725
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_281
timestamp 1676037725
transform 1 0 26956 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_337
timestamp 1676037725
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_349
timestamp 1676037725
transform 1 0 33212 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_359
timestamp 1676037725
transform 1 0 34132 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_393
timestamp 1676037725
transform 1 0 37260 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_405
timestamp 1676037725
transform 1 0 38364 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_417
timestamp 1676037725
transform 1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_439
timestamp 1676037725
transform 1 0 41492 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_447
timestamp 1676037725
transform 1 0 42228 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_449
timestamp 1676037725
transform 1 0 42412 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_461
timestamp 1676037725
transform 1 0 43516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1676037725
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_505
timestamp 1676037725
transform 1 0 47564 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_520
timestamp 1676037725
transform 1 0 48944 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1676037725
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1676037725
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_557
timestamp 1676037725
transform 1 0 52348 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_561
timestamp 1676037725
transform 1 0 52716 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_573
timestamp 1676037725
transform 1 0 53820 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_585
timestamp 1676037725
transform 1 0 54924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_589
timestamp 1676037725
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_597
timestamp 1676037725
transform 1 0 56028 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_604
timestamp 1676037725
transform 1 0 56672 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_617
timestamp 1676037725
transform 1 0 57868 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  Flash_238 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_239
timestamp 1676037725
transform 1 0 48668 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_240
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_241
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_242
timestamp 1676037725
transform 1 0 19412 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_243
timestamp 1676037725
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_244
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_245
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_246
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 42320 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 47472 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 52624 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 57776 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1676037725
transform 1 0 42596 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1676037725
transform 1 0 34132 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1676037725
transform 1 0 19320 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1676037725
transform 1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1676037725
transform 1 0 20976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1676037725
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1676037725
transform 1 0 21160 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0493_
timestamp 1676037725
transform 1 0 4876 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31280 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0498_
timestamp 1676037725
transform 1 0 5428 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0499_
timestamp 1676037725
transform 1 0 10212 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0500_
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0501_
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0502_
timestamp 1676037725
transform 1 0 12144 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0503_
timestamp 1676037725
transform 1 0 5428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0504_
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1676037725
transform 1 0 16928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30176 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0508_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0511_
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _0512_
timestamp 1676037725
transform 1 0 8740 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _0513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0514_
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0516_
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0517_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _0518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0519_
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0520_
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0522_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0523_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0524_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0525_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0527_
timestamp 1676037725
transform 1 0 14720 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0529_
timestamp 1676037725
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0531_
timestamp 1676037725
transform 1 0 14628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0532_
timestamp 1676037725
transform 1 0 15364 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0533_
timestamp 1676037725
transform 1 0 20240 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0534_
timestamp 1676037725
transform 1 0 19504 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0535_
timestamp 1676037725
transform 1 0 19780 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0536_
timestamp 1676037725
transform 1 0 24288 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0537_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0539_
timestamp 1676037725
transform 1 0 20148 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0540_
timestamp 1676037725
transform 1 0 21160 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0541_
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0542_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0543_
timestamp 1676037725
transform 1 0 18400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0545_
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0546_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0547_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0548_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0550_
timestamp 1676037725
transform 1 0 13892 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0551_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0553_
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0554_
timestamp 1676037725
transform 1 0 11960 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0555_
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0556_
timestamp 1676037725
transform 1 0 9844 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0557_
timestamp 1676037725
transform 1 0 26036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0558_
timestamp 1676037725
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0560_
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0561_
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0562_
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0563_
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0564_
timestamp 1676037725
transform 1 0 12696 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0565_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0566_
timestamp 1676037725
transform 1 0 9384 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0567_
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0568_
timestamp 1676037725
transform 1 0 28244 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0569_
timestamp 1676037725
transform 1 0 24748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0570_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0571_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0572_
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0573_
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0574_
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0575_
timestamp 1676037725
transform 1 0 11868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0576_
timestamp 1676037725
transform 1 0 29256 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0577_
timestamp 1676037725
transform 1 0 27324 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0578_
timestamp 1676037725
transform 1 0 36524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0579_
timestamp 1676037725
transform 1 0 33856 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0580_
timestamp 1676037725
transform 1 0 35604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0581_
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0582_
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0583_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0584_
timestamp 1676037725
transform 1 0 32384 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0585_
timestamp 1676037725
transform 1 0 31372 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0586_
timestamp 1676037725
transform 1 0 29164 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0587_
timestamp 1676037725
transform 1 0 37720 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0588_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0589_
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0590_
timestamp 1676037725
transform 1 0 20976 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0591_
timestamp 1676037725
transform 1 0 28704 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0592_
timestamp 1676037725
transform 1 0 10488 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0593_
timestamp 1676037725
transform 1 0 23460 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0594_
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0595_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0596_
timestamp 1676037725
transform 1 0 34960 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0597_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0598_
timestamp 1676037725
transform 1 0 31280 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1676037725
transform 1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _0601_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35696 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_4  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0605_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0606_
timestamp 1676037725
transform 1 0 31556 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0607_
timestamp 1676037725
transform 1 0 34868 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 1676037725
transform 1 0 33948 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0609_
timestamp 1676037725
transform 1 0 33856 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0610_
timestamp 1676037725
transform 1 0 33396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0611_
timestamp 1676037725
transform 1 0 36248 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35144 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0613_
timestamp 1676037725
transform 1 0 34868 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0614_
timestamp 1676037725
transform 1 0 35420 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0615_
timestamp 1676037725
transform 1 0 43884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0616_
timestamp 1676037725
transform 1 0 43700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0617_
timestamp 1676037725
transform 1 0 42596 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0618_
timestamp 1676037725
transform 1 0 42596 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 44804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 1676037725
transform 1 0 40020 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1676037725
transform 1 0 43608 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0623_
timestamp 1676037725
transform 1 0 41124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40020 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0625_
timestamp 1676037725
transform 1 0 37628 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0626_
timestamp 1676037725
transform 1 0 40020 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0627_
timestamp 1676037725
transform 1 0 39284 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0628_
timestamp 1676037725
transform 1 0 40848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1676037725
transform 1 0 45172 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0630_
timestamp 1676037725
transform 1 0 42596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1676037725
transform 1 0 43976 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0632_
timestamp 1676037725
transform 1 0 41400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1676037725
transform 1 0 38732 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0634_
timestamp 1676037725
transform 1 0 37628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1676037725
transform 1 0 35880 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0636_
timestamp 1676037725
transform 1 0 33212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0638_
timestamp 1676037725
transform 1 0 36248 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0639_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0640_
timestamp 1676037725
transform 1 0 38824 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0641_
timestamp 1676037725
transform 1 0 39008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1676037725
transform 1 0 39836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0644_
timestamp 1676037725
transform 1 0 38640 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0645_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1676037725
transform 1 0 43700 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0647_
timestamp 1676037725
transform 1 0 42964 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0648_
timestamp 1676037725
transform 1 0 38824 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0649_
timestamp 1676037725
transform 1 0 38548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 1676037725
transform 1 0 40664 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0651_
timestamp 1676037725
transform 1 0 39560 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0652_
timestamp 1676037725
transform 1 0 40112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0653_
timestamp 1676037725
transform 1 0 41124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0654_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0655_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1676037725
transform 1 0 38640 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0657_
timestamp 1676037725
transform 1 0 36524 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0658_
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0659_
timestamp 1676037725
transform 1 0 35420 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0660_
timestamp 1676037725
transform 1 0 32752 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0661_
timestamp 1676037725
transform 1 0 31648 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0662_
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0663_
timestamp 1676037725
transform 1 0 29808 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0664_
timestamp 1676037725
transform 1 0 29716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1676037725
transform 1 0 31464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0666_
timestamp 1676037725
transform 1 0 29900 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0667_
timestamp 1676037725
transform 1 0 32568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1676037725
transform 1 0 33948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1676037725
transform 1 0 37720 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0670_
timestamp 1676037725
transform 1 0 37444 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0671_
timestamp 1676037725
transform 1 0 33396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0672_
timestamp 1676037725
transform 1 0 30912 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0673_
timestamp 1676037725
transform 1 0 33856 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0675_
timestamp 1676037725
transform 1 0 32292 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0676_
timestamp 1676037725
transform 1 0 30912 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0678_
timestamp 1676037725
transform 1 0 29900 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0679_
timestamp 1676037725
transform 1 0 29716 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1676037725
transform 1 0 32844 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0683_
timestamp 1676037725
transform 1 0 31464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0684_
timestamp 1676037725
transform 1 0 30728 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0685_
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0686_
timestamp 1676037725
transform 1 0 35052 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0687_
timestamp 1676037725
transform 1 0 30544 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0688_
timestamp 1676037725
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0689_
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0690_
timestamp 1676037725
transform 1 0 29256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1676037725
transform 1 0 32384 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0693_
timestamp 1676037725
transform 1 0 29900 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0694_
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0695_
timestamp 1676037725
transform 1 0 33304 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1676037725
transform 1 0 33672 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0697_
timestamp 1676037725
transform 1 0 34224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0698_
timestamp 1676037725
transform 1 0 28060 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0699_
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0700_
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0701_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0702_
timestamp 1676037725
transform 1 0 37720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_2  _0703_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38456 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0704_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33120 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0705_
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0706_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0707_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0708_
timestamp 1676037725
transform 1 0 32292 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29624 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0711_
timestamp 1676037725
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0712_
timestamp 1676037725
transform 1 0 28336 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0713_
timestamp 1676037725
transform 1 0 25852 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0714_
timestamp 1676037725
transform 1 0 26128 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0715_
timestamp 1676037725
transform 1 0 34960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33580 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0717_
timestamp 1676037725
transform 1 0 35972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0718_
timestamp 1676037725
transform 1 0 36156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0719_
timestamp 1676037725
transform 1 0 34224 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0720_
timestamp 1676037725
transform 1 0 34408 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0721_
timestamp 1676037725
transform 1 0 34868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0722_
timestamp 1676037725
transform 1 0 37536 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35880 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0724_
timestamp 1676037725
transform 1 0 36524 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0725_
timestamp 1676037725
transform 1 0 40020 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0726_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38088 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0727_
timestamp 1676037725
transform 1 0 39836 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0728_
timestamp 1676037725
transform 1 0 38824 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41032 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0730_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0731_
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0732_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0733_
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0734_
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0737_
timestamp 1676037725
transform 1 0 18400 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0738_
timestamp 1676037725
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0739_
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0740_
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0741_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0742_
timestamp 1676037725
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0743_
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0744_
timestamp 1676037725
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0745_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1676037725
transform 1 0 17848 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0748_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0749_
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0750_
timestamp 1676037725
transform 1 0 23552 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0751_
timestamp 1676037725
transform 1 0 21896 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0752_
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0753_
timestamp 1676037725
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0754_
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _0756_
timestamp 1676037725
transform 1 0 23736 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0758_
timestamp 1676037725
transform 1 0 22724 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0759_
timestamp 1676037725
transform 1 0 27140 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1676037725
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 1676037725
transform 1 0 27508 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0763_
timestamp 1676037725
transform 1 0 27140 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0764_
timestamp 1676037725
transform 1 0 26496 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0765_
timestamp 1676037725
transform 1 0 25760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0766_
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0767_
timestamp 1676037725
transform 1 0 25668 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0768_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _0769_
timestamp 1676037725
transform 1 0 27508 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0770_
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0771_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0773_
timestamp 1676037725
transform 1 0 30544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0774_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0775_
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0776_
timestamp 1676037725
transform 1 0 36616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0777_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0778_
timestamp 1676037725
transform 1 0 36524 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 1676037725
transform 1 0 35788 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0780_
timestamp 1676037725
transform 1 0 37260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1676037725
transform 1 0 36616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0782_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0784_
timestamp 1676037725
transform 1 0 44712 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0785_
timestamp 1676037725
transform 1 0 45172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0786_
timestamp 1676037725
transform 1 0 38548 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0787_
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0788_
timestamp 1676037725
transform 1 0 44436 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0789_
timestamp 1676037725
transform 1 0 42412 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0790_
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0791_
timestamp 1676037725
transform 1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0792_
timestamp 1676037725
transform 1 0 45172 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _0793_
timestamp 1676037725
transform 1 0 42872 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0794_
timestamp 1676037725
transform 1 0 41400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0795_
timestamp 1676037725
transform 1 0 44436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0796_
timestamp 1676037725
transform 1 0 45172 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0797_
timestamp 1676037725
transform 1 0 41492 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0798_
timestamp 1676037725
transform 1 0 46460 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0799_
timestamp 1676037725
transform 1 0 45908 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0800_
timestamp 1676037725
transform 1 0 45540 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0801_
timestamp 1676037725
transform 1 0 45448 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47380 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0803_
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0804_
timestamp 1676037725
transform 1 0 44896 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0805_
timestamp 1676037725
transform 1 0 42596 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0806_
timestamp 1676037725
transform 1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _0807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0808_
timestamp 1676037725
transform 1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1676037725
transform 1 0 10212 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0810_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__and2b_1  _0812_
timestamp 1676037725
transform 1 0 10304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0813_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _0814_
timestamp 1676037725
transform 1 0 9844 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0815_
timestamp 1676037725
transform 1 0 4876 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0816_
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0817_
timestamp 1676037725
transform 1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1676037725
transform 1 0 12512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0819_
timestamp 1676037725
transform 1 0 12880 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0820_
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1676037725
transform 1 0 6808 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0822_
timestamp 1676037725
transform 1 0 7268 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0823_
timestamp 1676037725
transform 1 0 12144 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0824_
timestamp 1676037725
transform 1 0 10304 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp 1676037725
transform 1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0827_
timestamp 1676037725
transform 1 0 8004 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0828_
timestamp 1676037725
transform 1 0 11040 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0829_
timestamp 1676037725
transform 1 0 10488 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0830_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0831_
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0832_
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0833_
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0834_
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0835_
timestamp 1676037725
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0836_
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0837_
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0838_
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0839_
timestamp 1676037725
transform 1 0 16192 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0840_
timestamp 1676037725
transform 1 0 23276 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0841_
timestamp 1676037725
transform 1 0 17020 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0842_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0843_
timestamp 1676037725
transform 1 0 17296 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0845_
timestamp 1676037725
transform 1 0 15824 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0846_
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0847_
timestamp 1676037725
transform 1 0 20424 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1676037725
transform 1 0 20884 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0849_
timestamp 1676037725
transform 1 0 19872 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0851_
timestamp 1676037725
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0852_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0853_
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1676037725
transform 1 0 14444 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0855_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0856_
timestamp 1676037725
transform 1 0 27140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0857_
timestamp 1676037725
transform 1 0 23644 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0858_
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0859_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0861_
timestamp 1676037725
transform 1 0 16376 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0862_
timestamp 1676037725
transform 1 0 16928 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0863_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0864_
timestamp 1676037725
transform 1 0 27416 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0865_
timestamp 1676037725
transform 1 0 25668 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0866_
timestamp 1676037725
transform 1 0 25484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0867_
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0868_
timestamp 1676037725
transform 1 0 28336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0869_
timestamp 1676037725
transform 1 0 21620 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0870_
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0871_
timestamp 1676037725
transform 1 0 21620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0872_
timestamp 1676037725
transform 1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0873_
timestamp 1676037725
transform 1 0 20424 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0874_
timestamp 1676037725
transform 1 0 19412 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0875_
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0876_
timestamp 1676037725
transform 1 0 33120 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0877_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0878_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0879_
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0880_
timestamp 1676037725
transform 1 0 33212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0881_
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0882_
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0883_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0884_
timestamp 1676037725
transform 1 0 33856 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0885_
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0886_
timestamp 1676037725
transform 1 0 23552 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0887_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0888_
timestamp 1676037725
transform 1 0 25852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0889_
timestamp 1676037725
transform 1 0 36064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0890_
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0891_
timestamp 1676037725
transform 1 0 24380 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0893_
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0894_
timestamp 1676037725
transform 1 0 26772 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0895_
timestamp 1676037725
transform 1 0 25760 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0897_
timestamp 1676037725
transform 1 0 40020 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0898_
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0899_
timestamp 1676037725
transform 1 0 26404 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1676037725
transform 1 0 12788 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0901_
timestamp 1676037725
transform 1 0 39928 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0902_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0903_
timestamp 1676037725
transform 1 0 25760 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1676037725
transform 1 0 9844 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0905_
timestamp 1676037725
transform 1 0 43240 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0906_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0907_
timestamp 1676037725
transform 1 0 25760 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1676037725
transform 1 0 25116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0909_
timestamp 1676037725
transform 1 0 43700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0910_
timestamp 1676037725
transform 1 0 26036 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0911_
timestamp 1676037725
transform 1 0 25944 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1676037725
transform 1 0 24748 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0913_
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0914_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0915_
timestamp 1676037725
transform 1 0 23460 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _0917_
timestamp 1676037725
transform 1 0 43700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0918_
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0919_
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0920_
timestamp 1676037725
transform 1 0 22172 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0921_
timestamp 1676037725
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0922_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0923_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0924_
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0925_
timestamp 1676037725
transform 1 0 9476 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0926_
timestamp 1676037725
transform 1 0 4324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0927_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0928_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0929_
timestamp 1676037725
transform 1 0 3680 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0930_
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0931_
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1676037725
transform 1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0933_
timestamp 1676037725
transform 1 0 4416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0937_
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1676037725
transform 1 0 1932 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp 1676037725
transform 1 0 6992 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1676037725
transform 1 0 7360 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0943_
timestamp 1676037725
transform 1 0 2944 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 1676037725
transform 1 0 6624 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1676037725
transform 1 0 2208 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1676037725
transform 1 0 4416 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1676037725
transform 1 0 6256 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp 1676037725
transform 1 0 3772 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 1676037725
transform 1 0 10304 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1676037725
transform 1 0 7452 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1676037725
transform 1 0 10212 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0957_
timestamp 1676037725
transform 1 0 38548 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0959_
timestamp 1676037725
transform 1 0 5336 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _0963_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0964_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1676037725
transform 1 0 13340 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1676037725
transform 1 0 18768 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0969_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1676037725
transform 1 0 20884 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1676037725
transform 1 0 21344 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1676037725
transform 1 0 11500 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1676037725
transform 1 0 13248 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1676037725
transform 1 0 25852 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1676037725
transform 1 0 22632 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1676037725
transform 1 0 20976 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1676037725
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform 1 0 30360 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 28612 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1676037725
transform 1 0 29808 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1676037725
transform 1 0 40204 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1676037725
transform 1 0 28704 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1676037725
transform 1 0 18308 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1676037725
transform 1 0 36340 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1676037725
transform 1 0 41308 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1676037725
transform 1 0 41124 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1676037725
transform 1 0 38088 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1002_
timestamp 1676037725
transform 1 0 38640 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1676037725
transform 1 0 41216 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1676037725
transform 1 0 41032 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1005_
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1676037725
transform 1 0 38180 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1676037725
transform 1 0 33948 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1676037725
transform 1 0 35972 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1676037725
transform 1 0 40664 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1676037725
transform 1 0 40664 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1676037725
transform 1 0 41308 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1676037725
transform 1 0 41308 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1013_
timestamp 1676037725
transform 1 0 41492 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1014_
timestamp 1676037725
transform 1 0 39652 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1015_
timestamp 1676037725
transform 1 0 35328 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1676037725
transform 1 0 35328 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1676037725
transform 1 0 37168 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1676037725
transform 1 0 32016 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1022_
timestamp 1676037725
transform 1 0 28244 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1023_
timestamp 1676037725
transform 1 0 30268 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1024_
timestamp 1676037725
transform 1 0 33856 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1025_
timestamp 1676037725
transform 1 0 31924 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1026_
timestamp 1676037725
transform 1 0 35880 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1676037725
transform 1 0 28704 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1676037725
transform 1 0 25760 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1029_
timestamp 1676037725
transform 1 0 26128 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 29348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 32936 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1676037725
transform 1 0 32936 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1033_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27324 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1034_
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1035_
timestamp 1676037725
transform 1 0 29716 0 1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1676037725
transform 1 0 26220 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1038_
timestamp 1676037725
transform 1 0 36524 0 1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1039_
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1676037725
transform 1 0 36984 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1041_
timestamp 1676037725
transform 1 0 40572 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1042_
timestamp 1676037725
transform 1 0 40388 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1044_
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1045_
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1046_
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1047_
timestamp 1676037725
transform 1 0 13892 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 18952 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1049_
timestamp 1676037725
transform 1 0 22540 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1050_
timestamp 1676037725
transform 1 0 25944 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1052_
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1056_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1676037725
transform 1 0 36524 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1059_
timestamp 1676037725
transform 1 0 36616 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1676037725
transform 1 0 40204 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 40664 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1062_
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1676037725
transform 1 0 42136 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1676037725
transform 1 0 40296 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1676037725
transform 1 0 41124 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1066_
timestamp 1676037725
transform 1 0 11408 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1676037725
transform 1 0 10212 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1676037725
transform 1 0 4600 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1676037725
transform 1 0 12328 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1676037725
transform 1 0 17480 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1676037725
transform 1 0 17480 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1078_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1079_
timestamp 1676037725
transform 1 0 17940 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1676037725
transform 1 0 12972 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1676037725
transform 1 0 10764 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1676037725
transform 1 0 8280 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1676037725
transform 1 0 12144 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1087_
timestamp 1676037725
transform 1 0 24748 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1676037725
transform 1 0 24196 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1089_
timestamp 1676037725
transform 1 0 22356 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1091_
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1092_
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1093_
timestamp 1676037725
transform 1 0 5152 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1094_
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1095_
timestamp 1676037725
transform 1 0 8464 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1096_
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1097_
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1098_
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1676037725
transform 1 0 1656 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1676037725
transform 1 0 1656 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1676037725
transform 1 0 1656 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1676037725
transform 1 0 1656 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1676037725
transform 1 0 6808 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1676037725
transform 1 0 7636 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1676037725
transform 1 0 2668 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1676037725
transform 1 0 6348 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1676037725
transform 1 0 1840 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1676037725
transform 1 0 1932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1676037725
transform 1 0 1656 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1676037725
transform 1 0 4048 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1676037725
transform 1 0 5336 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1676037725
transform 1 0 10212 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1676037725
transform 1 0 7176 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1676037725
transform 1 0 2024 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1676037725
transform 1 0 9752 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1123_
timestamp 1676037725
transform 1 0 40756 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1124_
timestamp 1676037725
transform 1 0 5428 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1125_
timestamp 1676037725
transform 1 0 6900 0 -1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1126_
timestamp 1676037725
transform 1 0 1840 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1127_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1128_
timestamp 1676037725
transform 1 0 1748 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1139_
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1676037725
transform 1 0 9384 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1676037725
transform 1 0 14444 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1676037725
transform 1 0 14444 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1676037725
transform 1 0 15088 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1676037725
transform 1 0 30084 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1676037725
transform 1 0 30084 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1676037725
transform 1 0 35972 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1676037725
transform 1 0 36432 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1676037725
transform 1 0 29992 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1676037725
transform 1 0 30176 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1676037725
transform 1 0 36340 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1676037725
transform 1 0 36340 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout178 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout179
timestamp 1676037725
transform 1 0 19964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout180 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout181
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout182
timestamp 1676037725
transform 1 0 33304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout183
timestamp 1676037725
transform 1 0 37812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout184
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout185 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout186
timestamp 1676037725
transform 1 0 5888 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout187
timestamp 1676037725
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout188
timestamp 1676037725
transform 1 0 10120 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout189
timestamp 1676037725
transform 1 0 28888 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout190
timestamp 1676037725
transform 1 0 10672 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout191
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout192
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout193
timestamp 1676037725
transform 1 0 34960 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout194
timestamp 1676037725
transform 1 0 22080 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout195
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout196
timestamp 1676037725
transform 1 0 19504 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout197
timestamp 1676037725
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout198
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout199
timestamp 1676037725
transform 1 0 20976 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout200
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout201
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout202
timestamp 1676037725
transform 1 0 27968 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout203
timestamp 1676037725
transform 1 0 10120 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout204
timestamp 1676037725
transform 1 0 9476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout205
timestamp 1676037725
transform 1 0 10212 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout206
timestamp 1676037725
transform 1 0 29348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout207
timestamp 1676037725
transform 1 0 28520 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout208
timestamp 1676037725
transform 1 0 10396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout209
timestamp 1676037725
transform 1 0 33304 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout210
timestamp 1676037725
transform 1 0 7728 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout211
timestamp 1676037725
transform 1 0 7820 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout212
timestamp 1676037725
transform 1 0 2576 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout213
timestamp 1676037725
transform 1 0 8096 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout214
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout215
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout216
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout217
timestamp 1676037725
transform 1 0 9292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout218
timestamp 1676037725
transform 1 0 36984 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout219
timestamp 1676037725
transform 1 0 44068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout220
timestamp 1676037725
transform 1 0 10856 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout221
timestamp 1676037725
transform 1 0 9936 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout222
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout223
timestamp 1676037725
transform 1 0 15824 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout224
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout225
timestamp 1676037725
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout226
timestamp 1676037725
transform 1 0 32936 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout227
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout228
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout229
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout230
timestamp 1676037725
transform 1 0 35512 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout231
timestamp 1676037725
transform 1 0 28336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout232
timestamp 1676037725
transform 1 0 30636 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout233
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout234
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout235
timestamp 1676037725
transform 1 0 36432 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout236
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout237
timestamp 1676037725
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33764 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1676037725
transform 1 0 33120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 34592 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 38732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 45632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 47748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1676037725
transform 1 0 50324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1676037725
transform 1 0 51244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1676037725
transform 1 0 52900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1676037725
transform 1 0 53912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input23
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input25
timestamp 1676037725
transform 1 0 56672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1676037725
transform 1 0 55752 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1676037725
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1676037725
transform 1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1676037725
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1676037725
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1676037725
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 3772 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform 1 0 3128 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1676037725
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1676037725
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input60
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input63
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input64
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input65
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input68
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input69
timestamp 1676037725
transform 1 0 1564 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1676037725
transform 1 0 2300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1676037725
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1676037725
transform 1 0 2300 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input76
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1676037725
transform 1 0 3128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1676037725
transform 1 0 3128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input81
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1676037725
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output87
timestamp 1676037725
transform 1 0 3956 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output88
timestamp 1676037725
transform 1 0 27140 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output89
timestamp 1676037725
transform 1 0 56120 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output90
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output91
timestamp 1676037725
transform 1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output92
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output93
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output94
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output95
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output96
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output97
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output98
timestamp 1676037725
transform 1 0 23552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output99
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output100
timestamp 1676037725
transform 1 0 6992 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output101
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output102
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output103
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output104
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output105
timestamp 1676037725
transform 1 0 20332 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output106
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output107
timestamp 1676037725
transform 1 0 24932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1676037725
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output110
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output111
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output112
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output113
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output114
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output115
timestamp 1676037725
transform 1 0 30912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output116
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output117
timestamp 1676037725
transform 1 0 33672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output118
timestamp 1676037725
transform 1 0 35972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output119
timestamp 1676037725
transform 1 0 36432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output120
timestamp 1676037725
transform 1 0 37812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output121
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output122
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output123
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output124
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output125
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output126
timestamp 1676037725
transform 1 0 45172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output127
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output128
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output129
timestamp 1676037725
transform 1 0 48852 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output130
timestamp 1676037725
transform 1 0 50232 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output131
timestamp 1676037725
transform 1 0 51612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output132
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output133
timestamp 1676037725
transform 1 0 54832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output134
timestamp 1676037725
transform 1 0 10672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output135
timestamp 1676037725
transform 1 0 56396 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output136
timestamp 1676037725
transform 1 0 57132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output137
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output138
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output139
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output140
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output141
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output142
timestamp 1676037725
transform 1 0 25392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output143
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output144
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output145
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output146
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output147
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output148
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output149
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output150
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output151
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output152
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output153
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output154
timestamp 1676037725
transform 1 0 1564 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output155
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output156
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output157
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output158
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output159
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output160
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output161
timestamp 1676037725
transform 1 0 1564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output162
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output163
timestamp 1676037725
transform 1 0 1564 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output164
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output165
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output166
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output167
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output168
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output169
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output170
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output171
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output172
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output173
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output174
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output175
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output176
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output177
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
<< labels >>
flabel metal2 s 3882 41200 3938 42000 0 FreeSans 224 90 0 0 flash_csb
port 0 nsew signal tristate
flabel metal2 s 11334 41200 11390 42000 0 FreeSans 224 90 0 0 flash_io0_read
port 1 nsew signal input
flabel metal2 s 18786 41200 18842 42000 0 FreeSans 224 90 0 0 flash_io0_we
port 2 nsew signal tristate
flabel metal2 s 26238 41200 26294 42000 0 FreeSans 224 90 0 0 flash_io0_write
port 3 nsew signal tristate
flabel metal2 s 33690 41200 33746 42000 0 FreeSans 224 90 0 0 flash_io1_read
port 4 nsew signal input
flabel metal2 s 41142 41200 41198 42000 0 FreeSans 224 90 0 0 flash_io1_we
port 5 nsew signal tristate
flabel metal2 s 48594 41200 48650 42000 0 FreeSans 224 90 0 0 flash_io1_write
port 6 nsew signal tristate
flabel metal2 s 56046 41200 56102 42000 0 FreeSans 224 90 0 0 flash_sck
port 7 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 sram_addr0[0]
port 8 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 sram_addr0[1]
port 9 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 sram_addr0[2]
port 10 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 sram_addr0[3]
port 11 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 sram_addr0[4]
port 12 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 sram_addr0[5]
port 13 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 sram_addr0[6]
port 14 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 sram_addr0[7]
port 15 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 sram_addr0[8]
port 16 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 sram_addr1[0]
port 17 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 sram_addr1[1]
port 18 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 sram_addr1[2]
port 19 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 sram_addr1[3]
port 20 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 sram_addr1[4]
port 21 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 sram_addr1[5]
port 22 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 sram_addr1[6]
port 23 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 sram_addr1[7]
port 24 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 sram_addr1[8]
port 25 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 sram_clk0
port 26 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 sram_clk1
port 27 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 sram_csb0
port 28 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 sram_csb1
port 29 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 sram_din0[0]
port 30 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 sram_din0[10]
port 31 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 sram_din0[11]
port 32 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 sram_din0[12]
port 33 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 sram_din0[13]
port 34 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 sram_din0[14]
port 35 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 sram_din0[15]
port 36 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 sram_din0[16]
port 37 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 sram_din0[17]
port 38 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 sram_din0[18]
port 39 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 sram_din0[19]
port 40 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 sram_din0[1]
port 41 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 sram_din0[20]
port 42 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 sram_din0[21]
port 43 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 sram_din0[22]
port 44 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 sram_din0[23]
port 45 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 sram_din0[24]
port 46 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 sram_din0[25]
port 47 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 sram_din0[26]
port 48 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 sram_din0[27]
port 49 nsew signal tristate
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 sram_din0[28]
port 50 nsew signal tristate
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 sram_din0[29]
port 51 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 sram_din0[2]
port 52 nsew signal tristate
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 sram_din0[30]
port 53 nsew signal tristate
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 sram_din0[31]
port 54 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 sram_din0[3]
port 55 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 sram_din0[4]
port 56 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 sram_din0[5]
port 57 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 sram_din0[6]
port 58 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 sram_din0[7]
port 59 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 sram_din0[8]
port 60 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 sram_din0[9]
port 61 nsew signal tristate
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 sram_dout0[0]
port 62 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 sram_dout0[10]
port 63 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 sram_dout0[11]
port 64 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 sram_dout0[12]
port 65 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 sram_dout0[13]
port 66 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 sram_dout0[14]
port 67 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 sram_dout0[15]
port 68 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 sram_dout0[16]
port 69 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 sram_dout0[17]
port 70 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 sram_dout0[18]
port 71 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 sram_dout0[19]
port 72 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 sram_dout0[1]
port 73 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 sram_dout0[20]
port 74 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 sram_dout0[21]
port 75 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 sram_dout0[22]
port 76 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 sram_dout0[23]
port 77 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 sram_dout0[24]
port 78 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 sram_dout0[25]
port 79 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 sram_dout0[26]
port 80 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 sram_dout0[27]
port 81 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 sram_dout0[28]
port 82 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 sram_dout0[29]
port 83 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 sram_dout0[2]
port 84 nsew signal input
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 sram_dout0[30]
port 85 nsew signal input
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 sram_dout0[31]
port 86 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 sram_dout0[3]
port 87 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 sram_dout0[4]
port 88 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 sram_dout0[5]
port 89 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 sram_dout0[6]
port 90 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 sram_dout0[7]
port 91 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 sram_dout0[8]
port 92 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 sram_dout0[9]
port 93 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 sram_dout1[0]
port 94 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 sram_dout1[10]
port 95 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 sram_dout1[11]
port 96 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 sram_dout1[12]
port 97 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 sram_dout1[13]
port 98 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 sram_dout1[14]
port 99 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 sram_dout1[15]
port 100 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 sram_dout1[16]
port 101 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 sram_dout1[17]
port 102 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 sram_dout1[18]
port 103 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 sram_dout1[19]
port 104 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 sram_dout1[1]
port 105 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 sram_dout1[20]
port 106 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 sram_dout1[21]
port 107 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 sram_dout1[22]
port 108 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 sram_dout1[23]
port 109 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 sram_dout1[24]
port 110 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 sram_dout1[25]
port 111 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 sram_dout1[26]
port 112 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 sram_dout1[27]
port 113 nsew signal input
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 sram_dout1[28]
port 114 nsew signal input
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 sram_dout1[29]
port 115 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 sram_dout1[2]
port 116 nsew signal input
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 sram_dout1[30]
port 117 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 sram_dout1[31]
port 118 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 sram_dout1[3]
port 119 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 sram_dout1[4]
port 120 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 sram_dout1[5]
port 121 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 sram_dout1[6]
port 122 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 sram_dout1[7]
port 123 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 sram_dout1[8]
port 124 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 sram_dout1[9]
port 125 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 sram_web0
port 126 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 sram_wmask0[0]
port 127 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 sram_wmask0[1]
port 128 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 sram_wmask0[2]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 sram_wmask0[3]
port 130 nsew signal tristate
flabel metal4 s 4208 2128 4528 39760 0 FreeSans 1920 90 0 0 vccd1
port 131 nsew power bidirectional
flabel metal4 s 34928 2128 35248 39760 0 FreeSans 1920 90 0 0 vccd1
port 131 nsew power bidirectional
flabel metal4 s 19568 2128 19888 39760 0 FreeSans 1920 90 0 0 vssd1
port 132 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 39760 0 FreeSans 1920 90 0 0 vssd1
port 132 nsew ground bidirectional
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 wb_ack_o
port 133 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 wb_adr_i[0]
port 134 nsew signal input
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 wb_adr_i[10]
port 135 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 wb_adr_i[11]
port 136 nsew signal input
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 wb_adr_i[12]
port 137 nsew signal input
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 wb_adr_i[13]
port 138 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 wb_adr_i[14]
port 139 nsew signal input
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 wb_adr_i[15]
port 140 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 wb_adr_i[16]
port 141 nsew signal input
flabel metal3 s 0 26392 800 26512 0 FreeSans 480 0 0 0 wb_adr_i[17]
port 142 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 wb_adr_i[18]
port 143 nsew signal input
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 wb_adr_i[19]
port 144 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 wb_adr_i[1]
port 145 nsew signal input
flabel metal3 s 0 30064 800 30184 0 FreeSans 480 0 0 0 wb_adr_i[20]
port 146 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 wb_adr_i[21]
port 147 nsew signal input
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 wb_adr_i[22]
port 148 nsew signal input
flabel metal3 s 0 33736 800 33856 0 FreeSans 480 0 0 0 wb_adr_i[23]
port 149 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 wb_adr_i[2]
port 150 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 wb_adr_i[3]
port 151 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 wb_adr_i[4]
port 152 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 wb_adr_i[5]
port 153 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 wb_adr_i[6]
port 154 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 wb_adr_i[7]
port 155 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 wb_adr_i[8]
port 156 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 wb_adr_i[9]
port 157 nsew signal input
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 wb_clk_i
port 158 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 wb_cyc_i
port 159 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 wb_data_i[0]
port 160 nsew signal input
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 wb_data_i[10]
port 161 nsew signal input
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 wb_data_i[11]
port 162 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 wb_data_i[12]
port 163 nsew signal input
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 wb_data_i[13]
port 164 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 wb_data_i[14]
port 165 nsew signal input
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 wb_data_i[15]
port 166 nsew signal input
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 wb_data_i[16]
port 167 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 wb_data_i[17]
port 168 nsew signal input
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 wb_data_i[18]
port 169 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 wb_data_i[19]
port 170 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 wb_data_i[1]
port 171 nsew signal input
flabel metal3 s 0 30472 800 30592 0 FreeSans 480 0 0 0 wb_data_i[20]
port 172 nsew signal input
flabel metal3 s 0 31696 800 31816 0 FreeSans 480 0 0 0 wb_data_i[21]
port 173 nsew signal input
flabel metal3 s 0 32920 800 33040 0 FreeSans 480 0 0 0 wb_data_i[22]
port 174 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 wb_data_i[23]
port 175 nsew signal input
flabel metal3 s 0 34960 800 35080 0 FreeSans 480 0 0 0 wb_data_i[24]
port 176 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 wb_data_i[25]
port 177 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 wb_data_i[26]
port 178 nsew signal input
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 wb_data_i[27]
port 179 nsew signal input
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 wb_data_i[28]
port 180 nsew signal input
flabel metal3 s 0 39040 800 39160 0 FreeSans 480 0 0 0 wb_data_i[29]
port 181 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 wb_data_i[2]
port 182 nsew signal input
flabel metal3 s 0 39856 800 39976 0 FreeSans 480 0 0 0 wb_data_i[30]
port 183 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 wb_data_i[31]
port 184 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 wb_data_i[3]
port 185 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 wb_data_i[4]
port 186 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 wb_data_i[5]
port 187 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 wb_data_i[6]
port 188 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 wb_data_i[7]
port 189 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 wb_data_i[8]
port 190 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 wb_data_i[9]
port 191 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 wb_data_o[0]
port 192 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 wb_data_o[10]
port 193 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 wb_data_o[11]
port 194 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 wb_data_o[12]
port 195 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 wb_data_o[13]
port 196 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 wb_data_o[14]
port 197 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 wb_data_o[15]
port 198 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 wb_data_o[16]
port 199 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 wb_data_o[17]
port 200 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 wb_data_o[18]
port 201 nsew signal tristate
flabel metal3 s 0 29656 800 29776 0 FreeSans 480 0 0 0 wb_data_o[19]
port 202 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 wb_data_o[1]
port 203 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 wb_data_o[20]
port 204 nsew signal tristate
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 wb_data_o[21]
port 205 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 wb_data_o[22]
port 206 nsew signal tristate
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 wb_data_o[23]
port 207 nsew signal tristate
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 wb_data_o[24]
port 208 nsew signal tristate
flabel metal3 s 0 36184 800 36304 0 FreeSans 480 0 0 0 wb_data_o[25]
port 209 nsew signal tristate
flabel metal3 s 0 37000 800 37120 0 FreeSans 480 0 0 0 wb_data_o[26]
port 210 nsew signal tristate
flabel metal3 s 0 37816 800 37936 0 FreeSans 480 0 0 0 wb_data_o[27]
port 211 nsew signal tristate
flabel metal3 s 0 38632 800 38752 0 FreeSans 480 0 0 0 wb_data_o[28]
port 212 nsew signal tristate
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 wb_data_o[29]
port 213 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 wb_data_o[2]
port 214 nsew signal tristate
flabel metal3 s 0 40264 800 40384 0 FreeSans 480 0 0 0 wb_data_o[30]
port 215 nsew signal tristate
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 wb_data_o[31]
port 216 nsew signal tristate
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 wb_data_o[3]
port 217 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 wb_data_o[4]
port 218 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 wb_data_o[5]
port 219 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 wb_data_o[6]
port 220 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 wb_data_o[7]
port 221 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 wb_data_o[8]
port 222 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 wb_data_o[9]
port 223 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 wb_error_o
port 224 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 wb_rst_i
port 225 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 wb_sel_i[0]
port 226 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 wb_sel_i[1]
port 227 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 wb_sel_i[2]
port 228 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 wb_sel_i[3]
port 229 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 wb_stall_o
port 230 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 wb_stb_i
port 231 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 wb_we_i
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
<< end >>
