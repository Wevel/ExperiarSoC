magic
tech sky130A
magscale 1 2
timestamp 1651278039
<< viali >>
rect 2053 37417 2087 37451
rect 2697 37349 2731 37383
rect 1409 37213 1443 37247
rect 20085 37213 20119 37247
rect 35817 37213 35851 37247
rect 36461 37213 36495 37247
rect 37841 37213 37875 37247
rect 20269 37077 20303 37111
rect 36001 37077 36035 37111
rect 36645 37077 36679 37111
rect 37289 37077 37323 37111
rect 38025 37077 38059 37111
rect 36093 36873 36127 36907
rect 38025 36873 38059 36907
rect 1409 36737 1443 36771
rect 37381 36737 37415 36771
rect 37841 36737 37875 36771
rect 19441 36329 19475 36363
rect 38025 36329 38059 36363
rect 1409 36125 1443 36159
rect 19257 36125 19291 36159
rect 19901 36125 19935 36159
rect 36737 36125 36771 36159
rect 37381 36125 37415 36159
rect 37841 36125 37875 36159
rect 37197 35989 37231 36023
rect 37841 35649 37875 35683
rect 1409 35445 1443 35479
rect 38025 35445 38059 35479
rect 37841 35037 37875 35071
rect 37289 34901 37323 34935
rect 38025 34901 38059 34935
rect 1409 34425 1443 34459
rect 1409 33949 1443 33983
rect 37473 33949 37507 33983
rect 38117 33949 38151 33983
rect 37933 33813 37967 33847
rect 37841 33473 37875 33507
rect 38025 33269 38059 33303
rect 1409 32861 1443 32895
rect 37289 32861 37323 32895
rect 37841 32861 37875 32895
rect 38025 32725 38059 32759
rect 37473 32385 37507 32419
rect 38117 32385 38151 32419
rect 37933 32181 37967 32215
rect 1409 31773 1443 31807
rect 1409 31297 1443 31331
rect 2053 31297 2087 31331
rect 37841 31297 37875 31331
rect 1593 31093 1627 31127
rect 38025 31093 38059 31127
rect 1409 30685 1443 30719
rect 2053 30685 2087 30719
rect 37841 30685 37875 30719
rect 1593 30549 1627 30583
rect 37289 30549 37323 30583
rect 38025 30549 38059 30583
rect 37473 30209 37507 30243
rect 38117 30209 38151 30243
rect 1409 30005 1443 30039
rect 37933 30005 37967 30039
rect 1409 29597 1443 29631
rect 2053 29597 2087 29631
rect 1593 29461 1627 29495
rect 2513 29121 2547 29155
rect 2789 29121 2823 29155
rect 37841 29121 37875 29155
rect 2605 29053 2639 29087
rect 1409 28985 1443 29019
rect 2973 28985 3007 29019
rect 38025 28985 38059 29019
rect 2513 28917 2547 28951
rect 37841 28509 37875 28543
rect 37289 28373 37323 28407
rect 38025 28373 38059 28407
rect 1593 28169 1627 28203
rect 32137 28169 32171 28203
rect 1409 28033 1443 28067
rect 2053 28033 2087 28067
rect 33250 28033 33284 28067
rect 37473 28033 37507 28067
rect 38117 28033 38151 28067
rect 33517 27965 33551 27999
rect 37933 27829 37967 27863
rect 25789 27557 25823 27591
rect 33057 27557 33091 27591
rect 36093 27557 36127 27591
rect 1409 27421 1443 27455
rect 22293 27421 22327 27455
rect 24409 27421 24443 27455
rect 31033 27421 31067 27455
rect 32873 27421 32907 27455
rect 34713 27421 34747 27455
rect 37841 27421 37875 27455
rect 22538 27353 22572 27387
rect 24676 27353 24710 27387
rect 31278 27353 31312 27387
rect 34958 27353 34992 27387
rect 36829 27353 36863 27387
rect 23673 27285 23707 27319
rect 32413 27285 32447 27319
rect 33609 27285 33643 27319
rect 37289 27285 37323 27319
rect 38025 27285 38059 27319
rect 22477 27081 22511 27115
rect 24869 27081 24903 27115
rect 28365 27081 28399 27115
rect 30573 27081 30607 27115
rect 34161 27081 34195 27115
rect 37933 27081 37967 27115
rect 23182 27013 23216 27047
rect 29929 27013 29963 27047
rect 31033 27013 31067 27047
rect 1409 26945 1443 26979
rect 2053 26945 2087 26979
rect 22293 26945 22327 26979
rect 22937 26945 22971 26979
rect 25053 26945 25087 26979
rect 26985 26945 27019 26979
rect 27241 26945 27275 26979
rect 30389 26945 30423 26979
rect 32137 26945 32171 26979
rect 32393 26945 32427 26979
rect 33977 26945 34011 26979
rect 38117 26945 38151 26979
rect 31401 26809 31435 26843
rect 1593 26741 1627 26775
rect 24317 26741 24351 26775
rect 31493 26741 31527 26775
rect 33517 26741 33551 26775
rect 36645 26741 36679 26775
rect 37473 26741 37507 26775
rect 22385 26537 22419 26571
rect 23489 26537 23523 26571
rect 26433 26537 26467 26571
rect 30849 26537 30883 26571
rect 31953 26537 31987 26571
rect 34069 26537 34103 26571
rect 36277 26537 36311 26571
rect 23397 26469 23431 26503
rect 25053 26469 25087 26503
rect 30297 26469 30331 26503
rect 30941 26469 30975 26503
rect 33149 26469 33183 26503
rect 33885 26469 33919 26503
rect 38025 26469 38059 26503
rect 30389 26401 30423 26435
rect 32597 26401 32631 26435
rect 32689 26401 32723 26435
rect 1685 26333 1719 26367
rect 22569 26333 22603 26367
rect 26249 26333 26283 26367
rect 28273 26333 28307 26367
rect 31769 26333 31803 26367
rect 33609 26333 33643 26367
rect 36875 26333 36909 26367
rect 37013 26333 37047 26367
rect 37105 26333 37139 26367
rect 37288 26333 37322 26367
rect 37381 26333 37415 26367
rect 37841 26333 37875 26367
rect 2237 26265 2271 26299
rect 21925 26265 21959 26299
rect 23029 26265 23063 26299
rect 24409 26265 24443 26299
rect 28006 26265 28040 26299
rect 29929 26265 29963 26299
rect 31309 26265 31343 26299
rect 32781 26265 32815 26299
rect 34713 26265 34747 26299
rect 1501 26197 1535 26231
rect 26893 26197 26927 26231
rect 36737 26197 36771 26231
rect 22201 25993 22235 26027
rect 26985 25993 27019 26027
rect 27905 25993 27939 26027
rect 30849 25993 30883 26027
rect 32137 25993 32171 26027
rect 32597 25993 32631 26027
rect 31309 25925 31343 25959
rect 37657 25925 37691 25959
rect 1409 25857 1443 25891
rect 2329 25857 2363 25891
rect 23489 25857 23523 25891
rect 28089 25857 28123 25891
rect 30389 25857 30423 25891
rect 31217 25857 31251 25891
rect 32505 25857 32539 25891
rect 35633 25857 35667 25891
rect 36272 25857 36306 25891
rect 36369 25857 36403 25891
rect 36461 25857 36495 25891
rect 36644 25857 36678 25891
rect 36737 25857 36771 25891
rect 37560 25857 37594 25891
rect 37749 25857 37783 25891
rect 37932 25857 37966 25891
rect 38025 25857 38059 25891
rect 1685 25789 1719 25823
rect 22661 25789 22695 25823
rect 23581 25789 23615 25823
rect 23765 25789 23799 25823
rect 25237 25789 25271 25823
rect 25789 25789 25823 25823
rect 27445 25789 27479 25823
rect 31493 25789 31527 25823
rect 32689 25789 32723 25823
rect 22385 25721 22419 25755
rect 27077 25721 27111 25755
rect 33885 25721 33919 25755
rect 35081 25721 35115 25755
rect 21189 25653 21223 25687
rect 23121 25653 23155 25687
rect 24409 25653 24443 25687
rect 33333 25653 33367 25687
rect 36093 25653 36127 25687
rect 37381 25653 37415 25687
rect 22661 25449 22695 25483
rect 23121 25449 23155 25483
rect 24409 25449 24443 25483
rect 25697 25449 25731 25483
rect 28457 25449 28491 25483
rect 31585 25449 31619 25483
rect 1593 25381 1627 25415
rect 22569 25381 22603 25415
rect 36921 25381 36955 25415
rect 23581 25313 23615 25347
rect 23765 25313 23799 25347
rect 25053 25313 25087 25347
rect 32229 25313 32263 25347
rect 33333 25313 33367 25347
rect 35541 25313 35575 25347
rect 1409 25245 1443 25279
rect 2053 25245 2087 25279
rect 24869 25245 24903 25279
rect 27077 25245 27111 25279
rect 32045 25245 32079 25279
rect 37381 25245 37415 25279
rect 37474 25245 37508 25279
rect 37749 25245 37783 25279
rect 37846 25245 37880 25279
rect 22201 25177 22235 25211
rect 27322 25177 27356 25211
rect 31953 25177 31987 25211
rect 35786 25177 35820 25211
rect 37657 25177 37691 25211
rect 2697 25109 2731 25143
rect 21649 25109 21683 25143
rect 23489 25109 23523 25143
rect 24777 25109 24811 25143
rect 26249 25109 26283 25143
rect 30573 25109 30607 25143
rect 31125 25109 31159 25143
rect 32781 25109 32815 25143
rect 38025 25109 38059 25143
rect 26985 24905 27019 24939
rect 27353 24905 27387 24939
rect 1869 24769 1903 24803
rect 2697 24769 2731 24803
rect 23397 24769 23431 24803
rect 23581 24769 23615 24803
rect 26249 24769 26283 24803
rect 27445 24769 27479 24803
rect 28733 24769 28767 24803
rect 31401 24769 31435 24803
rect 35357 24769 35391 24803
rect 35624 24769 35658 24803
rect 37841 24769 37875 24803
rect 24593 24701 24627 24735
rect 27537 24701 27571 24735
rect 28273 24701 28307 24735
rect 2145 24633 2179 24667
rect 22753 24633 22787 24667
rect 36737 24633 36771 24667
rect 38025 24633 38059 24667
rect 22201 24565 22235 24599
rect 23213 24565 23247 24599
rect 24041 24565 24075 24599
rect 25145 24565 25179 24599
rect 26433 24565 26467 24599
rect 32505 24565 32539 24599
rect 37289 24565 37323 24599
rect 1501 24361 1535 24395
rect 24501 24361 24535 24395
rect 27169 24361 27203 24395
rect 35541 24361 35575 24395
rect 36001 24361 36035 24395
rect 36737 24361 36771 24395
rect 22109 24293 22143 24327
rect 24961 24293 24995 24327
rect 27077 24293 27111 24327
rect 27905 24293 27939 24327
rect 37381 24293 37415 24327
rect 22845 24225 22879 24259
rect 26709 24225 26743 24259
rect 1685 24157 1719 24191
rect 2145 24157 2179 24191
rect 2789 24157 2823 24191
rect 22549 24157 22583 24191
rect 22753 24157 22787 24191
rect 35357 24157 35391 24191
rect 36185 24157 36219 24191
rect 37841 24157 37875 24191
rect 22293 24089 22327 24123
rect 23673 24089 23707 24123
rect 23857 24089 23891 24123
rect 2329 24021 2363 24055
rect 22661 24021 22695 24055
rect 23489 24021 23523 24055
rect 28365 24021 28399 24055
rect 38025 24021 38059 24055
rect 22661 23817 22695 23851
rect 27445 23817 27479 23851
rect 22385 23749 22419 23783
rect 1685 23681 1719 23715
rect 2421 23681 2455 23715
rect 2513 23681 2547 23715
rect 2881 23681 2915 23715
rect 22155 23681 22189 23715
rect 22293 23681 22327 23715
rect 22477 23681 22511 23715
rect 23305 23681 23339 23715
rect 23489 23681 23523 23715
rect 23673 23681 23707 23715
rect 26433 23681 26467 23715
rect 27353 23681 27387 23715
rect 37473 23681 37507 23715
rect 38117 23681 38151 23715
rect 22017 23613 22051 23647
rect 24133 23613 24167 23647
rect 27537 23613 27571 23647
rect 28273 23613 28307 23647
rect 1501 23477 1535 23511
rect 2789 23477 2823 23511
rect 3065 23477 3099 23511
rect 3617 23477 3651 23511
rect 26985 23477 27019 23511
rect 28733 23477 28767 23511
rect 37933 23477 37967 23511
rect 24593 23273 24627 23307
rect 26709 23273 26743 23307
rect 29009 23273 29043 23307
rect 35173 23273 35207 23307
rect 26893 23205 26927 23239
rect 35081 23205 35115 23239
rect 2145 23137 2179 23171
rect 27169 23137 27203 23171
rect 27629 23137 27663 23171
rect 22477 23069 22511 23103
rect 22937 23069 22971 23103
rect 31401 23069 31435 23103
rect 37841 23069 37875 23103
rect 1869 23001 1903 23035
rect 2697 23001 2731 23035
rect 22293 23001 22327 23035
rect 22569 23001 22603 23035
rect 22661 23001 22695 23035
rect 22799 23001 22833 23035
rect 27874 23001 27908 23035
rect 31646 23001 31680 23035
rect 34713 23001 34747 23035
rect 23857 22933 23891 22967
rect 32781 22933 32815 22967
rect 38025 22933 38059 22967
rect 2329 22729 2363 22763
rect 24961 22729 24995 22763
rect 26433 22729 26467 22763
rect 27353 22729 27387 22763
rect 29469 22729 29503 22763
rect 31493 22729 31527 22763
rect 34161 22729 34195 22763
rect 34897 22729 34931 22763
rect 24225 22661 24259 22695
rect 37657 22661 37691 22695
rect 1685 22593 1719 22627
rect 2145 22593 2179 22627
rect 2789 22593 2823 22627
rect 24409 22593 24443 22627
rect 26249 22593 26283 22627
rect 27445 22593 27479 22627
rect 28641 22593 28675 22627
rect 31309 22593 31343 22627
rect 34989 22593 35023 22627
rect 35817 22593 35851 22627
rect 37468 22593 37502 22627
rect 37565 22593 37599 22627
rect 37785 22593 37819 22627
rect 37933 22593 37967 22627
rect 27261 22525 27295 22559
rect 28733 22525 28767 22559
rect 28825 22525 28859 22559
rect 32137 22525 32171 22559
rect 32597 22525 32631 22559
rect 33701 22525 33735 22559
rect 34805 22525 34839 22559
rect 28273 22457 28307 22491
rect 32229 22457 32263 22491
rect 34069 22457 34103 22491
rect 35357 22457 35391 22491
rect 37289 22457 37323 22491
rect 1501 22389 1535 22423
rect 3433 22389 3467 22423
rect 22753 22389 22787 22423
rect 24041 22389 24075 22423
rect 25697 22389 25731 22423
rect 27813 22389 27847 22423
rect 36001 22389 36035 22423
rect 34069 22185 34103 22219
rect 35173 22185 35207 22219
rect 37197 22185 37231 22219
rect 25881 22117 25915 22151
rect 28365 22117 28399 22151
rect 34989 22117 35023 22151
rect 2145 22049 2179 22083
rect 25513 22049 25547 22083
rect 28273 22049 28307 22083
rect 35817 22049 35851 22083
rect 22569 21981 22603 22015
rect 22845 21981 22879 22015
rect 23029 21981 23063 22015
rect 24409 21981 24443 22015
rect 24593 21981 24627 22015
rect 26433 21981 26467 22015
rect 32873 21981 32907 22015
rect 33517 21981 33551 22015
rect 34713 21981 34747 22015
rect 36084 21981 36118 22015
rect 37841 21981 37875 22015
rect 1869 21913 1903 21947
rect 2697 21913 2731 21947
rect 22727 21913 22761 21947
rect 22937 21913 22971 21947
rect 23673 21913 23707 21947
rect 26678 21913 26712 21947
rect 28733 21913 28767 21947
rect 30849 21913 30883 21947
rect 32628 21913 32662 21947
rect 23213 21845 23247 21879
rect 24777 21845 24811 21879
rect 25973 21845 26007 21879
rect 27813 21845 27847 21879
rect 30941 21845 30975 21879
rect 31493 21845 31527 21879
rect 33333 21845 33367 21879
rect 38025 21845 38059 21879
rect 26433 21641 26467 21675
rect 29837 21641 29871 21675
rect 32137 21641 32171 21675
rect 32597 21641 32631 21675
rect 34621 21641 34655 21675
rect 13829 21573 13863 21607
rect 24685 21573 24719 21607
rect 28181 21573 28215 21607
rect 28365 21573 28399 21607
rect 35081 21573 35115 21607
rect 36369 21573 36403 21607
rect 37657 21573 37691 21607
rect 1409 21505 1443 21539
rect 2053 21505 2087 21539
rect 14473 21505 14507 21539
rect 14749 21505 14783 21539
rect 18133 21505 18167 21539
rect 24501 21505 24535 21539
rect 26249 21505 26283 21539
rect 27353 21505 27387 21539
rect 29929 21505 29963 21539
rect 32505 21505 32539 21539
rect 33333 21505 33367 21539
rect 34069 21505 34103 21539
rect 34989 21505 35023 21539
rect 36272 21505 36306 21539
rect 36461 21505 36495 21539
rect 36644 21505 36678 21539
rect 36737 21505 36771 21539
rect 37427 21505 37461 21539
rect 37565 21505 37599 21539
rect 37840 21505 37874 21539
rect 37933 21505 37967 21539
rect 17877 21437 17911 21471
rect 27445 21437 27479 21471
rect 27537 21437 27571 21471
rect 31125 21437 31159 21471
rect 32781 21437 32815 21471
rect 35173 21437 35207 21471
rect 26985 21369 27019 21403
rect 31493 21369 31527 21403
rect 1593 21301 1627 21335
rect 14289 21301 14323 21335
rect 14657 21301 14691 21335
rect 17325 21301 17359 21335
rect 19257 21301 19291 21335
rect 24317 21301 24351 21335
rect 25237 21301 25271 21335
rect 31585 21301 31619 21335
rect 36093 21301 36127 21335
rect 37289 21301 37323 21335
rect 31953 21097 31987 21131
rect 34161 21097 34195 21131
rect 17877 21029 17911 21063
rect 26801 21029 26835 21063
rect 36829 21029 36863 21063
rect 2789 20961 2823 20995
rect 32597 20961 32631 20995
rect 35357 20961 35391 20995
rect 1685 20893 1719 20927
rect 14657 20893 14691 20927
rect 14933 20893 14967 20927
rect 15117 20893 15151 20927
rect 17785 20893 17819 20927
rect 18061 20893 18095 20927
rect 24777 20893 24811 20927
rect 32413 20893 32447 20927
rect 35081 20893 35115 20927
rect 36001 20893 36035 20927
rect 37008 20893 37042 20927
rect 37105 20893 37139 20927
rect 37380 20893 37414 20927
rect 37473 20893 37507 20927
rect 38117 20893 38151 20927
rect 24593 20825 24627 20859
rect 32321 20825 32355 20859
rect 37197 20825 37231 20859
rect 1501 20757 1535 20791
rect 2145 20757 2179 20791
rect 14473 20757 14507 20791
rect 15669 20757 15703 20791
rect 17233 20757 17267 20791
rect 18245 20757 18279 20791
rect 24409 20757 24443 20791
rect 31401 20757 31435 20791
rect 34713 20757 34747 20791
rect 35173 20757 35207 20791
rect 36185 20757 36219 20791
rect 37933 20757 37967 20791
rect 13553 20553 13587 20587
rect 15393 20553 15427 20587
rect 17417 20553 17451 20587
rect 19809 20553 19843 20587
rect 23489 20553 23523 20587
rect 23581 20553 23615 20587
rect 25237 20553 25271 20587
rect 27169 20553 27203 20587
rect 36737 20553 36771 20587
rect 14280 20485 14314 20519
rect 18144 20485 18178 20519
rect 22937 20485 22971 20519
rect 24685 20485 24719 20519
rect 37565 20485 37599 20519
rect 1869 20417 1903 20451
rect 2697 20417 2731 20451
rect 3341 20417 3375 20451
rect 17233 20417 17267 20451
rect 19993 20417 20027 20451
rect 20269 20417 20303 20451
rect 20453 20417 20487 20451
rect 23121 20417 23155 20451
rect 23673 20417 23707 20451
rect 24501 20417 24535 20451
rect 26985 20417 27019 20451
rect 30674 20417 30708 20451
rect 32781 20417 32815 20451
rect 37427 20417 37461 20451
rect 37657 20417 37691 20451
rect 37785 20417 37819 20451
rect 37933 20417 37967 20451
rect 14013 20349 14047 20383
rect 16129 20349 16163 20383
rect 16957 20349 16991 20383
rect 17877 20349 17911 20383
rect 23380 20349 23414 20383
rect 30941 20349 30975 20383
rect 33057 20349 33091 20383
rect 2145 20281 2179 20315
rect 29561 20281 29595 20315
rect 2881 20213 2915 20247
rect 17049 20213 17083 20247
rect 19257 20213 19291 20247
rect 24317 20213 24351 20247
rect 27721 20213 27755 20247
rect 37289 20213 37323 20247
rect 12909 20009 12943 20043
rect 16681 20009 16715 20043
rect 18061 20009 18095 20043
rect 23029 20009 23063 20043
rect 24593 20009 24627 20043
rect 29745 20009 29779 20043
rect 32965 20009 32999 20043
rect 27537 19941 27571 19975
rect 38025 19941 38059 19975
rect 22477 19873 22511 19907
rect 22569 19873 22603 19907
rect 23765 19873 23799 19907
rect 28181 19873 28215 19907
rect 1685 19805 1719 19839
rect 13093 19805 13127 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 15853 19805 15887 19839
rect 16497 19805 16531 19839
rect 16773 19805 16807 19839
rect 18245 19805 18279 19839
rect 18521 19805 18555 19839
rect 18705 19805 18739 19839
rect 22273 19805 22307 19839
rect 23469 19805 23503 19839
rect 24409 19805 24443 19839
rect 28365 19805 28399 19839
rect 28457 19805 28491 19839
rect 29561 19805 29595 19839
rect 37841 19805 37875 19839
rect 2697 19737 2731 19771
rect 15608 19737 15642 19771
rect 21833 19737 21867 19771
rect 22017 19737 22051 19771
rect 23213 19737 23247 19771
rect 23673 19737 23707 19771
rect 33057 19737 33091 19771
rect 1501 19669 1535 19703
rect 2145 19669 2179 19703
rect 3893 19669 3927 19703
rect 14473 19669 14507 19703
rect 16313 19669 16347 19703
rect 17509 19669 17543 19703
rect 19717 19669 19751 19703
rect 22385 19669 22419 19703
rect 23581 19669 23615 19703
rect 28825 19669 28859 19703
rect 32413 19669 32447 19703
rect 36277 19669 36311 19703
rect 37381 19669 37415 19703
rect 3065 19465 3099 19499
rect 15301 19465 15335 19499
rect 23489 19465 23523 19499
rect 29101 19465 29135 19499
rect 27629 19397 27663 19431
rect 1869 19329 1903 19363
rect 2697 19329 2731 19363
rect 3525 19329 3559 19363
rect 3709 19329 3743 19363
rect 13921 19329 13955 19363
rect 14188 19329 14222 19363
rect 20729 19329 20763 19363
rect 21005 19329 21039 19363
rect 21189 19329 21223 19363
rect 23121 19329 23155 19363
rect 23581 19329 23615 19363
rect 23673 19329 23707 19363
rect 27813 19329 27847 19363
rect 36461 19329 36495 19363
rect 37841 19329 37875 19363
rect 2789 19261 2823 19295
rect 19625 19261 19659 19295
rect 20913 19261 20947 19295
rect 23380 19261 23414 19295
rect 28641 19261 28675 19295
rect 36737 19261 36771 19295
rect 2145 19193 2179 19227
rect 18889 19193 18923 19227
rect 20821 19193 20855 19227
rect 22937 19193 22971 19227
rect 28917 19193 28951 19227
rect 2881 19125 2915 19159
rect 3893 19125 3927 19159
rect 16037 19125 16071 19159
rect 16681 19125 16715 19159
rect 27169 19125 27203 19159
rect 34805 19125 34839 19159
rect 35449 19125 35483 19159
rect 37289 19125 37323 19159
rect 38025 19125 38059 19159
rect 2789 18921 2823 18955
rect 3801 18921 3835 18955
rect 15393 18921 15427 18955
rect 19993 18921 20027 18955
rect 20177 18921 20211 18955
rect 21189 18921 21223 18955
rect 22201 18921 22235 18955
rect 20821 18853 20855 18887
rect 21833 18853 21867 18887
rect 2789 18785 2823 18819
rect 3893 18785 3927 18819
rect 35909 18785 35943 18819
rect 37197 18785 37231 18819
rect 1409 18717 1443 18751
rect 2881 18717 2915 18751
rect 3801 18717 3835 18751
rect 4077 18717 4111 18751
rect 14289 18717 14323 18751
rect 14749 18717 14783 18751
rect 14933 18717 14967 18751
rect 15209 18717 15243 18751
rect 19901 18717 19935 18751
rect 20033 18717 20067 18751
rect 20729 18717 20763 18751
rect 20913 18717 20947 18751
rect 21005 18717 21039 18751
rect 21741 18717 21775 18751
rect 21925 18717 21959 18751
rect 22017 18717 22051 18751
rect 27721 18717 27755 18751
rect 28181 18717 28215 18751
rect 28457 18717 28491 18751
rect 32413 18717 32447 18751
rect 36185 18717 36219 18751
rect 37473 18717 37507 18751
rect 38117 18717 38151 18751
rect 2421 18649 2455 18683
rect 13369 18649 13403 18683
rect 13553 18649 13587 18683
rect 19717 18649 19751 18683
rect 24869 18649 24903 18683
rect 25053 18649 25087 18683
rect 1593 18581 1627 18615
rect 3065 18581 3099 18615
rect 4261 18581 4295 18615
rect 11989 18581 12023 18615
rect 26893 18581 26927 18615
rect 31861 18581 31895 18615
rect 32597 18581 32631 18615
rect 34897 18581 34931 18615
rect 37933 18581 37967 18615
rect 2697 18377 2731 18411
rect 13461 18377 13495 18411
rect 14197 18377 14231 18411
rect 20269 18377 20303 18411
rect 21281 18377 21315 18411
rect 22293 18377 22327 18411
rect 2237 18309 2271 18343
rect 18797 18309 18831 18343
rect 25697 18309 25731 18343
rect 25881 18309 25915 18343
rect 1869 18241 1903 18275
rect 3249 18241 3283 18275
rect 3341 18241 3375 18275
rect 3525 18241 3559 18275
rect 9229 18241 9263 18275
rect 9505 18241 9539 18275
rect 9689 18241 9723 18275
rect 12357 18241 12391 18275
rect 13369 18241 13403 18275
rect 14381 18241 14415 18275
rect 14565 18241 14599 18275
rect 19809 18241 19843 18275
rect 20125 18241 20159 18275
rect 20821 18241 20855 18275
rect 20913 18241 20947 18275
rect 21097 18241 21131 18275
rect 21833 18241 21867 18275
rect 22109 18241 22143 18275
rect 26065 18241 26099 18275
rect 26985 18241 27019 18275
rect 30941 18241 30975 18275
rect 34529 18241 34563 18275
rect 35725 18241 35759 18275
rect 36461 18241 36495 18275
rect 37841 18241 37875 18275
rect 3985 18173 4019 18207
rect 12633 18173 12667 18207
rect 14657 18173 14691 18207
rect 19901 18173 19935 18207
rect 21925 18173 21959 18207
rect 24501 18173 24535 18207
rect 30021 18173 30055 18207
rect 30481 18173 30515 18207
rect 12449 18105 12483 18139
rect 21005 18105 21039 18139
rect 30297 18105 30331 18139
rect 35909 18105 35943 18139
rect 36645 18105 36679 18139
rect 9045 18037 9079 18071
rect 10149 18037 10183 18071
rect 10701 18037 10735 18071
rect 11713 18037 11747 18071
rect 12541 18037 12575 18071
rect 19349 18037 19383 18071
rect 19809 18037 19843 18071
rect 21833 18037 21867 18071
rect 22845 18037 22879 18071
rect 27169 18037 27203 18071
rect 31125 18037 31159 18071
rect 34713 18037 34747 18071
rect 37289 18037 37323 18071
rect 38025 18037 38059 18071
rect 1501 17833 1535 17867
rect 2329 17833 2363 17867
rect 4077 17833 4111 17867
rect 12173 17833 12207 17867
rect 14197 17833 14231 17867
rect 20637 17833 20671 17867
rect 20821 17833 20855 17867
rect 22017 17833 22051 17867
rect 28181 17833 28215 17867
rect 32413 17833 32447 17867
rect 37933 17833 37967 17867
rect 3939 17765 3973 17799
rect 7113 17765 7147 17799
rect 11437 17765 11471 17799
rect 12541 17765 12575 17799
rect 21649 17765 21683 17799
rect 24685 17765 24719 17799
rect 30481 17765 30515 17799
rect 36093 17765 36127 17799
rect 3157 17697 3191 17731
rect 4169 17697 4203 17731
rect 7205 17697 7239 17731
rect 9781 17697 9815 17731
rect 17141 17697 17175 17731
rect 20453 17697 20487 17731
rect 1685 17629 1719 17663
rect 2145 17629 2179 17663
rect 3065 17629 3099 17663
rect 3801 17629 3835 17663
rect 6837 17629 6871 17663
rect 6984 17629 7018 17663
rect 10057 17629 10091 17663
rect 11161 17629 11195 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 16865 17629 16899 17663
rect 19349 17629 19383 17663
rect 20361 17629 20395 17663
rect 20637 17629 20671 17663
rect 21557 17629 21591 17663
rect 21741 17629 21775 17663
rect 21833 17629 21867 17663
rect 24501 17629 24535 17663
rect 26065 17629 26099 17663
rect 28825 17629 28859 17663
rect 29009 17629 29043 17663
rect 31033 17629 31067 17663
rect 34713 17629 34747 17663
rect 36553 17629 36587 17663
rect 4537 17561 4571 17595
rect 7573 17561 7607 17595
rect 13185 17561 13219 17595
rect 13369 17561 13403 17595
rect 26332 17561 26366 17595
rect 29653 17561 29687 17595
rect 30113 17561 30147 17595
rect 31278 17561 31312 17595
rect 32965 17561 32999 17595
rect 33609 17561 33643 17595
rect 33793 17561 33827 17595
rect 34958 17561 34992 17595
rect 36798 17561 36832 17595
rect 6377 17493 6411 17527
rect 16129 17493 16163 17527
rect 19901 17493 19935 17527
rect 22477 17493 22511 17527
rect 25145 17493 25179 17527
rect 27445 17493 27479 17527
rect 30573 17493 30607 17527
rect 2145 17289 2179 17323
rect 3341 17289 3375 17323
rect 13369 17289 13403 17323
rect 14473 17289 14507 17323
rect 21833 17289 21867 17323
rect 23305 17289 23339 17323
rect 23765 17289 23799 17323
rect 30205 17289 30239 17323
rect 33701 17289 33735 17323
rect 35357 17289 35391 17323
rect 18521 17221 18555 17255
rect 18797 17221 18831 17255
rect 19007 17221 19041 17255
rect 25789 17221 25823 17255
rect 30665 17221 30699 17255
rect 34621 17221 34655 17255
rect 37933 17221 37967 17255
rect 1685 17153 1719 17187
rect 2789 17153 2823 17187
rect 7021 17153 7055 17187
rect 8484 17153 8518 17187
rect 10977 17153 11011 17187
rect 11805 17153 11839 17187
rect 12633 17153 12667 17187
rect 12817 17153 12851 17187
rect 13737 17153 13771 17187
rect 17141 17153 17175 17187
rect 18705 17153 18739 17187
rect 18890 17153 18924 17187
rect 19901 17153 19935 17187
rect 21097 17153 21131 17187
rect 22017 17153 22051 17187
rect 22293 17153 22327 17187
rect 22845 17153 22879 17187
rect 23029 17153 23063 17187
rect 23121 17153 23155 17187
rect 24869 17153 24903 17187
rect 25973 17153 26007 17187
rect 27721 17153 27755 17187
rect 30573 17153 30607 17187
rect 31585 17153 31619 17187
rect 34529 17153 34563 17187
rect 36461 17153 36495 17187
rect 37749 17153 37783 17187
rect 7168 17085 7202 17119
rect 7389 17085 7423 17119
rect 7757 17085 7791 17119
rect 8217 17085 8251 17119
rect 10701 17085 10735 17119
rect 13645 17085 13679 17119
rect 19165 17085 19199 17119
rect 19625 17085 19659 17119
rect 25145 17085 25179 17119
rect 27445 17085 27479 17119
rect 28365 17085 28399 17119
rect 30757 17085 30791 17119
rect 33241 17085 33275 17119
rect 34713 17085 34747 17119
rect 36737 17085 36771 17119
rect 9597 17017 9631 17051
rect 17325 17017 17359 17051
rect 22109 17017 22143 17051
rect 22201 17017 22235 17051
rect 25605 17017 25639 17051
rect 29009 17017 29043 17051
rect 33609 17017 33643 17051
rect 34161 17017 34195 17051
rect 1501 16949 1535 16983
rect 7297 16949 7331 16983
rect 12909 16949 12943 16983
rect 13553 16949 13587 16983
rect 15853 16949 15887 16983
rect 20913 16949 20947 16983
rect 22845 16949 22879 16983
rect 24685 16949 24719 16983
rect 25053 16949 25087 16983
rect 27537 16949 27571 16983
rect 27905 16949 27939 16983
rect 29653 16949 29687 16983
rect 31401 16949 31435 16983
rect 2145 16745 2179 16779
rect 6450 16745 6484 16779
rect 16221 16745 16255 16779
rect 16681 16745 16715 16779
rect 17693 16745 17727 16779
rect 22201 16745 22235 16779
rect 30481 16745 30515 16779
rect 32781 16745 32815 16779
rect 6561 16677 6595 16711
rect 21833 16677 21867 16711
rect 32321 16677 32355 16711
rect 33425 16677 33459 16711
rect 33977 16677 34011 16711
rect 6653 16609 6687 16643
rect 10977 16609 11011 16643
rect 11253 16609 11287 16643
rect 12357 16609 12391 16643
rect 14565 16609 14599 16643
rect 14841 16609 14875 16643
rect 16313 16609 16347 16643
rect 17325 16609 17359 16643
rect 17417 16609 17451 16643
rect 19809 16609 19843 16643
rect 20821 16609 20855 16643
rect 24501 16609 24535 16643
rect 27537 16609 27571 16643
rect 29929 16609 29963 16643
rect 30941 16609 30975 16643
rect 35173 16609 35207 16643
rect 35265 16609 35299 16643
rect 7941 16541 7975 16575
rect 8033 16541 8067 16575
rect 8217 16541 8251 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9413 16541 9447 16575
rect 9597 16541 9631 16575
rect 12449 16541 12483 16575
rect 13001 16541 13035 16575
rect 16221 16541 16255 16575
rect 16497 16541 16531 16575
rect 17233 16541 17267 16575
rect 17509 16541 17543 16575
rect 20085 16541 20119 16575
rect 21741 16541 21775 16575
rect 21925 16541 21959 16575
rect 22017 16541 22051 16575
rect 24768 16541 24802 16575
rect 26617 16541 26651 16575
rect 26893 16541 26927 16575
rect 27077 16541 27111 16575
rect 27804 16541 27838 16575
rect 30113 16541 30147 16575
rect 31208 16541 31242 16575
rect 35081 16541 35115 16575
rect 36001 16541 36035 16575
rect 37008 16541 37042 16575
rect 37197 16541 37231 16575
rect 37380 16541 37414 16575
rect 37473 16541 37507 16575
rect 38117 16541 38151 16575
rect 1869 16473 1903 16507
rect 2697 16473 2731 16507
rect 6285 16473 6319 16507
rect 7021 16473 7055 16507
rect 20637 16473 20671 16507
rect 37105 16473 37139 16507
rect 8401 16405 8435 16439
rect 12357 16405 12391 16439
rect 18613 16405 18647 16439
rect 22661 16405 22695 16439
rect 23305 16405 23339 16439
rect 25881 16405 25915 16439
rect 26433 16405 26467 16439
rect 28917 16405 28951 16439
rect 30021 16405 30055 16439
rect 34713 16405 34747 16439
rect 36185 16405 36219 16439
rect 36829 16405 36863 16439
rect 37933 16405 37967 16439
rect 6929 16201 6963 16235
rect 15117 16201 15151 16235
rect 21833 16201 21867 16235
rect 23305 16201 23339 16235
rect 24777 16201 24811 16235
rect 26433 16201 26467 16235
rect 27629 16201 27663 16235
rect 28181 16201 28215 16235
rect 14381 16133 14415 16167
rect 29469 16133 29503 16167
rect 1685 16065 1719 16099
rect 2145 16065 2179 16099
rect 2789 16065 2823 16099
rect 6837 16065 6871 16099
rect 8033 16065 8067 16099
rect 8300 16065 8334 16099
rect 10793 16065 10827 16099
rect 12265 16065 12299 16099
rect 13185 16065 13219 16099
rect 15209 16065 15243 16099
rect 15945 16065 15979 16099
rect 19073 16065 19107 16099
rect 21281 16065 21315 16099
rect 22017 16065 22051 16099
rect 22293 16065 22327 16099
rect 22845 16065 22879 16099
rect 23121 16065 23155 16099
rect 24961 16065 24995 16099
rect 25237 16065 25271 16099
rect 25421 16065 25455 16099
rect 25973 16065 26007 16099
rect 26249 16065 26283 16099
rect 26985 16065 27019 16099
rect 27169 16065 27203 16099
rect 27445 16065 27479 16099
rect 29285 16065 29319 16099
rect 33149 16065 33183 16099
rect 37565 16065 37599 16099
rect 7481 15997 7515 16031
rect 12909 15997 12943 16031
rect 16773 15997 16807 16031
rect 17049 15997 17083 16031
rect 18797 15997 18831 16031
rect 19533 15997 19567 16031
rect 22937 15997 22971 16031
rect 23857 15997 23891 16031
rect 33425 15997 33459 16031
rect 34529 15997 34563 16031
rect 35909 15997 35943 16031
rect 36185 15997 36219 16031
rect 37289 15997 37323 16031
rect 22109 15929 22143 15963
rect 22201 15929 22235 15963
rect 28641 15929 28675 15963
rect 34805 15929 34839 15963
rect 1501 15861 1535 15895
rect 2329 15861 2363 15895
rect 9413 15861 9447 15895
rect 9965 15861 9999 15895
rect 10885 15861 10919 15895
rect 11989 15861 12023 15895
rect 14473 15861 14507 15895
rect 15761 15861 15795 15895
rect 23121 15861 23155 15895
rect 26065 15861 26099 15895
rect 34989 15861 35023 15895
rect 2145 15657 2179 15691
rect 8953 15657 8987 15691
rect 9321 15657 9355 15691
rect 11897 15657 11931 15691
rect 13277 15657 13311 15691
rect 14749 15657 14783 15691
rect 16221 15657 16255 15691
rect 21833 15657 21867 15691
rect 23305 15657 23339 15691
rect 25145 15657 25179 15691
rect 35817 15657 35851 15691
rect 13185 15589 13219 15623
rect 16405 15589 16439 15623
rect 18705 15589 18739 15623
rect 22293 15589 22327 15623
rect 22845 15589 22879 15623
rect 10793 15521 10827 15555
rect 13001 15521 13035 15555
rect 16037 15521 16071 15555
rect 20085 15521 20119 15555
rect 20821 15521 20855 15555
rect 21925 15521 21959 15555
rect 9137 15453 9171 15487
rect 9413 15453 9447 15487
rect 12081 15453 12115 15487
rect 12449 15453 12483 15487
rect 12541 15453 12575 15487
rect 13277 15453 13311 15487
rect 14565 15453 14599 15487
rect 15485 15453 15519 15487
rect 16221 15453 16255 15487
rect 19809 15453 19843 15487
rect 20545 15453 20579 15487
rect 21833 15453 21867 15487
rect 22109 15453 22143 15487
rect 25789 15453 25823 15487
rect 35633 15453 35667 15487
rect 37008 15453 37042 15487
rect 37197 15453 37231 15487
rect 37380 15453 37414 15487
rect 37473 15453 37507 15487
rect 38117 15453 38151 15487
rect 1869 15385 1903 15419
rect 2697 15385 2731 15419
rect 12173 15385 12207 15419
rect 12265 15385 12299 15419
rect 15301 15385 15335 15419
rect 15945 15385 15979 15419
rect 17417 15385 17451 15419
rect 18521 15385 18555 15419
rect 24593 15385 24627 15419
rect 25973 15385 26007 15419
rect 27445 15385 27479 15419
rect 37105 15385 37139 15419
rect 8309 15317 8343 15351
rect 11345 15317 11379 15351
rect 17509 15317 17543 15351
rect 25605 15317 25639 15351
rect 26893 15317 26927 15351
rect 36829 15317 36863 15351
rect 37933 15317 37967 15351
rect 17325 15113 17359 15147
rect 35725 15113 35759 15147
rect 36737 15113 36771 15147
rect 38025 15113 38059 15147
rect 10977 15045 11011 15079
rect 12081 15045 12115 15079
rect 14565 15045 14599 15079
rect 18062 15045 18096 15079
rect 18291 15045 18325 15079
rect 25697 15045 25731 15079
rect 26341 15045 26375 15079
rect 37289 15045 37323 15079
rect 1409 14977 1443 15011
rect 2053 14977 2087 15011
rect 13369 14977 13403 15011
rect 15669 14977 15703 15011
rect 15945 14977 15979 15011
rect 16865 14977 16899 15011
rect 17141 14977 17175 15011
rect 17970 14967 18004 15001
rect 18153 14977 18187 15011
rect 21833 14977 21867 15011
rect 22017 14977 22051 15011
rect 22109 14977 22143 15011
rect 22845 14977 22879 15011
rect 34713 14977 34747 15011
rect 37841 14977 37875 15011
rect 15761 14909 15795 14943
rect 17049 14909 17083 14943
rect 18429 14909 18463 14943
rect 30297 14909 30331 14943
rect 12265 14841 12299 14875
rect 13185 14841 13219 14875
rect 14749 14841 14783 14875
rect 16957 14841 16991 14875
rect 18889 14841 18923 14875
rect 20729 14841 20763 14875
rect 22293 14841 22327 14875
rect 29929 14841 29963 14875
rect 1593 14773 1627 14807
rect 14013 14773 14047 14807
rect 15945 14773 15979 14807
rect 16129 14773 16163 14807
rect 17785 14773 17819 14807
rect 21189 14773 21223 14807
rect 21833 14773 21867 14807
rect 25145 14773 25179 14807
rect 29837 14773 29871 14807
rect 34897 14773 34931 14807
rect 15577 14569 15611 14603
rect 31769 14569 31803 14603
rect 34069 14569 34103 14603
rect 35173 14569 35207 14603
rect 38117 14569 38151 14603
rect 11897 14501 11931 14535
rect 13461 14501 13495 14535
rect 34989 14501 35023 14535
rect 36829 14501 36863 14535
rect 15393 14433 15427 14467
rect 16221 14433 16255 14467
rect 1685 14365 1719 14399
rect 12081 14365 12115 14399
rect 13277 14365 13311 14399
rect 15301 14365 15335 14399
rect 15577 14365 15611 14399
rect 17233 14365 17267 14399
rect 17693 14365 17727 14399
rect 18153 14365 18187 14399
rect 30389 14365 30423 14399
rect 36001 14365 36035 14399
rect 37008 14365 37042 14399
rect 37197 14365 37231 14399
rect 37380 14365 37414 14399
rect 37473 14365 37507 14399
rect 2145 14297 2179 14331
rect 12541 14297 12575 14331
rect 12725 14297 12759 14331
rect 14565 14297 14599 14331
rect 14749 14297 14783 14331
rect 17325 14297 17359 14331
rect 17417 14297 17451 14331
rect 17555 14297 17589 14331
rect 21649 14297 21683 14331
rect 30634 14297 30668 14331
rect 34713 14297 34747 14331
rect 37105 14297 37139 14331
rect 1501 14229 1535 14263
rect 9229 14229 9263 14263
rect 15761 14229 15795 14263
rect 17049 14229 17083 14263
rect 29653 14229 29687 14263
rect 36185 14229 36219 14263
rect 8953 14025 8987 14059
rect 15577 14025 15611 14059
rect 29377 14025 29411 14059
rect 29837 14025 29871 14059
rect 30205 14025 30239 14059
rect 33977 14025 34011 14059
rect 34437 14025 34471 14059
rect 36277 14025 36311 14059
rect 1685 13957 1719 13991
rect 2513 13957 2547 13991
rect 12449 13957 12483 13991
rect 12633 13957 12667 13991
rect 25881 13957 25915 13991
rect 30297 13957 30331 13991
rect 33149 13957 33183 13991
rect 34069 13957 34103 13991
rect 35142 13957 35176 13991
rect 1409 13889 1443 13923
rect 2789 13889 2823 13923
rect 7573 13889 7607 13923
rect 7840 13889 7874 13923
rect 9597 13889 9631 13923
rect 9781 13889 9815 13923
rect 9873 13889 9907 13923
rect 13369 13889 13403 13923
rect 14657 13889 14691 13923
rect 14933 13889 14967 13923
rect 15761 13889 15795 13923
rect 16037 13889 16071 13923
rect 16773 13889 16807 13923
rect 17049 13889 17083 13923
rect 26065 13889 26099 13923
rect 29193 13889 29227 13923
rect 31217 13889 31251 13923
rect 34897 13889 34931 13923
rect 37841 13889 37875 13923
rect 2605 13821 2639 13855
rect 13185 13821 13219 13855
rect 14841 13821 14875 13855
rect 16865 13821 16899 13855
rect 17877 13821 17911 13855
rect 25697 13821 25731 13855
rect 30481 13821 30515 13855
rect 33885 13821 33919 13855
rect 9413 13753 9447 13787
rect 15853 13753 15887 13787
rect 15945 13753 15979 13787
rect 16957 13753 16991 13787
rect 21833 13753 21867 13787
rect 2513 13685 2547 13719
rect 2973 13685 3007 13719
rect 10425 13685 10459 13719
rect 14933 13685 14967 13719
rect 15117 13685 15151 13719
rect 17233 13685 17267 13719
rect 31033 13685 31067 13719
rect 38025 13685 38059 13719
rect 2329 13481 2363 13515
rect 9597 13481 9631 13515
rect 12081 13481 12115 13515
rect 18705 13481 18739 13515
rect 19257 13481 19291 13515
rect 24685 13481 24719 13515
rect 28549 13481 28583 13515
rect 30205 13481 30239 13515
rect 32045 13481 32079 13515
rect 8401 13413 8435 13447
rect 26525 13413 26559 13447
rect 30021 13413 30055 13447
rect 34069 13413 34103 13447
rect 34713 13413 34747 13447
rect 4261 13345 4295 13379
rect 15577 13345 15611 13379
rect 15853 13345 15887 13379
rect 16865 13345 16899 13379
rect 21649 13345 21683 13379
rect 25237 13345 25271 13379
rect 29745 13345 29779 13379
rect 35265 13345 35299 13379
rect 1685 13277 1719 13311
rect 2145 13277 2179 13311
rect 2789 13277 2823 13311
rect 3801 13277 3835 13311
rect 4077 13277 4111 13311
rect 7021 13277 7055 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9413 13277 9447 13311
rect 10241 13277 10275 13311
rect 10517 13277 10551 13311
rect 10701 13277 10735 13311
rect 11713 13277 11747 13311
rect 12909 13277 12943 13311
rect 13093 13277 13127 13311
rect 13277 13277 13311 13311
rect 17325 13277 17359 13311
rect 19257 13277 19291 13311
rect 19349 13277 19383 13311
rect 20821 13277 20855 13311
rect 21005 13277 21039 13311
rect 21097 13277 21131 13311
rect 21557 13277 21591 13311
rect 21833 13277 21867 13311
rect 25329 13277 25363 13311
rect 25513 13277 25547 13311
rect 25697 13277 25731 13311
rect 30665 13277 30699 13311
rect 30932 13277 30966 13311
rect 35081 13277 35115 13311
rect 35909 13277 35943 13311
rect 37008 13277 37042 13311
rect 37197 13277 37231 13311
rect 37380 13277 37414 13311
rect 37473 13277 37507 13311
rect 38117 13277 38151 13311
rect 7288 13209 7322 13243
rect 10057 13209 10091 13243
rect 13461 13209 13495 13243
rect 17003 13209 17037 13243
rect 17141 13209 17175 13243
rect 17233 13209 17267 13243
rect 18061 13209 18095 13243
rect 20085 13209 20119 13243
rect 26157 13209 26191 13243
rect 26341 13209 26375 13243
rect 33701 13209 33735 13243
rect 35173 13209 35207 13243
rect 37105 13209 37139 13243
rect 1501 13141 1535 13175
rect 4353 13141 4387 13175
rect 11161 13141 11195 13175
rect 12081 13141 12115 13175
rect 12265 13141 12299 13175
rect 14197 13141 14231 13175
rect 17509 13141 17543 13175
rect 19625 13141 19659 13175
rect 20637 13141 20671 13175
rect 22017 13141 22051 13175
rect 22569 13141 22603 13175
rect 23857 13141 23891 13175
rect 34161 13141 34195 13175
rect 36829 13141 36863 13175
rect 37933 13141 37967 13175
rect 4169 12937 4203 12971
rect 12081 12937 12115 12971
rect 13645 12937 13679 12971
rect 27077 12937 27111 12971
rect 30021 12937 30055 12971
rect 30389 12937 30423 12971
rect 37381 12937 37415 12971
rect 2237 12869 2271 12903
rect 31309 12869 31343 12903
rect 1869 12801 1903 12835
rect 2697 12801 2731 12835
rect 3525 12801 3559 12835
rect 3672 12801 3706 12835
rect 7757 12801 7791 12835
rect 8024 12801 8058 12835
rect 9597 12801 9631 12835
rect 9781 12801 9815 12835
rect 9965 12801 9999 12835
rect 12265 12801 12299 12835
rect 12725 12801 12759 12835
rect 13461 12801 13495 12835
rect 14381 12801 14415 12835
rect 15669 12801 15703 12835
rect 15853 12801 15887 12835
rect 15945 12801 15979 12835
rect 16819 12801 16853 12835
rect 16957 12801 16991 12835
rect 17049 12801 17083 12835
rect 17141 12801 17175 12835
rect 18981 12801 19015 12835
rect 19901 12801 19935 12835
rect 20168 12801 20202 12835
rect 21833 12801 21867 12835
rect 22100 12801 22134 12835
rect 24308 12801 24342 12835
rect 26065 12801 26099 12835
rect 26249 12801 26283 12835
rect 26341 12801 26375 12835
rect 28825 12801 28859 12835
rect 29009 12801 29043 12835
rect 30481 12801 30515 12835
rect 33609 12801 33643 12835
rect 34437 12801 34471 12835
rect 35541 12801 35575 12835
rect 37841 12801 37875 12835
rect 3893 12733 3927 12767
rect 10057 12733 10091 12767
rect 10517 12733 10551 12767
rect 15761 12733 15795 12767
rect 16129 12733 16163 12767
rect 16681 12733 16715 12767
rect 17877 12733 17911 12767
rect 18705 12733 18739 12767
rect 24041 12733 24075 12767
rect 28273 12733 28307 12767
rect 28733 12733 28767 12767
rect 30573 12733 30607 12767
rect 34161 12733 34195 12767
rect 34345 12733 34379 12767
rect 12909 12665 12943 12699
rect 18889 12665 18923 12699
rect 3801 12597 3835 12631
rect 9137 12597 9171 12631
rect 14197 12597 14231 12631
rect 17325 12597 17359 12631
rect 18981 12597 19015 12631
rect 21281 12597 21315 12631
rect 23213 12597 23247 12631
rect 25421 12597 25455 12631
rect 25881 12597 25915 12631
rect 29193 12597 29227 12631
rect 31401 12597 31435 12631
rect 34805 12597 34839 12631
rect 35725 12597 35759 12631
rect 38025 12597 38059 12631
rect 1593 12393 1627 12427
rect 4077 12393 4111 12427
rect 4445 12393 4479 12427
rect 7941 12393 7975 12427
rect 9597 12393 9631 12427
rect 16497 12393 16531 12427
rect 19809 12393 19843 12427
rect 21741 12393 21775 12427
rect 24409 12393 24443 12427
rect 28641 12393 28675 12427
rect 37565 12393 37599 12427
rect 3939 12325 3973 12359
rect 8309 12325 8343 12359
rect 24777 12325 24811 12359
rect 34805 12325 34839 12359
rect 3157 12257 3191 12291
rect 4169 12257 4203 12291
rect 13461 12257 13495 12291
rect 20729 12257 20763 12291
rect 25421 12257 25455 12291
rect 34713 12257 34747 12291
rect 1409 12189 1443 12223
rect 2053 12189 2087 12223
rect 3065 12189 3099 12223
rect 8125 12189 8159 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 9413 12189 9447 12223
rect 13185 12189 13219 12223
rect 20453 12189 20487 12223
rect 21925 12189 21959 12223
rect 22201 12189 22235 12223
rect 22385 12189 22419 12223
rect 24593 12189 24627 12223
rect 24869 12189 24903 12223
rect 25688 12189 25722 12223
rect 27261 12189 27295 12223
rect 29561 12189 29595 12223
rect 29817 12189 29851 12223
rect 33977 12189 34011 12223
rect 35725 12189 35759 12223
rect 36185 12189 36219 12223
rect 3801 12121 3835 12155
rect 16405 12121 16439 12155
rect 23857 12121 23891 12155
rect 27506 12121 27540 12155
rect 35173 12121 35207 12155
rect 36430 12121 36464 12155
rect 7389 12053 7423 12087
rect 18613 12053 18647 12087
rect 26801 12053 26835 12087
rect 30941 12053 30975 12087
rect 34161 12053 34195 12087
rect 13277 11849 13311 11883
rect 14013 11849 14047 11883
rect 21833 11849 21867 11883
rect 24409 11849 24443 11883
rect 26157 11849 26191 11883
rect 28549 11849 28583 11883
rect 29101 11849 29135 11883
rect 13369 11781 13403 11815
rect 34774 11781 34808 11815
rect 37565 11781 37599 11815
rect 1685 11713 1719 11747
rect 9321 11713 9355 11747
rect 12449 11713 12483 11747
rect 22017 11713 22051 11747
rect 22293 11713 22327 11747
rect 22477 11713 22511 11747
rect 24593 11713 24627 11747
rect 24869 11713 24903 11747
rect 25053 11713 25087 11747
rect 25513 11713 25547 11747
rect 25697 11713 25731 11747
rect 25973 11713 26007 11747
rect 29285 11713 29319 11747
rect 29561 11713 29595 11747
rect 29745 11713 29779 11747
rect 30757 11713 30791 11747
rect 32597 11713 32631 11747
rect 32781 11713 32815 11747
rect 34069 11713 34103 11747
rect 34529 11713 34563 11747
rect 37289 11713 37323 11747
rect 37382 11713 37416 11747
rect 37657 11713 37691 11747
rect 37754 11713 37788 11747
rect 20453 11645 20487 11679
rect 20729 11645 20763 11679
rect 1501 11577 1535 11611
rect 2605 11577 2639 11611
rect 9873 11577 9907 11611
rect 35909 11577 35943 11611
rect 3065 11509 3099 11543
rect 9137 11509 9171 11543
rect 12265 11509 12299 11543
rect 30205 11509 30239 11543
rect 37933 11509 37967 11543
rect 2145 11305 2179 11339
rect 10149 11305 10183 11339
rect 12725 11305 12759 11339
rect 16313 11305 16347 11339
rect 16773 11305 16807 11339
rect 26065 11305 26099 11339
rect 36645 11305 36679 11339
rect 38025 11305 38059 11339
rect 12449 11237 12483 11271
rect 14841 11237 14875 11271
rect 25605 11237 25639 11271
rect 37289 11237 37323 11271
rect 14749 11169 14783 11203
rect 29561 11169 29595 11203
rect 30665 11169 30699 11203
rect 1869 11101 1903 11135
rect 2881 11101 2915 11135
rect 9505 11101 9539 11135
rect 12633 11101 12667 11135
rect 12725 11101 12759 11135
rect 12909 11101 12943 11135
rect 14657 11101 14691 11135
rect 14933 11101 14967 11135
rect 24961 11101 24995 11135
rect 25145 11101 25179 11135
rect 25421 11101 25455 11135
rect 30481 11101 30515 11135
rect 36001 11101 36035 11135
rect 36461 11101 36495 11135
rect 37105 11101 37139 11135
rect 37841 11101 37875 11135
rect 30573 11033 30607 11067
rect 2697 10965 2731 10999
rect 9413 10965 9447 10999
rect 15117 10965 15151 10999
rect 30113 10965 30147 10999
rect 9505 10761 9539 10795
rect 25697 10761 25731 10795
rect 37381 10761 37415 10795
rect 8861 10693 8895 10727
rect 11989 10693 12023 10727
rect 13553 10693 13587 10727
rect 15761 10693 15795 10727
rect 15853 10693 15887 10727
rect 29837 10693 29871 10727
rect 1685 10625 1719 10659
rect 11713 10625 11747 10659
rect 12817 10625 12851 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 15485 10625 15519 10659
rect 15623 10625 15657 10659
rect 15945 10625 15979 10659
rect 16865 10625 16899 10659
rect 19073 10625 19107 10659
rect 19257 10625 19291 10659
rect 20085 10625 20119 10659
rect 25237 10625 25271 10659
rect 37841 10625 37875 10659
rect 11897 10557 11931 10591
rect 17049 10557 17083 10591
rect 17141 10557 17175 10591
rect 17969 10489 18003 10523
rect 29653 10489 29687 10523
rect 1501 10421 1535 10455
rect 2145 10421 2179 10455
rect 2789 10421 2823 10455
rect 3249 10421 3283 10455
rect 8769 10421 8803 10455
rect 11529 10421 11563 10455
rect 11989 10421 12023 10455
rect 16129 10421 16163 10455
rect 16681 10421 16715 10455
rect 19901 10421 19935 10455
rect 22661 10421 22695 10455
rect 38025 10421 38059 10455
rect 2145 10217 2179 10251
rect 10701 10217 10735 10251
rect 11621 10217 11655 10251
rect 12725 10217 12759 10251
rect 14105 10217 14139 10251
rect 17601 10217 17635 10251
rect 22569 10217 22603 10251
rect 23765 10217 23799 10251
rect 27629 10217 27663 10251
rect 32597 10217 32631 10251
rect 35817 10217 35851 10251
rect 36277 10217 36311 10251
rect 18429 10149 18463 10183
rect 19257 10149 19291 10183
rect 30297 10149 30331 10183
rect 10609 10081 10643 10115
rect 11529 10081 11563 10115
rect 15853 10081 15887 10115
rect 18521 10081 18555 10115
rect 19993 10081 20027 10115
rect 21281 10081 21315 10115
rect 25513 10081 25547 10115
rect 37013 10081 37047 10115
rect 1869 10013 1903 10047
rect 7757 10013 7791 10047
rect 8033 10013 8067 10047
rect 8217 10013 8251 10047
rect 10701 10013 10735 10047
rect 11621 10013 11655 10047
rect 12909 10013 12943 10047
rect 13553 10013 13587 10047
rect 16129 10013 16163 10047
rect 16957 10013 16991 10047
rect 17141 10013 17175 10047
rect 17417 10013 17451 10047
rect 18245 10013 18279 10047
rect 19441 10013 19475 10047
rect 20269 10013 20303 10047
rect 24409 10013 24443 10047
rect 25605 10013 25639 10047
rect 25789 10013 25823 10047
rect 27813 10013 27847 10047
rect 31217 10013 31251 10047
rect 37289 10013 37323 10047
rect 10425 9945 10459 9979
rect 11345 9945 11379 9979
rect 26433 9945 26467 9979
rect 27997 9945 28031 9979
rect 30021 9945 30055 9979
rect 31462 9945 31496 9979
rect 2789 9877 2823 9911
rect 7573 9877 7607 9911
rect 10885 9877 10919 9911
rect 11805 9877 11839 9911
rect 13369 9877 13403 9911
rect 18061 9877 18095 9911
rect 22109 9877 22143 9911
rect 23121 9877 23155 9911
rect 24593 9877 24627 9911
rect 25973 9877 26007 9911
rect 30481 9877 30515 9911
rect 22385 9673 22419 9707
rect 23949 9673 23983 9707
rect 26985 9673 27019 9707
rect 30849 9673 30883 9707
rect 10517 9605 10551 9639
rect 14105 9605 14139 9639
rect 17684 9605 17718 9639
rect 22293 9605 22327 9639
rect 24685 9605 24719 9639
rect 27721 9605 27755 9639
rect 28365 9605 28399 9639
rect 31585 9605 31619 9639
rect 33149 9605 33183 9639
rect 33701 9605 33735 9639
rect 1409 9537 1443 9571
rect 2053 9537 2087 9571
rect 3045 9537 3079 9571
rect 4813 9537 4847 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 7205 9537 7239 9571
rect 7472 9537 7506 9571
rect 9229 9537 9263 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 10793 9537 10827 9571
rect 12081 9537 12115 9571
rect 12393 9537 12427 9571
rect 13093 9537 13127 9571
rect 13185 9537 13219 9571
rect 13369 9537 13403 9571
rect 19441 9537 19475 9571
rect 20453 9537 20487 9571
rect 23213 9537 23247 9571
rect 23397 9537 23431 9571
rect 24133 9537 24167 9571
rect 25513 9537 25547 9571
rect 25789 9537 25823 9571
rect 30665 9537 30699 9571
rect 31401 9537 31435 9571
rect 35173 9537 35207 9571
rect 36737 9537 36771 9571
rect 37289 9537 37323 9571
rect 2789 9469 2823 9503
rect 10609 9469 10643 9503
rect 12265 9469 12299 9503
rect 13921 9469 13955 9503
rect 17417 9469 17451 9503
rect 19625 9469 19659 9503
rect 19717 9469 19751 9503
rect 22937 9469 22971 9503
rect 37565 9469 37599 9503
rect 4169 9401 4203 9435
rect 8585 9401 8619 9435
rect 10977 9401 11011 9435
rect 12173 9401 12207 9435
rect 13277 9401 13311 9435
rect 1593 9333 1627 9367
rect 2237 9333 2271 9367
rect 4629 9333 4663 9367
rect 5825 9333 5859 9367
rect 9045 9333 9079 9367
rect 10793 9333 10827 9367
rect 11897 9333 11931 9367
rect 12909 9333 12943 9367
rect 18797 9333 18831 9367
rect 19257 9333 19291 9367
rect 20269 9333 20303 9367
rect 23029 9333 23063 9367
rect 25605 9333 25639 9367
rect 25973 9333 26007 9367
rect 28457 9333 28491 9367
rect 33793 9333 33827 9367
rect 35357 9333 35391 9367
rect 36507 9333 36541 9367
rect 2513 9129 2547 9163
rect 2973 9129 3007 9163
rect 22753 9129 22787 9163
rect 25513 9129 25547 9163
rect 27353 9129 27387 9163
rect 32321 9129 32355 9163
rect 11069 9061 11103 9095
rect 12173 9061 12207 9095
rect 18429 9061 18463 9095
rect 19257 9061 19291 9095
rect 20453 9061 20487 9095
rect 34989 9061 35023 9095
rect 2697 8993 2731 9027
rect 6653 8993 6687 9027
rect 11161 8993 11195 9027
rect 12265 8993 12299 9027
rect 14933 8993 14967 9027
rect 21373 8993 21407 9027
rect 22293 8993 22327 9027
rect 33149 8993 33183 9027
rect 2513 8925 2547 8959
rect 2789 8925 2823 8959
rect 3801 8925 3835 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 12081 8925 12115 8959
rect 12357 8925 12391 8959
rect 14657 8925 14691 8959
rect 16874 8925 16908 8959
rect 17141 8925 17175 8959
rect 17785 8925 17819 8959
rect 17969 8925 18003 8959
rect 18245 8925 18279 8959
rect 19441 8925 19475 8959
rect 19717 8925 19751 8959
rect 19901 8925 19935 8959
rect 22017 8925 22051 8959
rect 22201 8925 22235 8959
rect 22937 8925 22971 8959
rect 23213 8925 23247 8959
rect 23397 8925 23431 8959
rect 24869 8925 24903 8959
rect 25053 8925 25087 8959
rect 25329 8925 25363 8959
rect 25973 8925 26007 8959
rect 26240 8925 26274 8959
rect 30665 8925 30699 8959
rect 31677 8925 31711 8959
rect 33425 8925 33459 8959
rect 34713 8925 34747 8959
rect 36093 8925 36127 8959
rect 38117 8925 38151 8959
rect 1685 8857 1719 8891
rect 2053 8857 2087 8891
rect 4068 8857 4102 8891
rect 6920 8857 6954 8891
rect 10333 8857 10367 8891
rect 13001 8857 13035 8891
rect 36360 8857 36394 8891
rect 5181 8789 5215 8823
rect 8033 8789 8067 8823
rect 10241 8789 10275 8823
rect 11437 8789 11471 8823
rect 11897 8789 11931 8823
rect 15761 8789 15795 8823
rect 21833 8789 21867 8823
rect 27997 8789 28031 8823
rect 29745 8789 29779 8823
rect 30849 8789 30883 8823
rect 31585 8789 31619 8823
rect 35173 8789 35207 8823
rect 37473 8789 37507 8823
rect 37933 8789 37967 8823
rect 1501 8585 1535 8619
rect 4077 8585 4111 8619
rect 5641 8585 5675 8619
rect 7113 8585 7147 8619
rect 8033 8585 8067 8619
rect 25789 8585 25823 8619
rect 27353 8585 27387 8619
rect 30297 8585 30331 8619
rect 34437 8585 34471 8619
rect 36737 8585 36771 8619
rect 37381 8585 37415 8619
rect 9137 8517 9171 8551
rect 12174 8517 12208 8551
rect 12265 8517 12299 8551
rect 12403 8517 12437 8551
rect 14289 8517 14323 8551
rect 21925 8517 21959 8551
rect 23296 8517 23330 8551
rect 27537 8517 27571 8551
rect 30389 8517 30423 8551
rect 37749 8517 37783 8551
rect 1685 8449 1719 8483
rect 2697 8449 2731 8483
rect 2964 8449 2998 8483
rect 4721 8449 4755 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 12081 8449 12115 8483
rect 12541 8449 12575 8483
rect 13093 8449 13127 8483
rect 13369 8449 13403 8483
rect 14105 8449 14139 8483
rect 18797 8449 18831 8483
rect 19064 8449 19098 8483
rect 22134 8449 22168 8483
rect 22385 8449 22419 8483
rect 22486 8449 22520 8483
rect 25145 8449 25179 8483
rect 25329 8449 25363 8483
rect 25605 8449 25639 8483
rect 27721 8449 27755 8483
rect 34529 8449 34563 8483
rect 35357 8449 35391 8483
rect 35613 8449 35647 8483
rect 37560 8449 37594 8483
rect 37657 8449 37691 8483
rect 37932 8449 37966 8483
rect 38025 8449 38059 8483
rect 6653 8381 6687 8415
rect 7573 8381 7607 8415
rect 8493 8381 8527 8415
rect 13277 8381 13311 8415
rect 23029 8381 23063 8415
rect 28181 8381 28215 8415
rect 28457 8381 28491 8415
rect 30481 8381 30515 8415
rect 34345 8381 34379 8415
rect 2145 8313 2179 8347
rect 4537 8313 4571 8347
rect 8953 8313 8987 8347
rect 13185 8313 13219 8347
rect 13553 8313 13587 8347
rect 20177 8313 20211 8347
rect 21281 8313 21315 8347
rect 24409 8313 24443 8347
rect 33609 8313 33643 8347
rect 11897 8245 11931 8279
rect 29929 8245 29963 8279
rect 34897 8245 34931 8279
rect 2789 8041 2823 8075
rect 12633 8041 12667 8075
rect 13093 8041 13127 8075
rect 16589 8041 16623 8075
rect 32873 8041 32907 8075
rect 36093 8041 36127 8075
rect 38025 8041 38059 8075
rect 5365 7973 5399 8007
rect 27997 7973 28031 8007
rect 28641 7973 28675 8007
rect 30113 7973 30147 8007
rect 30297 7973 30331 8007
rect 32321 7973 32355 8007
rect 25973 7905 26007 7939
rect 29837 7905 29871 7939
rect 34069 7905 34103 7939
rect 35265 7905 35299 7939
rect 37381 7905 37415 7939
rect 1685 7837 1719 7871
rect 2973 7837 3007 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 4353 7837 4387 7871
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 12633 7837 12667 7871
rect 12817 7837 12851 7871
rect 12909 7837 12943 7871
rect 21557 7837 21591 7871
rect 26229 7837 26263 7871
rect 27813 7837 27847 7871
rect 30941 7837 30975 7871
rect 31197 7837 31231 7871
rect 35081 7837 35115 7871
rect 35909 7837 35943 7871
rect 37841 7837 37875 7871
rect 9321 7769 9355 7803
rect 9505 7769 9539 7803
rect 10149 7769 10183 7803
rect 21824 7769 21858 7803
rect 1501 7701 1535 7735
rect 2237 7701 2271 7735
rect 4169 7701 4203 7735
rect 7941 7701 7975 7735
rect 22937 7701 22971 7735
rect 23397 7701 23431 7735
rect 27353 7701 27387 7735
rect 34713 7701 34747 7735
rect 35173 7701 35207 7735
rect 3341 7497 3375 7531
rect 4261 7497 4295 7531
rect 6929 7497 6963 7531
rect 22661 7497 22695 7531
rect 34897 7497 34931 7531
rect 35357 7497 35391 7531
rect 36277 7497 36311 7531
rect 6377 7429 6411 7463
rect 29285 7429 29319 7463
rect 30205 7429 30239 7463
rect 34437 7429 34471 7463
rect 37657 7429 37691 7463
rect 37749 7429 37783 7463
rect 1409 7361 1443 7395
rect 3525 7361 3559 7395
rect 3801 7361 3835 7395
rect 4445 7361 4479 7395
rect 4629 7361 4663 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 9781 7361 9815 7395
rect 15209 7361 15243 7395
rect 15853 7361 15887 7395
rect 16865 7361 16899 7395
rect 17141 7361 17175 7395
rect 19533 7361 19567 7395
rect 19993 7361 20027 7395
rect 27721 7361 27755 7395
rect 27905 7361 27939 7395
rect 31033 7361 31067 7395
rect 37560 7361 37594 7395
rect 37877 7361 37911 7395
rect 38025 7361 38059 7395
rect 2881 7293 2915 7327
rect 4721 7293 4755 7327
rect 7941 7293 7975 7327
rect 9505 7293 9539 7327
rect 16129 7293 16163 7327
rect 19257 7293 19291 7327
rect 30297 7293 30331 7327
rect 30389 7293 30423 7327
rect 1593 7225 1627 7259
rect 16037 7225 16071 7259
rect 17049 7225 17083 7259
rect 34805 7225 34839 7259
rect 37381 7225 37415 7259
rect 2237 7157 2271 7191
rect 3709 7157 3743 7191
rect 5273 7157 5307 7191
rect 5733 7157 5767 7191
rect 7481 7157 7515 7191
rect 13277 7157 13311 7191
rect 15669 7157 15703 7191
rect 16681 7157 16715 7191
rect 27537 7157 27571 7191
rect 29837 7157 29871 7191
rect 31217 7157 31251 7191
rect 12265 6953 12299 6987
rect 15945 6953 15979 6987
rect 17049 6953 17083 6987
rect 32781 6953 32815 6987
rect 36645 6953 36679 6987
rect 38025 6953 38059 6987
rect 30113 6885 30147 6919
rect 6285 6817 6319 6851
rect 7021 6817 7055 6851
rect 11621 6817 11655 6851
rect 12817 6817 12851 6851
rect 23305 6817 23339 6851
rect 24501 6817 24535 6851
rect 29837 6817 29871 6851
rect 30297 6817 30331 6851
rect 30849 6817 30883 6851
rect 1685 6749 1719 6783
rect 2145 6749 2179 6783
rect 5181 6749 5215 6783
rect 7288 6749 7322 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 16129 6749 16163 6783
rect 16405 6749 16439 6783
rect 16506 6749 16540 6783
rect 17226 6743 17260 6777
rect 17509 6749 17543 6783
rect 17610 6749 17644 6783
rect 20453 6749 20487 6783
rect 23581 6749 23615 6783
rect 31116 6749 31150 6783
rect 36001 6749 36035 6783
rect 36461 6749 36495 6783
rect 37105 6749 37139 6783
rect 37841 6749 37875 6783
rect 4629 6681 4663 6715
rect 11759 6681 11793 6715
rect 11989 6681 12023 6715
rect 1501 6613 1535 6647
rect 2329 6613 2363 6647
rect 2789 6613 2823 6647
rect 4169 6613 4203 6647
rect 5733 6613 5767 6647
rect 8401 6613 8435 6647
rect 20637 6613 20671 6647
rect 32229 6613 32263 6647
rect 37289 6613 37323 6647
rect 2145 6409 2179 6443
rect 6929 6409 6963 6443
rect 7941 6409 7975 6443
rect 13185 6409 13219 6443
rect 1869 6341 1903 6375
rect 15862 6341 15896 6375
rect 19625 6341 19659 6375
rect 20269 6341 20303 6375
rect 23121 6341 23155 6375
rect 2881 6273 2915 6307
rect 8125 6273 8159 6307
rect 8401 6273 8435 6307
rect 8585 6273 8619 6307
rect 16129 6273 16163 6307
rect 21833 6273 21867 6307
rect 23305 6273 23339 6307
rect 23397 6273 23431 6307
rect 23581 6273 23615 6307
rect 23673 6273 23707 6307
rect 37841 6273 37875 6307
rect 22109 6205 22143 6239
rect 4721 6137 4755 6171
rect 34529 6137 34563 6171
rect 35909 6137 35943 6171
rect 37381 6137 37415 6171
rect 2697 6069 2731 6103
rect 3617 6069 3651 6103
rect 4261 6069 4295 6103
rect 5273 6069 5307 6103
rect 12633 6069 12667 6103
rect 13645 6069 13679 6103
rect 14749 6069 14783 6103
rect 20361 6069 20395 6103
rect 24225 6069 24259 6103
rect 35357 6069 35391 6103
rect 36369 6069 36403 6103
rect 38025 6069 38059 6103
rect 5549 5865 5583 5899
rect 6285 5865 6319 5899
rect 7389 5865 7423 5899
rect 11345 5865 11379 5899
rect 14197 5865 14231 5899
rect 19809 5865 19843 5899
rect 21649 5865 21683 5899
rect 22293 5865 22327 5899
rect 23305 5865 23339 5899
rect 24409 5865 24443 5899
rect 25789 5865 25823 5899
rect 28917 5865 28951 5899
rect 33425 5865 33459 5899
rect 36829 5865 36863 5899
rect 3801 5797 3835 5831
rect 4537 5797 4571 5831
rect 13185 5797 13219 5831
rect 36277 5797 36311 5831
rect 7481 5729 7515 5763
rect 11805 5729 11839 5763
rect 16589 5729 16623 5763
rect 26249 5729 26283 5763
rect 26525 5729 26559 5763
rect 34805 5729 34839 5763
rect 1685 5661 1719 5695
rect 2421 5661 2455 5695
rect 3157 5661 3191 5695
rect 3985 5661 4019 5695
rect 7205 5661 7239 5695
rect 10793 5661 10827 5695
rect 10885 5661 10919 5695
rect 11069 5661 11103 5695
rect 11161 5661 11195 5695
rect 12081 5661 12115 5695
rect 12265 5661 12299 5695
rect 13369 5661 13403 5695
rect 16333 5661 16367 5695
rect 19257 5661 19291 5695
rect 19349 5661 19383 5695
rect 19533 5661 19567 5695
rect 19625 5661 19659 5695
rect 22477 5661 22511 5695
rect 22569 5661 22603 5695
rect 22753 5661 22787 5695
rect 22845 5661 22879 5695
rect 23489 5661 23523 5695
rect 23581 5661 23615 5695
rect 23765 5661 23799 5695
rect 23857 5661 23891 5695
rect 24593 5661 24627 5695
rect 24685 5661 24719 5695
rect 24869 5661 24903 5695
rect 24961 5661 24995 5695
rect 35081 5661 35115 5695
rect 36093 5661 36127 5695
rect 37008 5661 37042 5695
rect 37096 5661 37130 5695
rect 37325 5661 37359 5695
rect 37473 5661 37507 5695
rect 38117 5661 38151 5695
rect 11943 5593 11977 5627
rect 12173 5593 12207 5627
rect 34989 5593 35023 5627
rect 37197 5593 37231 5627
rect 1501 5525 1535 5559
rect 2237 5525 2271 5559
rect 2973 5525 3007 5559
rect 7021 5525 7055 5559
rect 12449 5525 12483 5559
rect 15209 5525 15243 5559
rect 34161 5525 34195 5559
rect 35449 5525 35483 5559
rect 37933 5525 37967 5559
rect 3801 5321 3835 5355
rect 7389 5321 7423 5355
rect 10885 5321 10919 5355
rect 12909 5321 12943 5355
rect 14013 5321 14047 5355
rect 20545 5321 20579 5355
rect 23949 5321 23983 5355
rect 27261 5321 27295 5355
rect 28549 5321 28583 5355
rect 29377 5321 29411 5355
rect 32229 5321 32263 5355
rect 32873 5321 32907 5355
rect 12081 5253 12115 5287
rect 12173 5253 12207 5287
rect 13277 5253 13311 5287
rect 13415 5253 13449 5287
rect 15117 5253 15151 5287
rect 15301 5253 15335 5287
rect 27629 5253 27663 5287
rect 35173 5253 35207 5287
rect 37657 5253 37691 5287
rect 37749 5253 37783 5287
rect 1593 5185 1627 5219
rect 2329 5185 2363 5219
rect 2881 5185 2915 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4905 5185 4939 5219
rect 5181 5185 5215 5219
rect 5365 5185 5399 5219
rect 6653 5185 6687 5219
rect 6837 5185 6871 5219
rect 7573 5185 7607 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 10333 5185 10367 5219
rect 10425 5185 10459 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 11943 5185 11977 5219
rect 12265 5185 12299 5219
rect 13093 5185 13127 5219
rect 13185 5185 13219 5219
rect 17141 5185 17175 5219
rect 18245 5185 18279 5219
rect 19533 5185 19567 5219
rect 20729 5185 20763 5219
rect 20821 5185 20855 5219
rect 21005 5185 21039 5219
rect 21097 5185 21131 5219
rect 24133 5185 24167 5219
rect 24225 5185 24259 5219
rect 24409 5185 24443 5219
rect 24501 5185 24535 5219
rect 27445 5185 27479 5219
rect 30389 5185 30423 5219
rect 34345 5185 34379 5219
rect 34437 5185 34471 5219
rect 36093 5185 36127 5219
rect 37560 5185 37594 5219
rect 37932 5185 37966 5219
rect 38025 5185 38059 5219
rect 6929 5117 6963 5151
rect 11805 5117 11839 5151
rect 13553 5117 13587 5151
rect 17969 5117 18003 5151
rect 19257 5117 19291 5151
rect 21833 5117 21867 5151
rect 22109 5117 22143 5151
rect 28089 5117 28123 5151
rect 29469 5117 29503 5151
rect 29653 5117 29687 5151
rect 34621 5117 34655 5151
rect 35633 5117 35667 5151
rect 1777 5049 1811 5083
rect 28457 5049 28491 5083
rect 29009 5049 29043 5083
rect 33425 5049 33459 5083
rect 35449 5049 35483 5083
rect 37381 5049 37415 5083
rect 4721 4981 4755 5015
rect 6469 4981 6503 5015
rect 12449 4981 12483 5015
rect 17233 4981 17267 5015
rect 23213 4981 23247 5015
rect 25329 4981 25363 5015
rect 25789 4981 25823 5015
rect 30205 4981 30239 5015
rect 33977 4981 34011 5015
rect 36277 4981 36311 5015
rect 2789 4777 2823 4811
rect 3065 4777 3099 4811
rect 5825 4777 5859 4811
rect 8125 4777 8159 4811
rect 11069 4777 11103 4811
rect 15577 4777 15611 4811
rect 16589 4777 16623 4811
rect 17601 4777 17635 4811
rect 18613 4777 18647 4811
rect 22569 4777 22603 4811
rect 23305 4777 23339 4811
rect 24961 4777 24995 4811
rect 26801 4777 26835 4811
rect 27445 4777 27479 4811
rect 30941 4777 30975 4811
rect 37749 4777 37783 4811
rect 2145 4709 2179 4743
rect 14381 4709 14415 4743
rect 23581 4709 23615 4743
rect 25421 4709 25455 4743
rect 25697 4709 25731 4743
rect 25789 4709 25823 4743
rect 31677 4709 31711 4743
rect 33977 4709 34011 4743
rect 34713 4709 34747 4743
rect 4261 4641 4295 4675
rect 6745 4641 6779 4675
rect 19257 4641 19291 4675
rect 19533 4641 19567 4675
rect 28457 4641 28491 4675
rect 31401 4641 31435 4675
rect 32321 4641 32355 4675
rect 33609 4641 33643 4675
rect 35265 4641 35299 4675
rect 36369 4641 36403 4675
rect 2697 4573 2731 4607
rect 2881 4573 2915 4607
rect 3985 4573 4019 4607
rect 4169 4573 4203 4607
rect 4905 4573 4939 4607
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 7012 4573 7046 4607
rect 10517 4573 10551 4607
rect 10609 4573 10643 4607
rect 10793 4573 10827 4607
rect 10885 4573 10919 4607
rect 12541 4573 12575 4607
rect 12817 4573 12851 4607
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 14565 4573 14599 4607
rect 15761 4573 15795 4607
rect 15853 4573 15887 4607
rect 16037 4573 16071 4607
rect 16129 4573 16163 4607
rect 16773 4573 16807 4607
rect 16865 4573 16899 4607
rect 17049 4573 17083 4607
rect 17141 4573 17175 4607
rect 17785 4573 17819 4607
rect 17877 4573 17911 4607
rect 18061 4573 18095 4607
rect 18153 4573 18187 4607
rect 20729 4573 20763 4607
rect 21005 4573 21039 4607
rect 22017 4573 22051 4607
rect 22109 4573 22143 4607
rect 22293 4573 22327 4607
rect 22385 4573 22419 4607
rect 23489 4573 23523 4607
rect 23673 4573 23707 4607
rect 23765 4573 23799 4607
rect 24409 4573 24443 4607
rect 24501 4573 24535 4607
rect 24685 4573 24719 4607
rect 24777 4573 24811 4607
rect 25605 4573 25639 4607
rect 25881 4573 25915 4607
rect 26433 4573 26467 4607
rect 27813 4573 27847 4607
rect 28641 4573 28675 4607
rect 29561 4573 29595 4607
rect 29828 4573 29862 4607
rect 32965 4573 32999 4607
rect 36625 4573 36659 4607
rect 1869 4505 1903 4539
rect 4721 4505 4755 4539
rect 26617 4505 26651 4539
rect 27629 4505 27663 4539
rect 3801 4437 3835 4471
rect 8953 4437 8987 4471
rect 13553 4437 13587 4471
rect 14105 4437 14139 4471
rect 28549 4437 28583 4471
rect 29009 4437 29043 4471
rect 31861 4437 31895 4471
rect 33149 4437 33183 4471
rect 34069 4437 34103 4471
rect 35081 4437 35115 4471
rect 35173 4437 35207 4471
rect 13369 4233 13403 4267
rect 26341 4233 26375 4267
rect 31125 4233 31159 4267
rect 35725 4233 35759 4267
rect 3332 4165 3366 4199
rect 28365 4165 28399 4199
rect 30757 4165 30791 4199
rect 37749 4165 37783 4199
rect 1409 4097 1443 4131
rect 2605 4097 2639 4131
rect 5089 4097 5123 4131
rect 5273 4097 5307 4131
rect 7021 4097 7055 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 7665 4097 7699 4131
rect 9229 4097 9263 4131
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 10793 4097 10827 4131
rect 10977 4097 11011 4131
rect 13553 4097 13587 4131
rect 13645 4097 13679 4131
rect 13829 4097 13863 4131
rect 13921 4097 13955 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 16957 4097 16991 4131
rect 17141 4097 17175 4131
rect 17233 4097 17267 4131
rect 17969 4097 18003 4131
rect 19257 4097 19291 4131
rect 21005 4097 21039 4131
rect 22845 4097 22879 4131
rect 23029 4097 23063 4131
rect 23121 4097 23155 4131
rect 23305 4097 23339 4131
rect 23857 4097 23891 4131
rect 24041 4097 24075 4131
rect 24133 4097 24167 4131
rect 24317 4097 24351 4131
rect 24409 4097 24443 4131
rect 24869 4097 24903 4131
rect 25053 4097 25087 4131
rect 25329 4097 25363 4131
rect 29285 4097 29319 4131
rect 30665 4097 30699 4131
rect 32137 4097 32171 4131
rect 32873 4097 32907 4131
rect 34345 4097 34379 4131
rect 34612 4097 34646 4131
rect 36461 4097 36495 4131
rect 37560 4097 37594 4131
rect 37657 4097 37691 4131
rect 37877 4097 37911 4131
rect 38025 4097 38059 4131
rect 2145 4029 2179 4063
rect 3065 4029 3099 4063
rect 5365 4029 5399 4063
rect 11621 4029 11655 4063
rect 12081 4029 12115 4063
rect 12357 4029 12391 4063
rect 14381 4029 14415 4063
rect 18981 4029 19015 4063
rect 19717 4029 19751 4063
rect 19993 4029 20027 4063
rect 22385 4029 22419 4063
rect 23213 4029 23247 4063
rect 28825 4029 28859 4063
rect 30481 4029 30515 4063
rect 33425 4029 33459 4063
rect 33885 4029 33919 4063
rect 4445 3961 4479 3995
rect 25145 3961 25179 3995
rect 25237 3961 25271 3995
rect 28733 3961 28767 3995
rect 33609 3961 33643 3995
rect 37381 3961 37415 3995
rect 1593 3893 1627 3927
rect 2513 3893 2547 3927
rect 4905 3893 4939 3927
rect 6377 3893 6411 3927
rect 8217 3893 8251 3927
rect 8677 3893 8711 3927
rect 27905 3893 27939 3927
rect 29469 3893 29503 3927
rect 32321 3893 32355 3927
rect 36645 3893 36679 3927
rect 1777 3689 1811 3723
rect 2789 3689 2823 3723
rect 5181 3689 5215 3723
rect 7389 3689 7423 3723
rect 9873 3689 9907 3723
rect 10885 3689 10919 3723
rect 12909 3689 12943 3723
rect 15209 3689 15243 3723
rect 16681 3689 16715 3723
rect 17141 3689 17175 3723
rect 18153 3689 18187 3723
rect 22201 3689 22235 3723
rect 23305 3689 23339 3723
rect 23765 3689 23799 3723
rect 24961 3689 24995 3723
rect 25421 3689 25455 3723
rect 29561 3689 29595 3723
rect 30205 3689 30239 3723
rect 31033 3689 31067 3723
rect 32873 3689 32907 3723
rect 33425 3689 33459 3723
rect 36093 3689 36127 3723
rect 36553 3689 36587 3723
rect 10609 3621 10643 3655
rect 22569 3621 22603 3655
rect 24593 3621 24627 3655
rect 26985 3621 27019 3655
rect 34161 3621 34195 3655
rect 6009 3553 6043 3587
rect 10517 3553 10551 3587
rect 11529 3553 11563 3587
rect 17417 3553 17451 3587
rect 18521 3553 18555 3587
rect 19533 3553 19567 3587
rect 20637 3553 20671 3587
rect 20913 3553 20947 3587
rect 22477 3553 22511 3587
rect 24685 3553 24719 3587
rect 25697 3553 25731 3587
rect 32413 3553 32447 3587
rect 34713 3553 34747 3587
rect 2329 3485 2363 3519
rect 2973 3485 3007 3519
rect 3801 3485 3835 3519
rect 6276 3485 6310 3519
rect 7849 3485 7883 3519
rect 9413 3485 9447 3519
rect 9505 3485 9539 3519
rect 9597 3485 9631 3519
rect 9689 3485 9723 3519
rect 10425 3485 10459 3519
rect 10733 3485 10767 3519
rect 11805 3485 11839 3519
rect 17325 3485 17359 3519
rect 17509 3485 17543 3519
rect 17601 3485 17635 3519
rect 18337 3485 18371 3519
rect 18429 3485 18463 3519
rect 18613 3485 18647 3519
rect 19257 3485 19291 3519
rect 22385 3485 22419 3519
rect 22661 3485 22695 3519
rect 24501 3485 24535 3519
rect 24777 3485 24811 3519
rect 25605 3485 25639 3519
rect 25789 3485 25823 3519
rect 25881 3485 25915 3519
rect 28365 3485 28399 3519
rect 29009 3485 29043 3519
rect 32157 3485 32191 3519
rect 33977 3485 34011 3519
rect 37105 3485 37139 3519
rect 37841 3485 37875 3519
rect 1501 3417 1535 3451
rect 4068 3417 4102 3451
rect 34958 3417 34992 3451
rect 8033 3349 8067 3383
rect 13369 3349 13403 3383
rect 26433 3349 26467 3383
rect 28825 3349 28859 3383
rect 37289 3349 37323 3383
rect 38025 3349 38059 3383
rect 8033 3145 8067 3179
rect 10885 3145 10919 3179
rect 12081 3145 12115 3179
rect 14749 3145 14783 3179
rect 17233 3145 17267 3179
rect 18981 3145 19015 3179
rect 20453 3145 20487 3179
rect 21097 3145 21131 3179
rect 22753 3145 22787 3179
rect 24225 3145 24259 3179
rect 24685 3145 24719 3179
rect 26985 3145 27019 3179
rect 28181 3145 28215 3179
rect 33701 3145 33735 3179
rect 34529 3145 34563 3179
rect 35173 3145 35207 3179
rect 13829 3077 13863 3111
rect 29316 3077 29350 3111
rect 31585 3077 31619 3111
rect 1961 3009 1995 3043
rect 3249 3009 3283 3043
rect 4261 3009 4295 3043
rect 5365 3009 5399 3043
rect 6653 3009 6687 3043
rect 7389 3009 7423 3043
rect 7849 3009 7883 3043
rect 8493 3009 8527 3043
rect 9597 3009 9631 3043
rect 10425 3009 10459 3043
rect 10609 3009 10643 3043
rect 10701 3009 10735 3043
rect 11621 3009 11655 3043
rect 11805 3009 11839 3043
rect 11897 3009 11931 3043
rect 12725 3009 12759 3043
rect 13185 3009 13219 3043
rect 14565 3009 14599 3043
rect 15209 3009 15243 3043
rect 16129 3009 16163 3043
rect 17417 3009 17451 3043
rect 17601 3009 17635 3043
rect 17693 3009 17727 3043
rect 18521 3009 18555 3043
rect 18797 3009 18831 3043
rect 19533 3009 19567 3043
rect 19809 3009 19843 3043
rect 19993 3009 20027 3043
rect 20637 3009 20671 3043
rect 22937 3009 22971 3043
rect 23397 3009 23431 3043
rect 24041 3009 24075 3043
rect 24869 3009 24903 3043
rect 24961 3009 24995 3043
rect 25145 3009 25179 3043
rect 27169 3009 27203 3043
rect 27629 3009 27663 3043
rect 29561 3009 29595 3043
rect 32413 3009 32447 3043
rect 33057 3009 33091 3043
rect 33885 3009 33919 3043
rect 34345 3009 34379 3043
rect 34989 3009 35023 3043
rect 35725 3009 35759 3043
rect 36461 3009 36495 3043
rect 38117 3009 38151 3043
rect 2237 2941 2271 2975
rect 3525 2941 3559 2975
rect 18613 2941 18647 2975
rect 25697 2941 25731 2975
rect 37381 2941 37415 2975
rect 7205 2873 7239 2907
rect 10517 2873 10551 2907
rect 11713 2873 11747 2907
rect 12541 2873 12575 2907
rect 13369 2873 13403 2907
rect 17509 2873 17543 2907
rect 18705 2873 18739 2907
rect 19625 2873 19659 2907
rect 19717 2873 19751 2907
rect 21833 2873 21867 2907
rect 25053 2873 25087 2907
rect 30389 2873 30423 2907
rect 32873 2873 32907 2907
rect 36645 2873 36679 2907
rect 37933 2873 37967 2907
rect 4077 2805 4111 2839
rect 5181 2805 5215 2839
rect 6469 2805 6503 2839
rect 8677 2805 8711 2839
rect 9781 2805 9815 2839
rect 15945 2805 15979 2839
rect 16773 2805 16807 2839
rect 26249 2805 26283 2839
rect 30849 2805 30883 2839
rect 35909 2805 35943 2839
rect 3065 2601 3099 2635
rect 6469 2601 6503 2635
rect 10977 2601 11011 2635
rect 16865 2601 16899 2635
rect 10701 2533 10735 2567
rect 20821 2533 20855 2567
rect 33057 2533 33091 2567
rect 1961 2465 1995 2499
rect 28917 2465 28951 2499
rect 37289 2465 37323 2499
rect 2237 2397 2271 2431
rect 2789 2397 2823 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 5365 2397 5399 2431
rect 6653 2397 6687 2431
rect 7389 2397 7423 2431
rect 8125 2397 8159 2431
rect 9413 2397 9447 2431
rect 10517 2397 10551 2431
rect 10609 2397 10643 2431
rect 10793 2397 10827 2431
rect 11805 2397 11839 2431
rect 12541 2397 12575 2431
rect 13553 2397 13587 2431
rect 14381 2397 14415 2431
rect 15577 2397 15611 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 17601 2397 17635 2431
rect 18337 2397 18371 2431
rect 19349 2397 19383 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 22109 2397 22143 2431
rect 22569 2397 22603 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 25697 2397 25731 2431
rect 26157 2397 26191 2431
rect 27721 2397 27755 2431
rect 28181 2397 28215 2431
rect 29561 2397 29595 2431
rect 30297 2397 30331 2431
rect 31217 2397 31251 2431
rect 32137 2397 32171 2431
rect 32873 2397 32907 2431
rect 33609 2397 33643 2431
rect 34713 2397 34747 2431
rect 35633 2397 35667 2431
rect 36461 2397 36495 2431
rect 37565 2397 37599 2431
rect 9873 2329 9907 2363
rect 5181 2261 5215 2295
rect 7205 2261 7239 2295
rect 7941 2261 7975 2295
rect 9229 2261 9263 2295
rect 11621 2261 11655 2295
rect 12357 2261 12391 2295
rect 13369 2261 13403 2295
rect 14197 2261 14231 2295
rect 15393 2261 15427 2295
rect 17417 2261 17451 2295
rect 18153 2261 18187 2295
rect 19533 2261 19567 2295
rect 20269 2261 20303 2295
rect 21925 2261 21959 2295
rect 22753 2261 22787 2295
rect 23489 2261 23523 2295
rect 24593 2261 24627 2295
rect 25513 2261 25547 2295
rect 26341 2261 26375 2295
rect 27537 2261 27571 2295
rect 28365 2261 28399 2295
rect 29745 2261 29779 2295
rect 30481 2261 30515 2295
rect 31033 2261 31067 2295
rect 32321 2261 32355 2295
rect 33793 2261 33827 2295
rect 34897 2261 34931 2295
rect 35817 2261 35851 2295
rect 36645 2261 36679 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 2041 37451 2099 37457
rect 2041 37417 2053 37451
rect 2087 37448 2099 37451
rect 2774 37448 2780 37460
rect 2087 37420 2780 37448
rect 2087 37417 2099 37420
rect 2041 37411 2099 37417
rect 2774 37408 2780 37420
rect 2832 37408 2838 37460
rect 2685 37383 2743 37389
rect 2685 37349 2697 37383
rect 2731 37380 2743 37383
rect 2866 37380 2872 37392
rect 2731 37352 2872 37380
rect 2731 37349 2743 37352
rect 2685 37343 2743 37349
rect 2866 37340 2872 37352
rect 2924 37340 2930 37392
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 19426 37204 19432 37256
rect 19484 37244 19490 37256
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 19484 37216 20085 37244
rect 19484 37204 19490 37216
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 35802 37244 35808 37256
rect 35763 37216 35808 37244
rect 20073 37207 20131 37213
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 36078 37204 36084 37256
rect 36136 37244 36142 37256
rect 36449 37247 36507 37253
rect 36449 37244 36461 37247
rect 36136 37216 36461 37244
rect 36136 37204 36142 37216
rect 36449 37213 36461 37216
rect 36495 37213 36507 37247
rect 37829 37247 37887 37253
rect 37829 37244 37841 37247
rect 36449 37207 36507 37213
rect 37292 37216 37841 37244
rect 35710 37136 35716 37188
rect 35768 37176 35774 37188
rect 35768 37148 36676 37176
rect 35768 37136 35774 37148
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 35986 37108 35992 37120
rect 35947 37080 35992 37108
rect 20257 37071 20315 37077
rect 35986 37068 35992 37080
rect 36044 37068 36050 37120
rect 36648 37117 36676 37148
rect 37292 37120 37320 37216
rect 37829 37213 37841 37216
rect 37875 37213 37887 37247
rect 37829 37207 37887 37213
rect 36633 37111 36691 37117
rect 36633 37077 36645 37111
rect 36679 37077 36691 37111
rect 37274 37108 37280 37120
rect 37235 37080 37280 37108
rect 36633 37071 36691 37077
rect 37274 37068 37280 37080
rect 37332 37068 37338 37120
rect 38010 37108 38016 37120
rect 37971 37080 38016 37108
rect 38010 37068 38016 37080
rect 38068 37068 38074 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 35802 36864 35808 36916
rect 35860 36904 35866 36916
rect 36081 36907 36139 36913
rect 36081 36904 36093 36907
rect 35860 36876 36093 36904
rect 35860 36864 35866 36876
rect 36081 36873 36093 36876
rect 36127 36873 36139 36907
rect 36081 36867 36139 36873
rect 38013 36907 38071 36913
rect 38013 36873 38025 36907
rect 38059 36904 38071 36907
rect 38194 36904 38200 36916
rect 38059 36876 38200 36904
rect 38059 36873 38071 36876
rect 38013 36867 38071 36873
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1486 36768 1492 36780
rect 1443 36740 1492 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1486 36728 1492 36740
rect 1544 36728 1550 36780
rect 37369 36771 37427 36777
rect 37369 36737 37381 36771
rect 37415 36768 37427 36771
rect 37829 36771 37887 36777
rect 37829 36768 37841 36771
rect 37415 36740 37841 36768
rect 37415 36737 37427 36740
rect 37369 36731 37427 36737
rect 37829 36737 37841 36740
rect 37875 36768 37887 36771
rect 38194 36768 38200 36780
rect 37875 36740 38200 36768
rect 37875 36737 37887 36740
rect 37829 36731 37887 36737
rect 38194 36728 38200 36740
rect 38252 36728 38258 36780
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 19426 36360 19432 36372
rect 19387 36332 19432 36360
rect 19426 36320 19432 36332
rect 19484 36320 19490 36372
rect 38013 36363 38071 36369
rect 38013 36329 38025 36363
rect 38059 36360 38071 36363
rect 38102 36360 38108 36372
rect 38059 36332 38108 36360
rect 38059 36329 38071 36332
rect 38013 36323 38071 36329
rect 38102 36320 38108 36332
rect 38160 36320 38166 36372
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 18966 36116 18972 36168
rect 19024 36156 19030 36168
rect 19245 36159 19303 36165
rect 19245 36156 19257 36159
rect 19024 36128 19257 36156
rect 19024 36116 19030 36128
rect 19245 36125 19257 36128
rect 19291 36156 19303 36159
rect 19889 36159 19947 36165
rect 19889 36156 19901 36159
rect 19291 36128 19901 36156
rect 19291 36125 19303 36128
rect 19245 36119 19303 36125
rect 19889 36125 19901 36128
rect 19935 36125 19947 36159
rect 19889 36119 19947 36125
rect 36725 36159 36783 36165
rect 36725 36125 36737 36159
rect 36771 36156 36783 36159
rect 37366 36156 37372 36168
rect 36771 36128 37372 36156
rect 36771 36125 36783 36128
rect 36725 36119 36783 36125
rect 37366 36116 37372 36128
rect 37424 36116 37430 36168
rect 37829 36159 37887 36165
rect 37829 36125 37841 36159
rect 37875 36125 37887 36159
rect 37829 36119 37887 36125
rect 32122 36048 32128 36100
rect 32180 36088 32186 36100
rect 37844 36088 37872 36119
rect 32180 36060 37872 36088
rect 32180 36048 32186 36060
rect 36906 35980 36912 36032
rect 36964 36020 36970 36032
rect 37185 36023 37243 36029
rect 37185 36020 37197 36023
rect 36964 35992 37197 36020
rect 36964 35980 36970 35992
rect 37185 35989 37197 35992
rect 37231 35989 37243 36023
rect 37185 35983 37243 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 36998 35640 37004 35692
rect 37056 35680 37062 35692
rect 37829 35683 37887 35689
rect 37829 35680 37841 35683
rect 37056 35652 37841 35680
rect 37056 35640 37062 35652
rect 37829 35649 37841 35652
rect 37875 35649 37887 35683
rect 37829 35643 37887 35649
rect 1394 35476 1400 35488
rect 1355 35448 1400 35476
rect 1394 35436 1400 35448
rect 1452 35436 1458 35488
rect 38010 35476 38016 35488
rect 37971 35448 38016 35476
rect 38010 35436 38016 35448
rect 38068 35436 38074 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 37829 35071 37887 35077
rect 37829 35068 37841 35071
rect 37292 35040 37841 35068
rect 25774 34892 25780 34944
rect 25832 34932 25838 34944
rect 37292 34941 37320 35040
rect 37829 35037 37841 35040
rect 37875 35037 37887 35071
rect 37829 35031 37887 35037
rect 37277 34935 37335 34941
rect 37277 34932 37289 34935
rect 25832 34904 37289 34932
rect 25832 34892 25838 34904
rect 37277 34901 37289 34904
rect 37323 34901 37335 34935
rect 38010 34932 38016 34944
rect 37971 34904 38016 34932
rect 37277 34895 37335 34901
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1394 34456 1400 34468
rect 1355 34428 1400 34456
rect 1394 34416 1400 34428
rect 1452 34416 1458 34468
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 37461 33983 37519 33989
rect 37461 33949 37473 33983
rect 37507 33980 37519 33983
rect 38102 33980 38108 33992
rect 37507 33952 38108 33980
rect 37507 33949 37519 33952
rect 37461 33943 37519 33949
rect 38102 33940 38108 33952
rect 38160 33940 38166 33992
rect 37921 33847 37979 33853
rect 37921 33813 37933 33847
rect 37967 33844 37979 33847
rect 38286 33844 38292 33856
rect 37967 33816 38292 33844
rect 37967 33813 37979 33816
rect 37921 33807 37979 33813
rect 38286 33804 38292 33816
rect 38344 33804 38350 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 37550 33464 37556 33516
rect 37608 33504 37614 33516
rect 37829 33507 37887 33513
rect 37829 33504 37841 33507
rect 37608 33476 37841 33504
rect 37608 33464 37614 33476
rect 37829 33473 37841 33476
rect 37875 33473 37887 33507
rect 37829 33467 37887 33473
rect 38010 33300 38016 33312
rect 37971 33272 38016 33300
rect 38010 33260 38016 33272
rect 38068 33260 38074 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1394 32892 1400 32904
rect 1355 32864 1400 32892
rect 1394 32852 1400 32864
rect 1452 32852 1458 32904
rect 28350 32852 28356 32904
rect 28408 32892 28414 32904
rect 37277 32895 37335 32901
rect 37277 32892 37289 32895
rect 28408 32864 37289 32892
rect 28408 32852 28414 32864
rect 37277 32861 37289 32864
rect 37323 32892 37335 32895
rect 37829 32895 37887 32901
rect 37829 32892 37841 32895
rect 37323 32864 37841 32892
rect 37323 32861 37335 32864
rect 37277 32855 37335 32861
rect 37829 32861 37841 32864
rect 37875 32861 37887 32895
rect 37829 32855 37887 32861
rect 38010 32756 38016 32768
rect 37971 32728 38016 32756
rect 38010 32716 38016 32728
rect 38068 32716 38074 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 37461 32419 37519 32425
rect 37461 32385 37473 32419
rect 37507 32416 37519 32419
rect 38102 32416 38108 32428
rect 37507 32388 38108 32416
rect 37507 32385 37519 32388
rect 37461 32379 37519 32385
rect 38102 32376 38108 32388
rect 38160 32376 38166 32428
rect 37918 32212 37924 32224
rect 37879 32184 37924 32212
rect 37918 32172 37924 32184
rect 37976 32172 37982 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 35986 31764 35992 31816
rect 36044 31804 36050 31816
rect 38194 31804 38200 31816
rect 36044 31776 38200 31804
rect 36044 31764 36050 31776
rect 38194 31764 38200 31776
rect 38252 31764 38258 31816
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1397 31331 1455 31337
rect 1397 31297 1409 31331
rect 1443 31328 1455 31331
rect 1486 31328 1492 31340
rect 1443 31300 1492 31328
rect 1443 31297 1455 31300
rect 1397 31291 1455 31297
rect 1486 31288 1492 31300
rect 1544 31328 1550 31340
rect 2041 31331 2099 31337
rect 2041 31328 2053 31331
rect 1544 31300 2053 31328
rect 1544 31288 1550 31300
rect 2041 31297 2053 31300
rect 2087 31297 2099 31331
rect 37826 31328 37832 31340
rect 37787 31300 37832 31328
rect 2041 31291 2099 31297
rect 37826 31288 37832 31300
rect 37884 31288 37890 31340
rect 1581 31127 1639 31133
rect 1581 31093 1593 31127
rect 1627 31124 1639 31127
rect 2590 31124 2596 31136
rect 1627 31096 2596 31124
rect 1627 31093 1639 31096
rect 1581 31087 1639 31093
rect 2590 31084 2596 31096
rect 2648 31084 2654 31136
rect 38010 31124 38016 31136
rect 37971 31096 38016 31124
rect 38010 31084 38016 31096
rect 38068 31084 38074 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1394 30716 1400 30728
rect 1355 30688 1400 30716
rect 1394 30676 1400 30688
rect 1452 30716 1458 30728
rect 2041 30719 2099 30725
rect 2041 30716 2053 30719
rect 1452 30688 2053 30716
rect 1452 30676 1458 30688
rect 2041 30685 2053 30688
rect 2087 30685 2099 30719
rect 37829 30719 37887 30725
rect 37829 30716 37841 30719
rect 2041 30679 2099 30685
rect 37292 30688 37841 30716
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 2498 30580 2504 30592
rect 1627 30552 2504 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 2498 30540 2504 30552
rect 2556 30540 2562 30592
rect 28442 30540 28448 30592
rect 28500 30580 28506 30592
rect 37292 30589 37320 30688
rect 37829 30685 37841 30688
rect 37875 30685 37887 30719
rect 37829 30679 37887 30685
rect 37277 30583 37335 30589
rect 37277 30580 37289 30583
rect 28500 30552 37289 30580
rect 28500 30540 28506 30552
rect 37277 30549 37289 30552
rect 37323 30549 37335 30583
rect 38010 30580 38016 30592
rect 37971 30552 38016 30580
rect 37277 30543 37335 30549
rect 38010 30540 38016 30552
rect 38068 30540 38074 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 37461 30243 37519 30249
rect 37461 30209 37473 30243
rect 37507 30240 37519 30243
rect 38102 30240 38108 30252
rect 37507 30212 38108 30240
rect 37507 30209 37519 30212
rect 37461 30203 37519 30209
rect 38102 30200 38108 30212
rect 38160 30200 38166 30252
rect 1394 30036 1400 30048
rect 1355 30008 1400 30036
rect 1394 29996 1400 30008
rect 1452 29996 1458 30048
rect 37734 29996 37740 30048
rect 37792 30036 37798 30048
rect 37921 30039 37979 30045
rect 37921 30036 37933 30039
rect 37792 30008 37933 30036
rect 37792 29996 37798 30008
rect 37921 30005 37933 30008
rect 37967 30005 37979 30039
rect 37921 29999 37979 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29628 1458 29640
rect 2041 29631 2099 29637
rect 2041 29628 2053 29631
rect 1452 29600 2053 29628
rect 1452 29588 1458 29600
rect 2041 29597 2053 29600
rect 2087 29597 2099 29631
rect 2041 29591 2099 29597
rect 1578 29492 1584 29504
rect 1539 29464 1584 29492
rect 1578 29452 1584 29464
rect 1636 29452 1642 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1578 29180 1584 29232
rect 1636 29220 1642 29232
rect 1636 29192 2820 29220
rect 1636 29180 1642 29192
rect 2498 29152 2504 29164
rect 2459 29124 2504 29152
rect 2498 29112 2504 29124
rect 2556 29112 2562 29164
rect 2792 29161 2820 29192
rect 2777 29155 2835 29161
rect 2777 29121 2789 29155
rect 2823 29121 2835 29155
rect 2777 29115 2835 29121
rect 37829 29155 37887 29161
rect 37829 29121 37841 29155
rect 37875 29152 37887 29155
rect 38194 29152 38200 29164
rect 37875 29124 38200 29152
rect 37875 29121 37887 29124
rect 37829 29115 37887 29121
rect 38194 29112 38200 29124
rect 38252 29112 38258 29164
rect 2590 29084 2596 29096
rect 2551 29056 2596 29084
rect 2590 29044 2596 29056
rect 2648 29044 2654 29096
rect 1394 29016 1400 29028
rect 1355 28988 1400 29016
rect 1394 28976 1400 28988
rect 1452 28976 1458 29028
rect 2961 29019 3019 29025
rect 2961 28985 2973 29019
rect 3007 29016 3019 29019
rect 3510 29016 3516 29028
rect 3007 28988 3516 29016
rect 3007 28985 3019 28988
rect 2961 28979 3019 28985
rect 3510 28976 3516 28988
rect 3568 28976 3574 29028
rect 38010 29016 38016 29028
rect 37971 28988 38016 29016
rect 38010 28976 38016 28988
rect 38068 28976 38074 29028
rect 1578 28908 1584 28960
rect 1636 28948 1642 28960
rect 2501 28951 2559 28957
rect 2501 28948 2513 28951
rect 1636 28920 2513 28948
rect 1636 28908 1642 28920
rect 2501 28917 2513 28920
rect 2547 28917 2559 28951
rect 2501 28911 2559 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 37829 28543 37887 28549
rect 37829 28540 37841 28543
rect 37292 28512 37841 28540
rect 27614 28364 27620 28416
rect 27672 28404 27678 28416
rect 37292 28413 37320 28512
rect 37829 28509 37841 28512
rect 37875 28509 37887 28543
rect 37829 28503 37887 28509
rect 37277 28407 37335 28413
rect 37277 28404 37289 28407
rect 27672 28376 37289 28404
rect 27672 28364 27678 28376
rect 37277 28373 37289 28376
rect 37323 28373 37335 28407
rect 38010 28404 38016 28416
rect 37971 28376 38016 28404
rect 37277 28367 37335 28373
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 1578 28200 1584 28212
rect 1539 28172 1584 28200
rect 1578 28160 1584 28172
rect 1636 28160 1642 28212
rect 32122 28200 32128 28212
rect 32083 28172 32128 28200
rect 32122 28160 32128 28172
rect 32180 28200 32186 28212
rect 32858 28200 32864 28212
rect 32180 28172 32864 28200
rect 32180 28160 32186 28172
rect 32858 28160 32864 28172
rect 32916 28160 32922 28212
rect 1394 28064 1400 28076
rect 1355 28036 1400 28064
rect 1394 28024 1400 28036
rect 1452 28064 1458 28076
rect 2041 28067 2099 28073
rect 2041 28064 2053 28067
rect 1452 28036 2053 28064
rect 1452 28024 1458 28036
rect 2041 28033 2053 28036
rect 2087 28033 2099 28067
rect 33226 28064 33232 28076
rect 33284 28073 33290 28076
rect 33196 28036 33232 28064
rect 2041 28027 2099 28033
rect 33226 28024 33232 28036
rect 33284 28027 33296 28073
rect 37461 28067 37519 28073
rect 37461 28033 37473 28067
rect 37507 28064 37519 28067
rect 38102 28064 38108 28076
rect 37507 28036 38108 28064
rect 37507 28033 37519 28036
rect 37461 28027 37519 28033
rect 33284 28024 33290 28027
rect 38102 28024 38108 28036
rect 38160 28024 38166 28076
rect 33502 27996 33508 28008
rect 33463 27968 33508 27996
rect 33502 27956 33508 27968
rect 33560 27956 33566 28008
rect 37642 27820 37648 27872
rect 37700 27860 37706 27872
rect 37921 27863 37979 27869
rect 37921 27860 37933 27863
rect 37700 27832 37933 27860
rect 37700 27820 37706 27832
rect 37921 27829 37933 27832
rect 37967 27829 37979 27863
rect 37921 27823 37979 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 25774 27588 25780 27600
rect 25735 27560 25780 27588
rect 25774 27548 25780 27560
rect 25832 27548 25838 27600
rect 33045 27591 33103 27597
rect 33045 27557 33057 27591
rect 33091 27588 33103 27591
rect 33226 27588 33232 27600
rect 33091 27560 33232 27588
rect 33091 27557 33103 27560
rect 33045 27551 33103 27557
rect 33226 27548 33232 27560
rect 33284 27548 33290 27600
rect 36078 27588 36084 27600
rect 36039 27560 36084 27588
rect 36078 27548 36084 27560
rect 36136 27548 36142 27600
rect 32030 27480 32036 27532
rect 32088 27520 32094 27532
rect 32088 27492 32904 27520
rect 32088 27480 32094 27492
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27452 22339 27455
rect 22922 27452 22928 27464
rect 22327 27424 22928 27452
rect 22327 27421 22339 27424
rect 22281 27415 22339 27421
rect 22922 27412 22928 27424
rect 22980 27452 22986 27464
rect 24397 27455 24455 27461
rect 24397 27452 24409 27455
rect 22980 27424 24409 27452
rect 22980 27412 22986 27424
rect 24397 27421 24409 27424
rect 24443 27452 24455 27455
rect 26970 27452 26976 27464
rect 24443 27424 26976 27452
rect 24443 27421 24455 27424
rect 24397 27415 24455 27421
rect 26970 27412 26976 27424
rect 27028 27412 27034 27464
rect 32876 27461 32904 27492
rect 31021 27455 31079 27461
rect 31021 27421 31033 27455
rect 31067 27452 31079 27455
rect 32861 27455 32919 27461
rect 31067 27424 32812 27452
rect 31067 27421 31079 27424
rect 31021 27415 31079 27421
rect 22370 27344 22376 27396
rect 22428 27384 22434 27396
rect 22526 27387 22584 27393
rect 22526 27384 22538 27387
rect 22428 27356 22538 27384
rect 22428 27344 22434 27356
rect 22526 27353 22538 27356
rect 22572 27353 22584 27387
rect 22526 27347 22584 27353
rect 24664 27387 24722 27393
rect 24664 27353 24676 27387
rect 24710 27384 24722 27387
rect 24854 27384 24860 27396
rect 24710 27356 24860 27384
rect 24710 27353 24722 27356
rect 24664 27347 24722 27353
rect 24854 27344 24860 27356
rect 24912 27344 24918 27396
rect 30558 27344 30564 27396
rect 30616 27384 30622 27396
rect 31266 27387 31324 27393
rect 31266 27384 31278 27387
rect 30616 27356 31278 27384
rect 30616 27344 30622 27356
rect 31266 27353 31278 27356
rect 31312 27353 31324 27387
rect 32784 27384 32812 27424
rect 32861 27421 32873 27455
rect 32907 27421 32919 27455
rect 32861 27415 32919 27421
rect 33502 27412 33508 27464
rect 33560 27452 33566 27464
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 33560 27424 34713 27452
rect 33560 27412 33566 27424
rect 34701 27421 34713 27424
rect 34747 27452 34759 27455
rect 35342 27452 35348 27464
rect 34747 27424 35348 27452
rect 34747 27421 34759 27424
rect 34701 27415 34759 27421
rect 35342 27412 35348 27424
rect 35400 27412 35406 27464
rect 37274 27412 37280 27464
rect 37332 27452 37338 27464
rect 37829 27455 37887 27461
rect 37829 27452 37841 27455
rect 37332 27424 37841 27452
rect 37332 27412 37338 27424
rect 37829 27421 37841 27424
rect 37875 27421 37887 27455
rect 37829 27415 37887 27421
rect 33520 27384 33548 27412
rect 32784 27356 33548 27384
rect 31266 27347 31324 27353
rect 34146 27344 34152 27396
rect 34204 27384 34210 27396
rect 34946 27387 35004 27393
rect 34946 27384 34958 27387
rect 34204 27356 34958 27384
rect 34204 27344 34210 27356
rect 34946 27353 34958 27356
rect 34992 27353 35004 27387
rect 36817 27387 36875 27393
rect 36817 27384 36829 27387
rect 34946 27347 35004 27353
rect 35866 27356 36829 27384
rect 23658 27316 23664 27328
rect 23619 27288 23664 27316
rect 23658 27276 23664 27288
rect 23716 27276 23722 27328
rect 32401 27319 32459 27325
rect 32401 27285 32413 27319
rect 32447 27316 32459 27319
rect 32950 27316 32956 27328
rect 32447 27288 32956 27316
rect 32447 27285 32459 27288
rect 32401 27279 32459 27285
rect 32950 27276 32956 27288
rect 33008 27276 33014 27328
rect 33594 27316 33600 27328
rect 33555 27288 33600 27316
rect 33594 27276 33600 27288
rect 33652 27276 33658 27328
rect 33686 27276 33692 27328
rect 33744 27316 33750 27328
rect 35866 27316 35894 27356
rect 36817 27353 36829 27356
rect 36863 27384 36875 27387
rect 37458 27384 37464 27396
rect 36863 27356 37464 27384
rect 36863 27353 36875 27356
rect 36817 27347 36875 27353
rect 37458 27344 37464 27356
rect 37516 27344 37522 27396
rect 33744 27288 35894 27316
rect 33744 27276 33750 27288
rect 37182 27276 37188 27328
rect 37240 27316 37246 27328
rect 37277 27319 37335 27325
rect 37277 27316 37289 27319
rect 37240 27288 37289 27316
rect 37240 27276 37246 27288
rect 37277 27285 37289 27288
rect 37323 27285 37335 27319
rect 38010 27316 38016 27328
rect 37971 27288 38016 27316
rect 37277 27279 37335 27285
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 22465 27115 22523 27121
rect 22465 27081 22477 27115
rect 22511 27081 22523 27115
rect 24854 27112 24860 27124
rect 24815 27084 24860 27112
rect 22465 27075 22523 27081
rect 22480 27044 22508 27075
rect 24854 27072 24860 27084
rect 24912 27072 24918 27124
rect 28350 27112 28356 27124
rect 28311 27084 28356 27112
rect 28350 27072 28356 27084
rect 28408 27072 28414 27124
rect 30558 27112 30564 27124
rect 30519 27084 30564 27112
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 31294 27112 31300 27124
rect 31036 27084 31300 27112
rect 23170 27047 23228 27053
rect 23170 27044 23182 27047
rect 22480 27016 23182 27044
rect 23170 27013 23182 27016
rect 23216 27013 23228 27047
rect 27522 27044 27528 27056
rect 23170 27007 23228 27013
rect 26988 27016 27528 27044
rect 26988 26988 27016 27016
rect 27522 27004 27528 27016
rect 27580 27004 27586 27056
rect 31036 27053 31064 27084
rect 31294 27072 31300 27084
rect 31352 27112 31358 27124
rect 33594 27112 33600 27124
rect 31352 27084 33600 27112
rect 31352 27072 31358 27084
rect 33594 27072 33600 27084
rect 33652 27072 33658 27124
rect 34146 27112 34152 27124
rect 34107 27084 34152 27112
rect 34146 27072 34152 27084
rect 34204 27072 34210 27124
rect 36630 27072 36636 27124
rect 36688 27112 36694 27124
rect 37921 27115 37979 27121
rect 37921 27112 37933 27115
rect 36688 27084 37933 27112
rect 36688 27072 36694 27084
rect 37921 27081 37933 27084
rect 37967 27081 37979 27115
rect 37921 27075 37979 27081
rect 29917 27047 29975 27053
rect 29917 27013 29929 27047
rect 29963 27044 29975 27047
rect 31021 27047 31079 27053
rect 31021 27044 31033 27047
rect 29963 27016 31033 27044
rect 29963 27013 29975 27016
rect 29917 27007 29975 27013
rect 31021 27013 31033 27016
rect 31067 27013 31079 27047
rect 33502 27044 33508 27056
rect 31021 27007 31079 27013
rect 32140 27016 33508 27044
rect 1394 26976 1400 26988
rect 1355 26948 1400 26976
rect 1394 26936 1400 26948
rect 1452 26976 1458 26988
rect 2041 26979 2099 26985
rect 2041 26976 2053 26979
rect 1452 26948 2053 26976
rect 1452 26936 1458 26948
rect 2041 26945 2053 26948
rect 2087 26945 2099 26979
rect 22278 26976 22284 26988
rect 22239 26948 22284 26976
rect 2041 26939 2099 26945
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 22922 26976 22928 26988
rect 22883 26948 22928 26976
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 23474 26936 23480 26988
rect 23532 26976 23538 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 23532 26948 25053 26976
rect 23532 26936 23538 26948
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 26970 26976 26976 26988
rect 26931 26948 26976 26976
rect 25041 26939 25099 26945
rect 26970 26936 26976 26948
rect 27028 26936 27034 26988
rect 27062 26936 27068 26988
rect 27120 26976 27126 26988
rect 27229 26979 27287 26985
rect 27229 26976 27241 26979
rect 27120 26948 27241 26976
rect 27120 26936 27126 26948
rect 27229 26945 27241 26948
rect 27275 26945 27287 26979
rect 27229 26939 27287 26945
rect 30377 26979 30435 26985
rect 30377 26945 30389 26979
rect 30423 26976 30435 26979
rect 30834 26976 30840 26988
rect 30423 26948 30840 26976
rect 30423 26945 30435 26948
rect 30377 26939 30435 26945
rect 30834 26936 30840 26948
rect 30892 26936 30898 26988
rect 32140 26985 32168 27016
rect 33502 27004 33508 27016
rect 33560 27004 33566 27056
rect 35986 27004 35992 27056
rect 36044 27044 36050 27056
rect 38378 27044 38384 27056
rect 36044 27016 38384 27044
rect 36044 27004 36050 27016
rect 38378 27004 38384 27016
rect 38436 27004 38442 27056
rect 32125 26979 32183 26985
rect 32125 26945 32137 26979
rect 32171 26945 32183 26979
rect 32125 26939 32183 26945
rect 32214 26936 32220 26988
rect 32272 26976 32278 26988
rect 32381 26979 32439 26985
rect 32381 26976 32393 26979
rect 32272 26948 32393 26976
rect 32272 26936 32278 26948
rect 32381 26945 32393 26948
rect 32427 26945 32439 26979
rect 32381 26939 32439 26945
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26976 34023 26979
rect 34146 26976 34152 26988
rect 34011 26948 34152 26976
rect 34011 26945 34023 26948
rect 33965 26939 34023 26945
rect 34146 26936 34152 26948
rect 34204 26936 34210 26988
rect 37182 26936 37188 26988
rect 37240 26976 37246 26988
rect 38105 26979 38163 26985
rect 38105 26976 38117 26979
rect 37240 26948 38117 26976
rect 37240 26936 37246 26948
rect 38105 26945 38117 26948
rect 38151 26945 38163 26979
rect 38105 26939 38163 26945
rect 31128 26880 31892 26908
rect 31128 26840 31156 26880
rect 31386 26840 31392 26852
rect 28276 26812 31156 26840
rect 31347 26812 31392 26840
rect 1581 26775 1639 26781
rect 1581 26741 1593 26775
rect 1627 26772 1639 26775
rect 2866 26772 2872 26784
rect 1627 26744 2872 26772
rect 1627 26741 1639 26744
rect 1581 26735 1639 26741
rect 2866 26732 2872 26744
rect 2924 26732 2930 26784
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 24305 26775 24363 26781
rect 24305 26772 24317 26775
rect 23624 26744 24317 26772
rect 23624 26732 23630 26744
rect 24305 26741 24317 26744
rect 24351 26772 24363 26775
rect 28276 26772 28304 26812
rect 31386 26800 31392 26812
rect 31444 26800 31450 26852
rect 24351 26744 28304 26772
rect 31481 26775 31539 26781
rect 24351 26741 24363 26744
rect 24305 26735 24363 26741
rect 31481 26741 31493 26775
rect 31527 26772 31539 26775
rect 31754 26772 31760 26784
rect 31527 26744 31760 26772
rect 31527 26741 31539 26744
rect 31481 26735 31539 26741
rect 31754 26732 31760 26744
rect 31812 26732 31818 26784
rect 31864 26772 31892 26880
rect 33502 26868 33508 26920
rect 33560 26908 33566 26920
rect 36998 26908 37004 26920
rect 33560 26880 37004 26908
rect 33560 26868 33566 26880
rect 36998 26868 37004 26880
rect 37056 26868 37062 26920
rect 37366 26868 37372 26920
rect 37424 26868 37430 26920
rect 37384 26840 37412 26868
rect 33060 26812 37412 26840
rect 33060 26772 33088 26812
rect 33502 26772 33508 26784
rect 31864 26744 33088 26772
rect 33463 26744 33508 26772
rect 33502 26732 33508 26744
rect 33560 26732 33566 26784
rect 36633 26775 36691 26781
rect 36633 26741 36645 26775
rect 36679 26772 36691 26775
rect 37090 26772 37096 26784
rect 36679 26744 37096 26772
rect 36679 26741 36691 26744
rect 36633 26735 36691 26741
rect 37090 26732 37096 26744
rect 37148 26732 37154 26784
rect 37366 26732 37372 26784
rect 37424 26772 37430 26784
rect 37461 26775 37519 26781
rect 37461 26772 37473 26775
rect 37424 26744 37473 26772
rect 37424 26732 37430 26744
rect 37461 26741 37473 26744
rect 37507 26772 37519 26775
rect 38378 26772 38384 26784
rect 37507 26744 38384 26772
rect 37507 26741 37519 26744
rect 37461 26735 37519 26741
rect 38378 26732 38384 26744
rect 38436 26732 38442 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 22370 26568 22376 26580
rect 22331 26540 22376 26568
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 23474 26568 23480 26580
rect 23435 26540 23480 26568
rect 23474 26528 23480 26540
rect 23532 26528 23538 26580
rect 26421 26571 26479 26577
rect 26421 26537 26433 26571
rect 26467 26568 26479 26571
rect 27062 26568 27068 26580
rect 26467 26540 27068 26568
rect 26467 26537 26479 26540
rect 26421 26531 26479 26537
rect 27062 26528 27068 26540
rect 27120 26528 27126 26580
rect 30834 26568 30840 26580
rect 27356 26540 30420 26568
rect 30795 26540 30840 26568
rect 23382 26500 23388 26512
rect 23343 26472 23388 26500
rect 23382 26460 23388 26472
rect 23440 26460 23446 26512
rect 24670 26460 24676 26512
rect 24728 26500 24734 26512
rect 25041 26503 25099 26509
rect 25041 26500 25053 26503
rect 24728 26472 25053 26500
rect 24728 26460 24734 26472
rect 25041 26469 25053 26472
rect 25087 26500 25099 26503
rect 27356 26500 27384 26540
rect 30282 26500 30288 26512
rect 25087 26472 27384 26500
rect 30243 26472 30288 26500
rect 25087 26469 25099 26472
rect 25041 26463 25099 26469
rect 30282 26460 30288 26472
rect 30340 26460 30346 26512
rect 30392 26500 30420 26540
rect 30834 26528 30840 26540
rect 30892 26528 30898 26580
rect 31941 26571 31999 26577
rect 31941 26537 31953 26571
rect 31987 26568 31999 26571
rect 32214 26568 32220 26580
rect 31987 26540 32220 26568
rect 31987 26537 31999 26540
rect 31941 26531 31999 26537
rect 32214 26528 32220 26540
rect 32272 26528 32278 26580
rect 34057 26571 34115 26577
rect 32324 26540 34008 26568
rect 30926 26500 30932 26512
rect 30392 26472 30788 26500
rect 30887 26472 30932 26500
rect 30377 26435 30435 26441
rect 30377 26401 30389 26435
rect 30423 26401 30435 26435
rect 30760 26432 30788 26472
rect 30926 26460 30932 26472
rect 30984 26460 30990 26512
rect 32324 26432 32352 26540
rect 33137 26503 33195 26509
rect 33137 26469 33149 26503
rect 33183 26500 33195 26503
rect 33873 26503 33931 26509
rect 33873 26500 33885 26503
rect 33183 26472 33885 26500
rect 33183 26469 33195 26472
rect 33137 26463 33195 26469
rect 33873 26469 33885 26472
rect 33919 26469 33931 26503
rect 33980 26500 34008 26540
rect 34057 26537 34069 26571
rect 34103 26568 34115 26571
rect 34146 26568 34152 26580
rect 34103 26540 34152 26568
rect 34103 26537 34115 26540
rect 34057 26531 34115 26537
rect 34146 26528 34152 26540
rect 34204 26528 34210 26580
rect 35986 26568 35992 26580
rect 35866 26540 35992 26568
rect 35866 26500 35894 26540
rect 35986 26528 35992 26540
rect 36044 26528 36050 26580
rect 36262 26568 36268 26580
rect 36175 26540 36268 26568
rect 36262 26528 36268 26540
rect 36320 26568 36326 26580
rect 37366 26568 37372 26580
rect 36320 26540 37372 26568
rect 36320 26528 36326 26540
rect 37366 26528 37372 26540
rect 37424 26528 37430 26580
rect 33980 26472 35894 26500
rect 33873 26463 33931 26469
rect 37090 26460 37096 26512
rect 37148 26500 37154 26512
rect 38010 26500 38016 26512
rect 37148 26472 37412 26500
rect 37971 26472 38016 26500
rect 37148 26460 37154 26472
rect 32582 26432 32588 26444
rect 30760 26404 32352 26432
rect 32543 26404 32588 26432
rect 30377 26395 30435 26401
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 22557 26367 22615 26373
rect 1719 26336 2268 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 2240 26308 2268 26336
rect 22557 26333 22569 26367
rect 22603 26364 22615 26367
rect 22646 26364 22652 26376
rect 22603 26336 22652 26364
rect 22603 26333 22615 26336
rect 22557 26327 22615 26333
rect 22646 26324 22652 26336
rect 22704 26324 22710 26376
rect 26234 26324 26240 26376
rect 26292 26364 26298 26376
rect 26292 26336 26337 26364
rect 26292 26324 26298 26336
rect 27522 26324 27528 26376
rect 27580 26364 27586 26376
rect 28261 26367 28319 26373
rect 28261 26364 28273 26367
rect 27580 26336 28273 26364
rect 27580 26324 27586 26336
rect 28261 26333 28273 26336
rect 28307 26333 28319 26367
rect 30392 26364 30420 26395
rect 32582 26392 32588 26404
rect 32640 26392 32646 26444
rect 32677 26435 32735 26441
rect 32677 26401 32689 26435
rect 32723 26432 32735 26435
rect 36078 26432 36084 26444
rect 32723 26404 36084 26432
rect 32723 26401 32735 26404
rect 32677 26395 32735 26401
rect 36078 26392 36084 26404
rect 36136 26392 36142 26444
rect 36538 26392 36544 26444
rect 36596 26432 36602 26444
rect 36596 26404 37136 26432
rect 36596 26392 36602 26404
rect 31754 26364 31760 26376
rect 30392 26336 31432 26364
rect 31715 26336 31760 26364
rect 28261 26327 28319 26333
rect 2222 26296 2228 26308
rect 2183 26268 2228 26296
rect 2222 26256 2228 26268
rect 2280 26256 2286 26308
rect 21913 26299 21971 26305
rect 21913 26265 21925 26299
rect 21959 26296 21971 26299
rect 22922 26296 22928 26308
rect 21959 26268 22928 26296
rect 21959 26265 21971 26268
rect 21913 26259 21971 26265
rect 22922 26256 22928 26268
rect 22980 26296 22986 26308
rect 23017 26299 23075 26305
rect 23017 26296 23029 26299
rect 22980 26268 23029 26296
rect 22980 26256 22986 26268
rect 23017 26265 23029 26268
rect 23063 26296 23075 26299
rect 24397 26299 24455 26305
rect 24397 26296 24409 26299
rect 23063 26268 24409 26296
rect 23063 26265 23075 26268
rect 23017 26259 23075 26265
rect 24397 26265 24409 26268
rect 24443 26265 24455 26299
rect 27614 26296 27620 26308
rect 24397 26259 24455 26265
rect 26896 26268 27620 26296
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 23750 26188 23756 26240
rect 23808 26228 23814 26240
rect 24670 26228 24676 26240
rect 23808 26200 24676 26228
rect 23808 26188 23814 26200
rect 24670 26188 24676 26200
rect 24728 26188 24734 26240
rect 26896 26237 26924 26268
rect 27614 26256 27620 26268
rect 27672 26256 27678 26308
rect 27890 26256 27896 26308
rect 27948 26296 27954 26308
rect 27994 26299 28052 26305
rect 27994 26296 28006 26299
rect 27948 26268 28006 26296
rect 27948 26256 27954 26268
rect 27994 26265 28006 26268
rect 28040 26265 28052 26299
rect 27994 26259 28052 26265
rect 29917 26299 29975 26305
rect 29917 26265 29929 26299
rect 29963 26296 29975 26299
rect 31294 26296 31300 26308
rect 29963 26268 31300 26296
rect 29963 26265 29975 26268
rect 29917 26259 29975 26265
rect 31294 26256 31300 26268
rect 31352 26256 31358 26308
rect 31404 26296 31432 26336
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 33594 26364 33600 26376
rect 33555 26336 33600 26364
rect 33594 26324 33600 26336
rect 33652 26324 33658 26376
rect 36262 26324 36268 26376
rect 36320 26364 36326 26376
rect 36863 26367 36921 26373
rect 36863 26364 36875 26367
rect 36320 26336 36875 26364
rect 36320 26324 36326 26336
rect 36863 26333 36875 26336
rect 36909 26333 36921 26367
rect 36998 26364 37004 26376
rect 36959 26336 37004 26364
rect 36863 26327 36921 26333
rect 36998 26324 37004 26336
rect 37056 26324 37062 26376
rect 37108 26373 37136 26404
rect 37384 26373 37412 26472
rect 38010 26460 38016 26472
rect 38068 26460 38074 26512
rect 37093 26367 37151 26373
rect 37093 26333 37105 26367
rect 37139 26333 37151 26367
rect 37093 26327 37151 26333
rect 37276 26367 37334 26373
rect 37276 26333 37288 26367
rect 37322 26333 37334 26367
rect 37276 26327 37334 26333
rect 37369 26367 37427 26373
rect 37369 26333 37381 26367
rect 37415 26333 37427 26367
rect 37369 26327 37427 26333
rect 32030 26296 32036 26308
rect 31404 26268 32036 26296
rect 32030 26256 32036 26268
rect 32088 26256 32094 26308
rect 32769 26299 32827 26305
rect 32769 26265 32781 26299
rect 32815 26296 32827 26299
rect 33134 26296 33140 26308
rect 32815 26268 33140 26296
rect 32815 26265 32827 26268
rect 32769 26259 32827 26265
rect 33134 26256 33140 26268
rect 33192 26256 33198 26308
rect 34701 26299 34759 26305
rect 34701 26296 34713 26299
rect 33704 26268 34713 26296
rect 26881 26231 26939 26237
rect 26881 26197 26893 26231
rect 26927 26228 26939 26231
rect 26927 26200 26961 26228
rect 26927 26197 26939 26200
rect 26881 26191 26939 26197
rect 32582 26188 32588 26240
rect 32640 26228 32646 26240
rect 33704 26228 33732 26268
rect 34701 26265 34713 26268
rect 34747 26265 34759 26299
rect 37292 26296 37320 26327
rect 37458 26324 37464 26376
rect 37516 26364 37522 26376
rect 37829 26367 37887 26373
rect 37829 26364 37841 26367
rect 37516 26336 37841 26364
rect 37516 26324 37522 26336
rect 37829 26333 37841 26336
rect 37875 26333 37887 26367
rect 37829 26327 37887 26333
rect 38286 26324 38292 26376
rect 38344 26324 38350 26376
rect 38304 26296 38332 26324
rect 37292 26268 38332 26296
rect 34701 26259 34759 26265
rect 36722 26228 36728 26240
rect 32640 26200 33732 26228
rect 36683 26200 36728 26228
rect 32640 26188 32646 26200
rect 36722 26188 36728 26200
rect 36780 26188 36786 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 22189 26027 22247 26033
rect 22189 25993 22201 26027
rect 22235 26024 22247 26027
rect 22278 26024 22284 26036
rect 22235 25996 22284 26024
rect 22235 25993 22247 25996
rect 22189 25987 22247 25993
rect 22278 25984 22284 25996
rect 22336 25984 22342 26036
rect 26234 25984 26240 26036
rect 26292 26024 26298 26036
rect 26973 26027 27031 26033
rect 26973 26024 26985 26027
rect 26292 25996 26985 26024
rect 26292 25984 26298 25996
rect 26973 25993 26985 25996
rect 27019 25993 27031 26027
rect 27890 26024 27896 26036
rect 27851 25996 27896 26024
rect 26973 25987 27031 25993
rect 27890 25984 27896 25996
rect 27948 25984 27954 26036
rect 30837 26027 30895 26033
rect 30837 25993 30849 26027
rect 30883 26024 30895 26027
rect 30926 26024 30932 26036
rect 30883 25996 30932 26024
rect 30883 25993 30895 25996
rect 30837 25987 30895 25993
rect 30926 25984 30932 25996
rect 30984 25984 30990 26036
rect 31386 25984 31392 26036
rect 31444 26024 31450 26036
rect 32125 26027 32183 26033
rect 32125 26024 32137 26027
rect 31444 25996 32137 26024
rect 31444 25984 31450 25996
rect 32125 25993 32137 25996
rect 32171 25993 32183 26027
rect 32125 25987 32183 25993
rect 32585 26027 32643 26033
rect 32585 25993 32597 26027
rect 32631 26024 32643 26027
rect 33502 26024 33508 26036
rect 32631 25996 33508 26024
rect 32631 25993 32643 25996
rect 32585 25987 32643 25993
rect 33502 25984 33508 25996
rect 33560 25984 33566 26036
rect 37550 26024 37556 26036
rect 35866 25996 37556 26024
rect 31297 25959 31355 25965
rect 31297 25925 31309 25959
rect 31343 25956 31355 25959
rect 32950 25956 32956 25968
rect 31343 25928 32956 25956
rect 31343 25925 31355 25928
rect 31297 25919 31355 25925
rect 32950 25916 32956 25928
rect 33008 25956 33014 25968
rect 35866 25956 35894 25996
rect 37550 25984 37556 25996
rect 37608 26024 37614 26036
rect 37608 25996 37688 26024
rect 37608 25984 37614 25996
rect 36906 25956 36912 25968
rect 33008 25928 35894 25956
rect 36648 25928 36912 25956
rect 33008 25916 33014 25928
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25888 1458 25900
rect 2317 25891 2375 25897
rect 2317 25888 2329 25891
rect 1452 25860 2329 25888
rect 1452 25848 1458 25860
rect 2317 25857 2329 25860
rect 2363 25857 2375 25891
rect 21174 25888 21180 25900
rect 2317 25851 2375 25857
rect 6886 25860 21180 25888
rect 1673 25823 1731 25829
rect 1673 25789 1685 25823
rect 1719 25820 1731 25823
rect 6886 25820 6914 25860
rect 21174 25848 21180 25860
rect 21232 25888 21238 25900
rect 23477 25891 23535 25897
rect 23477 25888 23489 25891
rect 21232 25860 23489 25888
rect 21232 25848 21238 25860
rect 23477 25857 23489 25860
rect 23523 25888 23535 25891
rect 28074 25888 28080 25900
rect 23523 25860 27936 25888
rect 28035 25860 28080 25888
rect 23523 25857 23535 25860
rect 23477 25851 23535 25857
rect 1719 25792 6914 25820
rect 1719 25789 1731 25792
rect 1673 25783 1731 25789
rect 22462 25780 22468 25832
rect 22520 25820 22526 25832
rect 22649 25823 22707 25829
rect 22649 25820 22661 25823
rect 22520 25792 22661 25820
rect 22520 25780 22526 25792
rect 22649 25789 22661 25792
rect 22695 25820 22707 25823
rect 22922 25820 22928 25832
rect 22695 25792 22928 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 22922 25780 22928 25792
rect 22980 25780 22986 25832
rect 23569 25823 23627 25829
rect 23569 25789 23581 25823
rect 23615 25820 23627 25823
rect 23658 25820 23664 25832
rect 23615 25792 23664 25820
rect 23615 25789 23627 25792
rect 23569 25783 23627 25789
rect 23658 25780 23664 25792
rect 23716 25780 23722 25832
rect 23753 25823 23811 25829
rect 23753 25789 23765 25823
rect 23799 25820 23811 25823
rect 25225 25823 25283 25829
rect 25225 25820 25237 25823
rect 23799 25792 25237 25820
rect 23799 25789 23811 25792
rect 23753 25783 23811 25789
rect 25225 25789 25237 25792
rect 25271 25820 25283 25823
rect 25777 25823 25835 25829
rect 25777 25820 25789 25823
rect 25271 25792 25789 25820
rect 25271 25789 25283 25792
rect 25225 25783 25283 25789
rect 25777 25789 25789 25792
rect 25823 25820 25835 25823
rect 26234 25820 26240 25832
rect 25823 25792 26240 25820
rect 25823 25789 25835 25792
rect 25777 25783 25835 25789
rect 26234 25780 26240 25792
rect 26292 25780 26298 25832
rect 27430 25820 27436 25832
rect 27391 25792 27436 25820
rect 27430 25780 27436 25792
rect 27488 25780 27494 25832
rect 22373 25755 22431 25761
rect 22373 25721 22385 25755
rect 22419 25752 22431 25755
rect 23014 25752 23020 25764
rect 22419 25724 23020 25752
rect 22419 25721 22431 25724
rect 22373 25715 22431 25721
rect 23014 25712 23020 25724
rect 23072 25712 23078 25764
rect 27062 25752 27068 25764
rect 27023 25724 27068 25752
rect 27062 25712 27068 25724
rect 27120 25712 27126 25764
rect 27908 25752 27936 25860
rect 28074 25848 28080 25860
rect 28132 25848 28138 25900
rect 30374 25888 30380 25900
rect 30287 25860 30380 25888
rect 30374 25848 30380 25860
rect 30432 25888 30438 25900
rect 31205 25891 31263 25897
rect 31205 25888 31217 25891
rect 30432 25860 31217 25888
rect 30432 25848 30438 25860
rect 31205 25857 31217 25860
rect 31251 25857 31263 25891
rect 31205 25851 31263 25857
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25888 32551 25891
rect 32766 25888 32772 25900
rect 32539 25860 32772 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 32766 25848 32772 25860
rect 32824 25848 32830 25900
rect 36262 25897 36268 25900
rect 35621 25891 35679 25897
rect 35621 25857 35633 25891
rect 35667 25888 35679 25891
rect 36260 25888 36268 25897
rect 35667 25860 36268 25888
rect 35667 25857 35679 25860
rect 35621 25851 35679 25857
rect 36260 25851 36268 25860
rect 36262 25848 36268 25851
rect 36320 25848 36326 25900
rect 36357 25891 36415 25897
rect 36357 25857 36369 25891
rect 36403 25857 36415 25891
rect 36357 25851 36415 25857
rect 36449 25891 36507 25897
rect 36449 25857 36461 25891
rect 36495 25888 36507 25891
rect 36538 25888 36544 25900
rect 36495 25860 36544 25888
rect 36495 25857 36507 25860
rect 36449 25851 36507 25857
rect 31481 25823 31539 25829
rect 31481 25789 31493 25823
rect 31527 25820 31539 25823
rect 32582 25820 32588 25832
rect 31527 25792 32588 25820
rect 31527 25789 31539 25792
rect 31481 25783 31539 25789
rect 32582 25780 32588 25792
rect 32640 25820 32646 25832
rect 32677 25823 32735 25829
rect 32677 25820 32689 25823
rect 32640 25792 32689 25820
rect 32640 25780 32646 25792
rect 32677 25789 32689 25792
rect 32723 25789 32735 25823
rect 32677 25783 32735 25789
rect 32858 25780 32864 25832
rect 32916 25820 32922 25832
rect 36372 25820 36400 25851
rect 36538 25848 36544 25860
rect 36596 25848 36602 25900
rect 36648 25897 36676 25928
rect 36906 25916 36912 25928
rect 36964 25916 36970 25968
rect 37660 25965 37688 25996
rect 37645 25959 37703 25965
rect 37645 25925 37657 25959
rect 37691 25925 37703 25959
rect 37645 25919 37703 25925
rect 37826 25916 37832 25968
rect 37884 25956 37890 25968
rect 38194 25956 38200 25968
rect 37884 25928 38200 25956
rect 37884 25916 37890 25928
rect 38194 25916 38200 25928
rect 38252 25916 38258 25968
rect 36632 25891 36690 25897
rect 36632 25857 36644 25891
rect 36678 25857 36690 25891
rect 36632 25851 36690 25857
rect 36725 25891 36783 25897
rect 36725 25857 36737 25891
rect 36771 25888 36783 25891
rect 37090 25888 37096 25900
rect 36771 25860 37096 25888
rect 36771 25857 36783 25860
rect 36725 25851 36783 25857
rect 32916 25792 36400 25820
rect 32916 25780 32922 25792
rect 33134 25752 33140 25764
rect 27908 25724 33140 25752
rect 33134 25712 33140 25724
rect 33192 25752 33198 25764
rect 33873 25755 33931 25761
rect 33873 25752 33885 25755
rect 33192 25724 33885 25752
rect 33192 25712 33198 25724
rect 33873 25721 33885 25724
rect 33919 25721 33931 25755
rect 33873 25715 33931 25721
rect 35069 25755 35127 25761
rect 35069 25721 35081 25755
rect 35115 25752 35127 25755
rect 36262 25752 36268 25764
rect 35115 25724 36268 25752
rect 35115 25721 35127 25724
rect 35069 25715 35127 25721
rect 36262 25712 36268 25724
rect 36320 25752 36326 25764
rect 36740 25752 36768 25851
rect 37090 25848 37096 25860
rect 37148 25848 37154 25900
rect 37550 25897 37556 25900
rect 37548 25888 37556 25897
rect 37511 25860 37556 25888
rect 37548 25851 37556 25860
rect 37550 25848 37556 25851
rect 37608 25848 37614 25900
rect 37737 25891 37795 25897
rect 37737 25857 37749 25891
rect 37783 25857 37795 25891
rect 37918 25888 37924 25900
rect 37879 25860 37924 25888
rect 37737 25851 37795 25857
rect 36998 25780 37004 25832
rect 37056 25820 37062 25832
rect 37752 25820 37780 25851
rect 37918 25848 37924 25860
rect 37976 25848 37982 25900
rect 38013 25891 38071 25897
rect 38013 25857 38025 25891
rect 38059 25888 38071 25891
rect 38059 25860 38424 25888
rect 38059 25857 38071 25860
rect 38013 25851 38071 25857
rect 37056 25792 37780 25820
rect 37056 25780 37062 25792
rect 36320 25724 37504 25752
rect 36320 25712 36326 25724
rect 21174 25684 21180 25696
rect 21135 25656 21180 25684
rect 21174 25644 21180 25656
rect 21232 25644 21238 25696
rect 22554 25644 22560 25696
rect 22612 25684 22618 25696
rect 23109 25687 23167 25693
rect 23109 25684 23121 25687
rect 22612 25656 23121 25684
rect 22612 25644 22618 25656
rect 23109 25653 23121 25656
rect 23155 25653 23167 25687
rect 24394 25684 24400 25696
rect 24355 25656 24400 25684
rect 23109 25647 23167 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 32582 25644 32588 25696
rect 32640 25684 32646 25696
rect 33321 25687 33379 25693
rect 33321 25684 33333 25687
rect 32640 25656 33333 25684
rect 32640 25644 32646 25656
rect 33321 25653 33333 25656
rect 33367 25653 33379 25687
rect 36078 25684 36084 25696
rect 36039 25656 36084 25684
rect 33321 25647 33379 25653
rect 36078 25644 36084 25656
rect 36136 25644 36142 25696
rect 37366 25684 37372 25696
rect 37327 25656 37372 25684
rect 37366 25644 37372 25656
rect 37424 25644 37430 25696
rect 37476 25684 37504 25724
rect 37550 25712 37556 25764
rect 37608 25752 37614 25764
rect 37826 25752 37832 25764
rect 37608 25724 37832 25752
rect 37608 25712 37614 25724
rect 37826 25712 37832 25724
rect 37884 25752 37890 25764
rect 38286 25752 38292 25764
rect 37884 25724 38292 25752
rect 37884 25712 37890 25724
rect 38286 25712 38292 25724
rect 38344 25712 38350 25764
rect 38396 25684 38424 25860
rect 37476 25656 38424 25684
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 22646 25480 22652 25492
rect 22607 25452 22652 25480
rect 22646 25440 22652 25452
rect 22704 25440 22710 25492
rect 23014 25440 23020 25492
rect 23072 25480 23078 25492
rect 23109 25483 23167 25489
rect 23109 25480 23121 25483
rect 23072 25452 23121 25480
rect 23072 25440 23078 25452
rect 23109 25449 23121 25452
rect 23155 25449 23167 25483
rect 23109 25443 23167 25449
rect 23382 25440 23388 25492
rect 23440 25480 23446 25492
rect 24397 25483 24455 25489
rect 24397 25480 24409 25483
rect 23440 25452 24409 25480
rect 23440 25440 23446 25452
rect 24397 25449 24409 25452
rect 24443 25449 24455 25483
rect 24397 25443 24455 25449
rect 25685 25483 25743 25489
rect 25685 25449 25697 25483
rect 25731 25480 25743 25483
rect 25774 25480 25780 25492
rect 25731 25452 25780 25480
rect 25731 25449 25743 25452
rect 25685 25443 25743 25449
rect 25774 25440 25780 25452
rect 25832 25440 25838 25492
rect 28442 25480 28448 25492
rect 28403 25452 28448 25480
rect 28442 25440 28448 25452
rect 28500 25440 28506 25492
rect 30282 25440 30288 25492
rect 30340 25480 30346 25492
rect 31573 25483 31631 25489
rect 31573 25480 31585 25483
rect 30340 25452 31585 25480
rect 30340 25440 30346 25452
rect 31573 25449 31585 25452
rect 31619 25449 31631 25483
rect 31573 25443 31631 25449
rect 36170 25440 36176 25492
rect 36228 25480 36234 25492
rect 36228 25452 37780 25480
rect 36228 25440 36234 25452
rect 1581 25415 1639 25421
rect 1581 25381 1593 25415
rect 1627 25412 1639 25415
rect 2774 25412 2780 25424
rect 1627 25384 2780 25412
rect 1627 25381 1639 25384
rect 1581 25375 1639 25381
rect 2774 25372 2780 25384
rect 2832 25372 2838 25424
rect 22554 25412 22560 25424
rect 22515 25384 22560 25412
rect 22554 25372 22560 25384
rect 22612 25372 22618 25424
rect 36909 25415 36967 25421
rect 36909 25381 36921 25415
rect 36955 25412 36967 25415
rect 37274 25412 37280 25424
rect 36955 25384 37280 25412
rect 36955 25381 36967 25384
rect 36909 25375 36967 25381
rect 23566 25344 23572 25356
rect 23527 25316 23572 25344
rect 23566 25304 23572 25316
rect 23624 25304 23630 25356
rect 23753 25347 23811 25353
rect 23753 25313 23765 25347
rect 23799 25344 23811 25347
rect 25041 25347 25099 25353
rect 25041 25344 25053 25347
rect 23799 25316 25053 25344
rect 23799 25313 23811 25316
rect 23753 25307 23811 25313
rect 25041 25313 25053 25316
rect 25087 25344 25099 25347
rect 26234 25344 26240 25356
rect 25087 25316 26240 25344
rect 25087 25313 25099 25316
rect 25041 25307 25099 25313
rect 26234 25304 26240 25316
rect 26292 25304 26298 25356
rect 32217 25347 32275 25353
rect 32217 25313 32229 25347
rect 32263 25344 32275 25347
rect 32582 25344 32588 25356
rect 32263 25316 32588 25344
rect 32263 25313 32275 25316
rect 32217 25307 32275 25313
rect 32582 25304 32588 25316
rect 32640 25344 32646 25356
rect 33321 25347 33379 25353
rect 33321 25344 33333 25347
rect 32640 25316 33333 25344
rect 32640 25304 32646 25316
rect 33321 25313 33333 25316
rect 33367 25313 33379 25347
rect 33321 25307 33379 25313
rect 35342 25304 35348 25356
rect 35400 25344 35406 25356
rect 35529 25347 35587 25353
rect 35529 25344 35541 25347
rect 35400 25316 35541 25344
rect 35400 25304 35406 25316
rect 35529 25313 35541 25316
rect 35575 25313 35587 25347
rect 35529 25307 35587 25313
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25276 1458 25288
rect 2041 25279 2099 25285
rect 2041 25276 2053 25279
rect 1452 25248 2053 25276
rect 1452 25236 1458 25248
rect 2041 25245 2053 25248
rect 2087 25245 2099 25279
rect 2041 25239 2099 25245
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 24857 25279 24915 25285
rect 24857 25276 24869 25279
rect 24544 25248 24869 25276
rect 24544 25236 24550 25248
rect 24857 25245 24869 25248
rect 24903 25276 24915 25279
rect 25774 25276 25780 25288
rect 24903 25248 25780 25276
rect 24903 25245 24915 25248
rect 24857 25239 24915 25245
rect 25774 25236 25780 25248
rect 25832 25236 25838 25288
rect 27065 25279 27123 25285
rect 26252 25248 27016 25276
rect 22189 25211 22247 25217
rect 22189 25177 22201 25211
rect 22235 25208 22247 25211
rect 22462 25208 22468 25220
rect 22235 25180 22468 25208
rect 22235 25177 22247 25180
rect 22189 25171 22247 25177
rect 22462 25168 22468 25180
rect 22520 25168 22526 25220
rect 24670 25208 24676 25220
rect 23492 25180 24676 25208
rect 2682 25140 2688 25152
rect 2643 25112 2688 25140
rect 2682 25100 2688 25112
rect 2740 25100 2746 25152
rect 21634 25140 21640 25152
rect 21595 25112 21640 25140
rect 21634 25100 21640 25112
rect 21692 25140 21698 25152
rect 23492 25149 23520 25180
rect 24670 25168 24676 25180
rect 24728 25208 24734 25220
rect 26252 25208 26280 25248
rect 24728 25180 26280 25208
rect 24728 25168 24734 25180
rect 23477 25143 23535 25149
rect 23477 25140 23489 25143
rect 21692 25112 23489 25140
rect 21692 25100 21698 25112
rect 23477 25109 23489 25112
rect 23523 25109 23535 25143
rect 23477 25103 23535 25109
rect 24394 25100 24400 25152
rect 24452 25140 24458 25152
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 24452 25112 24777 25140
rect 24452 25100 24458 25112
rect 24765 25109 24777 25112
rect 24811 25140 24823 25143
rect 25866 25140 25872 25152
rect 24811 25112 25872 25140
rect 24811 25109 24823 25112
rect 24765 25103 24823 25109
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 26988 25140 27016 25248
rect 27065 25245 27077 25279
rect 27111 25276 27123 25279
rect 32033 25279 32091 25285
rect 27111 25248 27568 25276
rect 27111 25245 27123 25248
rect 27065 25239 27123 25245
rect 27540 25220 27568 25248
rect 32033 25245 32045 25279
rect 32079 25276 32091 25279
rect 32858 25276 32864 25288
rect 32079 25248 32864 25276
rect 32079 25245 32091 25248
rect 32033 25239 32091 25245
rect 32858 25236 32864 25248
rect 32916 25236 32922 25288
rect 36924 25276 36952 25375
rect 37274 25372 37280 25384
rect 37332 25372 37338 25424
rect 35912 25248 36952 25276
rect 35912 25220 35940 25248
rect 37182 25236 37188 25288
rect 37240 25276 37246 25288
rect 37369 25279 37427 25285
rect 37369 25276 37381 25279
rect 37240 25248 37381 25276
rect 37240 25236 37246 25248
rect 37369 25245 37381 25248
rect 37415 25245 37427 25279
rect 37369 25239 37427 25245
rect 37458 25236 37464 25288
rect 37516 25276 37522 25288
rect 37752 25285 37780 25452
rect 37737 25279 37795 25285
rect 37516 25248 37561 25276
rect 37516 25236 37522 25248
rect 37737 25245 37749 25279
rect 37783 25245 37795 25279
rect 37737 25239 37795 25245
rect 37826 25236 37832 25288
rect 37884 25285 37890 25288
rect 37884 25276 37892 25285
rect 37884 25248 37929 25276
rect 37884 25239 37892 25248
rect 37884 25236 37890 25239
rect 27338 25217 27344 25220
rect 27310 25211 27344 25217
rect 27310 25177 27322 25211
rect 27310 25171 27344 25177
rect 27338 25168 27344 25171
rect 27396 25168 27402 25220
rect 27522 25168 27528 25220
rect 27580 25168 27586 25220
rect 31941 25211 31999 25217
rect 31941 25208 31953 25211
rect 30484 25180 31953 25208
rect 30484 25152 30512 25180
rect 31941 25177 31953 25180
rect 31987 25177 31999 25211
rect 31941 25171 31999 25177
rect 35526 25168 35532 25220
rect 35584 25208 35590 25220
rect 35774 25211 35832 25217
rect 35774 25208 35786 25211
rect 35584 25180 35786 25208
rect 35584 25168 35590 25180
rect 35774 25177 35786 25180
rect 35820 25177 35832 25211
rect 35774 25171 35832 25177
rect 35894 25168 35900 25220
rect 35952 25168 35958 25220
rect 36538 25168 36544 25220
rect 36596 25208 36602 25220
rect 36998 25208 37004 25220
rect 36596 25180 37004 25208
rect 36596 25168 36602 25180
rect 36998 25168 37004 25180
rect 37056 25208 37062 25220
rect 37645 25211 37703 25217
rect 37645 25208 37657 25211
rect 37056 25180 37657 25208
rect 37056 25168 37062 25180
rect 37645 25177 37657 25180
rect 37691 25177 37703 25211
rect 37645 25171 37703 25177
rect 30466 25140 30472 25152
rect 26292 25112 26337 25140
rect 26988 25112 30472 25140
rect 26292 25100 26298 25112
rect 30466 25100 30472 25112
rect 30524 25100 30530 25152
rect 30561 25143 30619 25149
rect 30561 25109 30573 25143
rect 30607 25140 30619 25143
rect 31113 25143 31171 25149
rect 31113 25140 31125 25143
rect 30607 25112 31125 25140
rect 30607 25109 30619 25112
rect 30561 25103 30619 25109
rect 31113 25109 31125 25112
rect 31159 25140 31171 25143
rect 31294 25140 31300 25152
rect 31159 25112 31300 25140
rect 31159 25109 31171 25112
rect 31113 25103 31171 25109
rect 31294 25100 31300 25112
rect 31352 25100 31358 25152
rect 32766 25140 32772 25152
rect 32727 25112 32772 25140
rect 32766 25100 32772 25112
rect 32824 25100 32830 25152
rect 37274 25100 37280 25152
rect 37332 25140 37338 25152
rect 38013 25143 38071 25149
rect 38013 25140 38025 25143
rect 37332 25112 38025 25140
rect 37332 25100 37338 25112
rect 38013 25109 38025 25112
rect 38059 25109 38071 25143
rect 38013 25103 38071 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 26973 24939 27031 24945
rect 26973 24905 26985 24939
rect 27019 24936 27031 24939
rect 27062 24936 27068 24948
rect 27019 24908 27068 24936
rect 27019 24905 27031 24908
rect 26973 24899 27031 24905
rect 27062 24896 27068 24908
rect 27120 24896 27126 24948
rect 27341 24939 27399 24945
rect 27341 24905 27353 24939
rect 27387 24936 27399 24939
rect 27706 24936 27712 24948
rect 27387 24908 27712 24936
rect 27387 24905 27399 24908
rect 27341 24899 27399 24905
rect 27706 24896 27712 24908
rect 27764 24936 27770 24948
rect 28258 24936 28264 24948
rect 27764 24908 28264 24936
rect 27764 24896 27770 24908
rect 28258 24896 28264 24908
rect 28316 24896 28322 24948
rect 25866 24828 25872 24880
rect 25924 24868 25930 24880
rect 32766 24868 32772 24880
rect 25924 24840 32772 24868
rect 25924 24828 25930 24840
rect 32766 24828 32772 24840
rect 32824 24828 32830 24880
rect 1854 24800 1860 24812
rect 1815 24772 1860 24800
rect 1854 24760 1860 24772
rect 1912 24800 1918 24812
rect 2685 24803 2743 24809
rect 2685 24800 2697 24803
rect 1912 24772 2697 24800
rect 1912 24760 1918 24772
rect 2685 24769 2697 24772
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24769 23443 24803
rect 23385 24763 23443 24769
rect 23569 24803 23627 24809
rect 23569 24769 23581 24803
rect 23615 24800 23627 24803
rect 23842 24800 23848 24812
rect 23615 24772 23848 24800
rect 23615 24769 23627 24772
rect 23569 24763 23627 24769
rect 23400 24732 23428 24763
rect 23842 24760 23848 24772
rect 23900 24760 23906 24812
rect 26234 24760 26240 24812
rect 26292 24800 26298 24812
rect 27433 24803 27491 24809
rect 26292 24772 26337 24800
rect 26292 24760 26298 24772
rect 27433 24769 27445 24803
rect 27479 24800 27491 24803
rect 28350 24800 28356 24812
rect 27479 24772 28356 24800
rect 27479 24769 27491 24772
rect 27433 24763 27491 24769
rect 23658 24732 23664 24744
rect 23400 24704 23664 24732
rect 23658 24692 23664 24704
rect 23716 24732 23722 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 23716 24704 24593 24732
rect 23716 24692 23722 24704
rect 24581 24701 24593 24704
rect 24627 24701 24639 24735
rect 24581 24695 24639 24701
rect 24854 24692 24860 24744
rect 24912 24732 24918 24744
rect 27448 24732 27476 24763
rect 28350 24760 28356 24772
rect 28408 24800 28414 24812
rect 28721 24803 28779 24809
rect 28721 24800 28733 24803
rect 28408 24772 28733 24800
rect 28408 24760 28414 24772
rect 28721 24769 28733 24772
rect 28767 24769 28779 24803
rect 28721 24763 28779 24769
rect 30466 24760 30472 24812
rect 30524 24800 30530 24812
rect 31389 24803 31447 24809
rect 31389 24800 31401 24803
rect 30524 24772 31401 24800
rect 30524 24760 30530 24772
rect 31389 24769 31401 24772
rect 31435 24769 31447 24803
rect 35342 24800 35348 24812
rect 35303 24772 35348 24800
rect 31389 24763 31447 24769
rect 35342 24760 35348 24772
rect 35400 24760 35406 24812
rect 35612 24803 35670 24809
rect 35612 24769 35624 24803
rect 35658 24800 35670 24803
rect 35986 24800 35992 24812
rect 35658 24772 35992 24800
rect 35658 24769 35670 24772
rect 35612 24763 35670 24769
rect 35986 24760 35992 24772
rect 36044 24760 36050 24812
rect 37550 24760 37556 24812
rect 37608 24800 37614 24812
rect 37829 24803 37887 24809
rect 37829 24800 37841 24803
rect 37608 24772 37841 24800
rect 37608 24760 37614 24772
rect 37829 24769 37841 24772
rect 37875 24769 37887 24803
rect 37829 24763 37887 24769
rect 24912 24704 27476 24732
rect 27525 24735 27583 24741
rect 24912 24692 24918 24704
rect 27525 24701 27537 24735
rect 27571 24701 27583 24735
rect 28258 24732 28264 24744
rect 28171 24704 28264 24732
rect 27525 24695 27583 24701
rect 2133 24667 2191 24673
rect 2133 24633 2145 24667
rect 2179 24664 2191 24667
rect 21634 24664 21640 24676
rect 2179 24636 21640 24664
rect 2179 24633 2191 24636
rect 2133 24627 2191 24633
rect 21634 24624 21640 24636
rect 21692 24624 21698 24676
rect 22741 24667 22799 24673
rect 22741 24633 22753 24667
rect 22787 24664 22799 24667
rect 23014 24664 23020 24676
rect 22787 24636 23020 24664
rect 22787 24633 22799 24636
rect 22741 24627 22799 24633
rect 23014 24624 23020 24636
rect 23072 24624 23078 24676
rect 26326 24624 26332 24676
rect 26384 24664 26390 24676
rect 27154 24664 27160 24676
rect 26384 24636 27160 24664
rect 26384 24624 26390 24636
rect 27154 24624 27160 24636
rect 27212 24664 27218 24676
rect 27540 24664 27568 24695
rect 28258 24692 28264 24704
rect 28316 24732 28322 24744
rect 30374 24732 30380 24744
rect 28316 24704 30380 24732
rect 28316 24692 28322 24704
rect 30374 24692 30380 24704
rect 30432 24692 30438 24744
rect 37458 24732 37464 24744
rect 36740 24704 37464 24732
rect 36740 24673 36768 24704
rect 37458 24692 37464 24704
rect 37516 24732 37522 24744
rect 38102 24732 38108 24744
rect 37516 24704 38108 24732
rect 37516 24692 37522 24704
rect 38102 24692 38108 24704
rect 38160 24692 38166 24744
rect 27212 24636 27568 24664
rect 36725 24667 36783 24673
rect 27212 24624 27218 24636
rect 36725 24633 36737 24667
rect 36771 24633 36783 24667
rect 38010 24664 38016 24676
rect 37971 24636 38016 24664
rect 36725 24627 36783 24633
rect 38010 24624 38016 24636
rect 38068 24624 38074 24676
rect 22189 24599 22247 24605
rect 22189 24565 22201 24599
rect 22235 24596 22247 24599
rect 22462 24596 22468 24608
rect 22235 24568 22468 24596
rect 22235 24565 22247 24568
rect 22189 24559 22247 24565
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 22830 24556 22836 24608
rect 22888 24596 22894 24608
rect 23201 24599 23259 24605
rect 23201 24596 23213 24599
rect 22888 24568 23213 24596
rect 22888 24556 22894 24568
rect 23201 24565 23213 24568
rect 23247 24565 23259 24599
rect 23201 24559 23259 24565
rect 23842 24556 23848 24608
rect 23900 24596 23906 24608
rect 24029 24599 24087 24605
rect 24029 24596 24041 24599
rect 23900 24568 24041 24596
rect 23900 24556 23906 24568
rect 24029 24565 24041 24568
rect 24075 24596 24087 24599
rect 25133 24599 25191 24605
rect 25133 24596 25145 24599
rect 24075 24568 25145 24596
rect 24075 24565 24087 24568
rect 24029 24559 24087 24565
rect 25133 24565 25145 24568
rect 25179 24565 25191 24599
rect 25133 24559 25191 24565
rect 26421 24599 26479 24605
rect 26421 24565 26433 24599
rect 26467 24596 26479 24599
rect 27338 24596 27344 24608
rect 26467 24568 27344 24596
rect 26467 24565 26479 24568
rect 26421 24559 26479 24565
rect 27338 24556 27344 24568
rect 27396 24556 27402 24608
rect 32493 24599 32551 24605
rect 32493 24565 32505 24599
rect 32539 24596 32551 24599
rect 32582 24596 32588 24608
rect 32539 24568 32588 24596
rect 32539 24565 32551 24568
rect 32493 24559 32551 24565
rect 32582 24556 32588 24568
rect 32640 24556 32646 24608
rect 37182 24556 37188 24608
rect 37240 24596 37246 24608
rect 37277 24599 37335 24605
rect 37277 24596 37289 24599
rect 37240 24568 37289 24596
rect 37240 24556 37246 24568
rect 37277 24565 37289 24568
rect 37323 24565 37335 24599
rect 37277 24559 37335 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1486 24392 1492 24404
rect 1447 24364 1492 24392
rect 1486 24352 1492 24364
rect 1544 24352 1550 24404
rect 24486 24392 24492 24404
rect 24447 24364 24492 24392
rect 24486 24352 24492 24364
rect 24544 24352 24550 24404
rect 27157 24395 27215 24401
rect 27157 24361 27169 24395
rect 27203 24392 27215 24395
rect 28074 24392 28080 24404
rect 27203 24364 28080 24392
rect 27203 24361 27215 24364
rect 27157 24355 27215 24361
rect 28074 24352 28080 24364
rect 28132 24352 28138 24404
rect 35526 24392 35532 24404
rect 35487 24364 35532 24392
rect 35526 24352 35532 24364
rect 35584 24352 35590 24404
rect 35986 24392 35992 24404
rect 35947 24364 35992 24392
rect 35986 24352 35992 24364
rect 36044 24352 36050 24404
rect 36262 24352 36268 24404
rect 36320 24392 36326 24404
rect 36725 24395 36783 24401
rect 36725 24392 36737 24395
rect 36320 24364 36737 24392
rect 36320 24352 36326 24364
rect 36725 24361 36737 24364
rect 36771 24392 36783 24395
rect 37182 24392 37188 24404
rect 36771 24364 37188 24392
rect 36771 24361 36783 24364
rect 36725 24355 36783 24361
rect 37182 24352 37188 24364
rect 37240 24352 37246 24404
rect 2222 24284 2228 24336
rect 2280 24324 2286 24336
rect 22097 24327 22155 24333
rect 22097 24324 22109 24327
rect 2280 24296 22109 24324
rect 2280 24284 2286 24296
rect 22097 24293 22109 24296
rect 22143 24293 22155 24327
rect 22097 24287 22155 24293
rect 23566 24284 23572 24336
rect 23624 24324 23630 24336
rect 24949 24327 25007 24333
rect 24949 24324 24961 24327
rect 23624 24296 24961 24324
rect 23624 24284 23630 24296
rect 24949 24293 24961 24296
rect 24995 24293 25007 24327
rect 27062 24324 27068 24336
rect 27023 24296 27068 24324
rect 24949 24287 25007 24293
rect 27062 24284 27068 24296
rect 27120 24284 27126 24336
rect 27890 24324 27896 24336
rect 27803 24296 27896 24324
rect 27890 24284 27896 24296
rect 27948 24324 27954 24336
rect 28442 24324 28448 24336
rect 27948 24296 28448 24324
rect 27948 24284 27954 24296
rect 28442 24284 28448 24296
rect 28500 24284 28506 24336
rect 37274 24324 37280 24336
rect 31036 24296 37280 24324
rect 2682 24256 2688 24268
rect 1688 24228 2688 24256
rect 1688 24197 1716 24228
rect 2682 24216 2688 24228
rect 2740 24256 2746 24268
rect 22646 24256 22652 24268
rect 2740 24228 22652 24256
rect 2740 24216 2746 24228
rect 22646 24216 22652 24228
rect 22704 24216 22710 24268
rect 22830 24256 22836 24268
rect 22791 24228 22836 24256
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 26697 24259 26755 24265
rect 26697 24225 26709 24259
rect 26743 24256 26755 24259
rect 27430 24256 27436 24268
rect 26743 24228 27436 24256
rect 26743 24225 26755 24228
rect 26697 24219 26755 24225
rect 27430 24216 27436 24228
rect 27488 24216 27494 24268
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24157 1731 24191
rect 2130 24188 2136 24200
rect 2091 24160 2136 24188
rect 1673 24151 1731 24157
rect 2130 24148 2136 24160
rect 2188 24188 2194 24200
rect 2777 24191 2835 24197
rect 2777 24188 2789 24191
rect 2188 24160 2789 24188
rect 2188 24148 2194 24160
rect 2777 24157 2789 24160
rect 2823 24157 2835 24191
rect 2777 24151 2835 24157
rect 22537 24191 22595 24197
rect 22537 24157 22549 24191
rect 22583 24188 22595 24191
rect 22741 24191 22799 24197
rect 22583 24160 22692 24188
rect 22583 24157 22595 24160
rect 22537 24151 22595 24157
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 22281 24123 22339 24129
rect 22281 24120 22293 24123
rect 21876 24092 22293 24120
rect 21876 24080 21882 24092
rect 22281 24089 22293 24092
rect 22327 24089 22339 24123
rect 22664 24120 22692 24160
rect 22741 24157 22753 24191
rect 22787 24188 22799 24191
rect 31036 24188 31064 24296
rect 37274 24284 37280 24296
rect 37332 24284 37338 24336
rect 37369 24327 37427 24333
rect 37369 24293 37381 24327
rect 37415 24324 37427 24327
rect 37826 24324 37832 24336
rect 37415 24296 37832 24324
rect 37415 24293 37427 24296
rect 37369 24287 37427 24293
rect 37826 24284 37832 24296
rect 37884 24324 37890 24336
rect 38286 24324 38292 24336
rect 37884 24296 38292 24324
rect 37884 24284 37890 24296
rect 38286 24284 38292 24296
rect 38344 24284 38350 24336
rect 36722 24256 36728 24268
rect 22787 24160 31064 24188
rect 31128 24228 36728 24256
rect 22787 24157 22799 24160
rect 22741 24151 22799 24157
rect 23014 24120 23020 24132
rect 22664 24092 23020 24120
rect 22281 24083 22339 24089
rect 23014 24080 23020 24092
rect 23072 24080 23078 24132
rect 23661 24123 23719 24129
rect 23661 24089 23673 24123
rect 23707 24089 23719 24123
rect 23842 24120 23848 24132
rect 23803 24092 23848 24120
rect 23661 24083 23719 24089
rect 2317 24055 2375 24061
rect 2317 24021 2329 24055
rect 2363 24052 2375 24055
rect 2406 24052 2412 24064
rect 2363 24024 2412 24052
rect 2363 24021 2375 24024
rect 2317 24015 2375 24021
rect 2406 24012 2412 24024
rect 2464 24012 2470 24064
rect 22554 24012 22560 24064
rect 22612 24052 22618 24064
rect 22649 24055 22707 24061
rect 22649 24052 22661 24055
rect 22612 24024 22661 24052
rect 22612 24012 22618 24024
rect 22649 24021 22661 24024
rect 22695 24021 22707 24055
rect 23474 24052 23480 24064
rect 23435 24024 23480 24052
rect 22649 24015 22707 24021
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 23676 24052 23704 24083
rect 23842 24080 23848 24092
rect 23900 24080 23906 24132
rect 28902 24080 28908 24132
rect 28960 24120 28966 24132
rect 31128 24120 31156 24228
rect 36722 24216 36728 24228
rect 36780 24216 36786 24268
rect 34514 24148 34520 24200
rect 34572 24188 34578 24200
rect 35345 24191 35403 24197
rect 35345 24188 35357 24191
rect 34572 24160 35357 24188
rect 34572 24148 34578 24160
rect 35345 24157 35357 24160
rect 35391 24157 35403 24191
rect 36170 24188 36176 24200
rect 36131 24160 36176 24188
rect 35345 24151 35403 24157
rect 36170 24148 36176 24160
rect 36228 24148 36234 24200
rect 37366 24188 37372 24200
rect 36556 24160 37372 24188
rect 36556 24120 36584 24160
rect 37366 24148 37372 24160
rect 37424 24148 37430 24200
rect 37829 24191 37887 24197
rect 37829 24157 37841 24191
rect 37875 24157 37887 24191
rect 37829 24151 37887 24157
rect 37844 24120 37872 24151
rect 28960 24092 31156 24120
rect 31211 24092 36584 24120
rect 36648 24092 37872 24120
rect 28960 24080 28966 24092
rect 24486 24052 24492 24064
rect 23676 24024 24492 24052
rect 24486 24012 24492 24024
rect 24544 24012 24550 24064
rect 27154 24012 27160 24064
rect 27212 24052 27218 24064
rect 28353 24055 28411 24061
rect 28353 24052 28365 24055
rect 27212 24024 28365 24052
rect 27212 24012 27218 24024
rect 28353 24021 28365 24024
rect 28399 24021 28411 24055
rect 28353 24015 28411 24021
rect 28626 24012 28632 24064
rect 28684 24052 28690 24064
rect 31211 24052 31239 24092
rect 28684 24024 31239 24052
rect 28684 24012 28690 24024
rect 31386 24012 31392 24064
rect 31444 24052 31450 24064
rect 36648 24052 36676 24092
rect 38010 24052 38016 24064
rect 31444 24024 36676 24052
rect 37971 24024 38016 24052
rect 31444 24012 31450 24024
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 22646 23848 22652 23860
rect 22607 23820 22652 23848
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 24946 23808 24952 23860
rect 25004 23848 25010 23860
rect 27433 23851 27491 23857
rect 27433 23848 27445 23851
rect 25004 23820 27445 23848
rect 25004 23808 25010 23820
rect 27433 23817 27445 23820
rect 27479 23848 27491 23851
rect 27890 23848 27896 23860
rect 27479 23820 27896 23848
rect 27479 23817 27491 23820
rect 27433 23811 27491 23817
rect 27890 23808 27896 23820
rect 27948 23808 27954 23860
rect 28994 23808 29000 23860
rect 29052 23848 29058 23860
rect 31386 23848 31392 23860
rect 29052 23820 31392 23848
rect 29052 23808 29058 23820
rect 31386 23808 31392 23820
rect 31444 23808 31450 23860
rect 22373 23783 22431 23789
rect 22373 23749 22385 23783
rect 22419 23780 22431 23783
rect 36078 23780 36084 23792
rect 22419 23752 36084 23780
rect 22419 23749 22431 23752
rect 22373 23743 22431 23749
rect 36078 23740 36084 23752
rect 36136 23740 36142 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23681 1731 23715
rect 2406 23712 2412 23724
rect 2367 23684 2412 23712
rect 1673 23675 1731 23681
rect 1688 23644 1716 23675
rect 2406 23672 2412 23684
rect 2464 23672 2470 23724
rect 2498 23672 2504 23724
rect 2556 23712 2562 23724
rect 2866 23712 2872 23724
rect 2556 23684 2601 23712
rect 2827 23684 2872 23712
rect 2556 23672 2562 23684
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 22094 23672 22100 23724
rect 22152 23721 22158 23724
rect 22152 23715 22201 23721
rect 22152 23681 22155 23715
rect 22189 23681 22201 23715
rect 22152 23675 22201 23681
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 22465 23715 22523 23721
rect 22465 23681 22477 23715
rect 22511 23712 22523 23715
rect 23293 23715 23351 23721
rect 23293 23712 23305 23715
rect 22511 23684 23305 23712
rect 22511 23681 22523 23684
rect 22465 23675 22523 23681
rect 23293 23681 23305 23684
rect 23339 23681 23351 23715
rect 23293 23675 23351 23681
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 23566 23712 23572 23724
rect 23523 23684 23572 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 22152 23672 22158 23675
rect 1688 23616 3648 23644
rect 3620 23520 3648 23616
rect 21634 23604 21640 23656
rect 21692 23644 21698 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21692 23616 22017 23644
rect 21692 23604 21698 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22296 23644 22324 23675
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 23661 23715 23719 23721
rect 23661 23681 23673 23715
rect 23707 23712 23719 23715
rect 23842 23712 23848 23724
rect 23707 23684 23848 23712
rect 23707 23681 23719 23684
rect 23661 23675 23719 23681
rect 23842 23672 23848 23684
rect 23900 23712 23906 23724
rect 25038 23712 25044 23724
rect 23900 23684 25044 23712
rect 23900 23672 23906 23684
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23712 26479 23715
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 26467 23684 27353 23712
rect 26467 23681 26479 23684
rect 26421 23675 26479 23681
rect 27341 23681 27353 23684
rect 27387 23712 27399 23715
rect 34146 23712 34152 23724
rect 27387 23684 34152 23712
rect 27387 23681 27399 23684
rect 27341 23675 27399 23681
rect 22646 23644 22652 23656
rect 22296 23616 22652 23644
rect 22005 23607 22063 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 23584 23644 23612 23672
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 23584 23616 24133 23644
rect 24121 23613 24133 23616
rect 24167 23613 24179 23647
rect 24121 23607 24179 23613
rect 16942 23536 16948 23588
rect 17000 23576 17006 23588
rect 26436 23576 26464 23675
rect 34146 23672 34152 23684
rect 34204 23672 34210 23724
rect 37461 23715 37519 23721
rect 37461 23681 37473 23715
rect 37507 23712 37519 23715
rect 38102 23712 38108 23724
rect 37507 23684 38108 23712
rect 37507 23681 37519 23684
rect 37461 23675 37519 23681
rect 38102 23672 38108 23684
rect 38160 23672 38166 23724
rect 27525 23647 27583 23653
rect 27525 23613 27537 23647
rect 27571 23613 27583 23647
rect 27525 23607 27583 23613
rect 28261 23647 28319 23653
rect 28261 23613 28273 23647
rect 28307 23644 28319 23647
rect 28810 23644 28816 23656
rect 28307 23616 28816 23644
rect 28307 23613 28319 23616
rect 28261 23607 28319 23613
rect 17000 23548 26464 23576
rect 17000 23536 17006 23548
rect 27338 23536 27344 23588
rect 27396 23576 27402 23588
rect 27540 23576 27568 23607
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 27396 23548 27568 23576
rect 27396 23536 27402 23548
rect 27614 23536 27620 23588
rect 27672 23576 27678 23588
rect 27672 23548 28764 23576
rect 27672 23536 27678 23548
rect 28736 23520 28764 23548
rect 1486 23508 1492 23520
rect 1447 23480 1492 23508
rect 1486 23468 1492 23480
rect 1544 23468 1550 23520
rect 2774 23508 2780 23520
rect 2735 23480 2780 23508
rect 2774 23468 2780 23480
rect 2832 23468 2838 23520
rect 3053 23511 3111 23517
rect 3053 23477 3065 23511
rect 3099 23508 3111 23511
rect 3326 23508 3332 23520
rect 3099 23480 3332 23508
rect 3099 23477 3111 23480
rect 3053 23471 3111 23477
rect 3326 23468 3332 23480
rect 3384 23468 3390 23520
rect 3602 23508 3608 23520
rect 3563 23480 3608 23508
rect 3602 23468 3608 23480
rect 3660 23468 3666 23520
rect 26878 23468 26884 23520
rect 26936 23508 26942 23520
rect 26973 23511 27031 23517
rect 26973 23508 26985 23511
rect 26936 23480 26985 23508
rect 26936 23468 26942 23480
rect 26973 23477 26985 23480
rect 27019 23477 27031 23511
rect 28718 23508 28724 23520
rect 28679 23480 28724 23508
rect 26973 23471 27031 23477
rect 28718 23468 28724 23480
rect 28776 23468 28782 23520
rect 37826 23468 37832 23520
rect 37884 23508 37890 23520
rect 37921 23511 37979 23517
rect 37921 23508 37933 23511
rect 37884 23480 37933 23508
rect 37884 23468 37890 23480
rect 37921 23477 37933 23480
rect 37967 23477 37979 23511
rect 37921 23471 37979 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 24581 23307 24639 23313
rect 24581 23273 24593 23307
rect 24627 23304 24639 23307
rect 24854 23304 24860 23316
rect 24627 23276 24860 23304
rect 24627 23273 24639 23276
rect 24581 23267 24639 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 26234 23264 26240 23316
rect 26292 23304 26298 23316
rect 26697 23307 26755 23313
rect 26697 23304 26709 23307
rect 26292 23276 26709 23304
rect 26292 23264 26298 23276
rect 26697 23273 26709 23276
rect 26743 23273 26755 23307
rect 26697 23267 26755 23273
rect 28997 23307 29055 23313
rect 28997 23273 29009 23307
rect 29043 23304 29055 23307
rect 29454 23304 29460 23316
rect 29043 23276 29460 23304
rect 29043 23273 29055 23276
rect 28997 23267 29055 23273
rect 29454 23264 29460 23276
rect 29512 23304 29518 23316
rect 33686 23304 33692 23316
rect 29512 23276 33692 23304
rect 29512 23264 29518 23276
rect 33686 23264 33692 23276
rect 33744 23264 33750 23316
rect 35161 23307 35219 23313
rect 35161 23273 35173 23307
rect 35207 23304 35219 23307
rect 36170 23304 36176 23316
rect 35207 23276 36176 23304
rect 35207 23273 35219 23276
rect 35161 23267 35219 23273
rect 36170 23264 36176 23276
rect 36228 23264 36234 23316
rect 24394 23236 24400 23248
rect 6886 23208 24400 23236
rect 2133 23171 2191 23177
rect 2133 23137 2145 23171
rect 2179 23168 2191 23171
rect 6886 23168 6914 23208
rect 24394 23196 24400 23208
rect 24452 23196 24458 23248
rect 26878 23236 26884 23248
rect 26839 23208 26884 23236
rect 26878 23196 26884 23208
rect 26936 23196 26942 23248
rect 35066 23236 35072 23248
rect 35027 23208 35072 23236
rect 35066 23196 35072 23208
rect 35124 23196 35130 23248
rect 23474 23168 23480 23180
rect 2179 23140 6914 23168
rect 22480 23140 23480 23168
rect 2179 23137 2191 23140
rect 2133 23131 2191 23137
rect 22480 23109 22508 23140
rect 23474 23128 23480 23140
rect 23532 23128 23538 23180
rect 26234 23128 26240 23180
rect 26292 23168 26298 23180
rect 27157 23171 27215 23177
rect 27157 23168 27169 23171
rect 26292 23140 27169 23168
rect 26292 23128 26298 23140
rect 27157 23137 27169 23140
rect 27203 23168 27215 23171
rect 27430 23168 27436 23180
rect 27203 23140 27436 23168
rect 27203 23137 27215 23140
rect 27157 23131 27215 23137
rect 27430 23128 27436 23140
rect 27488 23128 27494 23180
rect 27614 23168 27620 23180
rect 27575 23140 27620 23168
rect 27614 23128 27620 23140
rect 27672 23128 27678 23180
rect 22465 23103 22523 23109
rect 22465 23069 22477 23103
rect 22511 23069 22523 23103
rect 22922 23100 22928 23112
rect 22883 23072 22928 23100
rect 22465 23063 22523 23069
rect 22922 23060 22928 23072
rect 22980 23060 22986 23112
rect 28902 23100 28908 23112
rect 26206 23072 28908 23100
rect 1854 23032 1860 23044
rect 1815 23004 1860 23032
rect 1854 22992 1860 23004
rect 1912 23032 1918 23044
rect 2685 23035 2743 23041
rect 2685 23032 2697 23035
rect 1912 23004 2697 23032
rect 1912 22992 1918 23004
rect 2685 23001 2697 23004
rect 2731 23001 2743 23035
rect 2685 22995 2743 23001
rect 3602 22992 3608 23044
rect 3660 23032 3666 23044
rect 22281 23035 22339 23041
rect 22281 23032 22293 23035
rect 3660 23004 22293 23032
rect 3660 22992 3666 23004
rect 22281 23001 22293 23004
rect 22327 23001 22339 23035
rect 22281 22995 22339 23001
rect 22557 23035 22615 23041
rect 22557 23001 22569 23035
rect 22603 23001 22615 23035
rect 22557 22995 22615 23001
rect 22572 22964 22600 22995
rect 22646 22992 22652 23044
rect 22704 23032 22710 23044
rect 22787 23035 22845 23041
rect 22704 23004 22749 23032
rect 22704 22992 22710 23004
rect 22787 23001 22799 23035
rect 22833 23032 22845 23035
rect 23198 23032 23204 23044
rect 22833 23004 23204 23032
rect 22833 23001 22845 23004
rect 22787 22995 22845 23001
rect 23198 22992 23204 23004
rect 23256 22992 23262 23044
rect 26206 23032 26234 23072
rect 28902 23060 28908 23072
rect 28960 23060 28966 23112
rect 31386 23100 31392 23112
rect 31347 23072 31392 23100
rect 31386 23060 31392 23072
rect 31444 23060 31450 23112
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23100 37887 23103
rect 37918 23100 37924 23112
rect 37875 23072 37924 23100
rect 37875 23069 37887 23072
rect 37829 23063 37887 23069
rect 37918 23060 37924 23072
rect 37976 23060 37982 23112
rect 23676 23004 26234 23032
rect 23676 22964 23704 23004
rect 27246 22992 27252 23044
rect 27304 23032 27310 23044
rect 27862 23035 27920 23041
rect 27862 23032 27874 23035
rect 27304 23004 27874 23032
rect 27304 22992 27310 23004
rect 27862 23001 27874 23004
rect 27908 23001 27920 23035
rect 27862 22995 27920 23001
rect 31478 22992 31484 23044
rect 31536 23032 31542 23044
rect 31634 23035 31692 23041
rect 31634 23032 31646 23035
rect 31536 23004 31646 23032
rect 31536 22992 31542 23004
rect 31634 23001 31646 23004
rect 31680 23001 31692 23035
rect 31634 22995 31692 23001
rect 34606 22992 34612 23044
rect 34664 23032 34670 23044
rect 34701 23035 34759 23041
rect 34701 23032 34713 23035
rect 34664 23004 34713 23032
rect 34664 22992 34670 23004
rect 34701 23001 34713 23004
rect 34747 23001 34759 23035
rect 34701 22995 34759 23001
rect 22572 22936 23704 22964
rect 23845 22967 23903 22973
rect 23845 22933 23857 22967
rect 23891 22964 23903 22967
rect 25038 22964 25044 22976
rect 23891 22936 25044 22964
rect 23891 22933 23903 22936
rect 23845 22927 23903 22933
rect 25038 22924 25044 22936
rect 25096 22924 25102 22976
rect 26786 22924 26792 22976
rect 26844 22964 26850 22976
rect 27614 22964 27620 22976
rect 26844 22936 27620 22964
rect 26844 22924 26850 22936
rect 27614 22924 27620 22936
rect 27672 22924 27678 22976
rect 32766 22964 32772 22976
rect 32679 22936 32772 22964
rect 32766 22924 32772 22936
rect 32824 22964 32830 22976
rect 37550 22964 37556 22976
rect 32824 22936 37556 22964
rect 32824 22924 32830 22936
rect 37550 22924 37556 22936
rect 37608 22924 37614 22976
rect 38010 22964 38016 22976
rect 37971 22936 38016 22964
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2317 22763 2375 22769
rect 2317 22729 2329 22763
rect 2363 22760 2375 22763
rect 2498 22760 2504 22772
rect 2363 22732 2504 22760
rect 2363 22729 2375 22732
rect 2317 22723 2375 22729
rect 2498 22720 2504 22732
rect 2556 22720 2562 22772
rect 24946 22760 24952 22772
rect 24907 22732 24952 22760
rect 24946 22720 24952 22732
rect 25004 22720 25010 22772
rect 26421 22763 26479 22769
rect 26421 22729 26433 22763
rect 26467 22760 26479 22763
rect 27246 22760 27252 22772
rect 26467 22732 27252 22760
rect 26467 22729 26479 22732
rect 26421 22723 26479 22729
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 27341 22763 27399 22769
rect 27341 22729 27353 22763
rect 27387 22760 27399 22763
rect 27614 22760 27620 22772
rect 27387 22732 27620 22760
rect 27387 22729 27399 22732
rect 27341 22723 27399 22729
rect 27614 22720 27620 22732
rect 27672 22760 27678 22772
rect 29454 22760 29460 22772
rect 27672 22732 29460 22760
rect 27672 22720 27678 22732
rect 29454 22720 29460 22732
rect 29512 22720 29518 22772
rect 31478 22760 31484 22772
rect 31439 22732 31484 22760
rect 31478 22720 31484 22732
rect 31536 22720 31542 22772
rect 34149 22763 34207 22769
rect 34149 22729 34161 22763
rect 34195 22760 34207 22763
rect 34514 22760 34520 22772
rect 34195 22732 34520 22760
rect 34195 22729 34207 22732
rect 34149 22723 34207 22729
rect 34514 22720 34520 22732
rect 34572 22720 34578 22772
rect 34885 22763 34943 22769
rect 34885 22729 34897 22763
rect 34931 22760 34943 22763
rect 37458 22760 37464 22772
rect 34931 22732 37464 22760
rect 34931 22729 34943 22732
rect 34885 22723 34943 22729
rect 37458 22720 37464 22732
rect 37516 22760 37522 22772
rect 38378 22760 38384 22772
rect 37516 22732 38384 22760
rect 37516 22720 37522 22732
rect 38378 22720 38384 22732
rect 38436 22720 38442 22772
rect 24213 22695 24271 22701
rect 24213 22661 24225 22695
rect 24259 22692 24271 22695
rect 24854 22692 24860 22704
rect 24259 22664 24860 22692
rect 24259 22661 24271 22664
rect 24213 22655 24271 22661
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 28258 22692 28264 22704
rect 26252 22664 28264 22692
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22593 1731 22627
rect 2130 22624 2136 22636
rect 2091 22596 2136 22624
rect 1673 22587 1731 22593
rect 1688 22556 1716 22587
rect 2130 22584 2136 22596
rect 2188 22624 2194 22636
rect 2777 22627 2835 22633
rect 2777 22624 2789 22627
rect 2188 22596 2789 22624
rect 2188 22584 2194 22596
rect 2777 22593 2789 22596
rect 2823 22593 2835 22627
rect 24394 22624 24400 22636
rect 24355 22596 24400 22624
rect 2777 22587 2835 22593
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 26252 22633 26280 22664
rect 28258 22652 28264 22664
rect 28316 22652 28322 22704
rect 33962 22692 33968 22704
rect 28552 22664 33968 22692
rect 26237 22627 26295 22633
rect 26237 22593 26249 22627
rect 26283 22593 26295 22627
rect 27433 22627 27491 22633
rect 27433 22624 27445 22627
rect 26237 22587 26295 22593
rect 26988 22596 27445 22624
rect 1688 22528 3464 22556
rect 3436 22432 3464 22528
rect 25222 22516 25228 22568
rect 25280 22556 25286 22568
rect 26786 22556 26792 22568
rect 25280 22528 26792 22556
rect 25280 22516 25286 22528
rect 26786 22516 26792 22528
rect 26844 22516 26850 22568
rect 26988 22488 27016 22596
rect 27433 22593 27445 22596
rect 27479 22624 27491 22627
rect 28552 22624 28580 22664
rect 33962 22652 33968 22664
rect 34020 22652 34026 22704
rect 37366 22652 37372 22704
rect 37424 22692 37430 22704
rect 37645 22695 37703 22701
rect 37645 22692 37657 22695
rect 37424 22664 37657 22692
rect 37424 22652 37430 22664
rect 37645 22661 37657 22664
rect 37691 22661 37703 22695
rect 37645 22655 37703 22661
rect 27479 22596 28580 22624
rect 28629 22627 28687 22633
rect 27479 22593 27491 22596
rect 27433 22587 27491 22593
rect 28629 22593 28641 22627
rect 28675 22624 28687 22627
rect 28902 22624 28908 22636
rect 28675 22596 28908 22624
rect 28675 22593 28687 22596
rect 28629 22587 28687 22593
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 31297 22627 31355 22633
rect 31297 22593 31309 22627
rect 31343 22593 31355 22627
rect 31297 22587 31355 22593
rect 27249 22559 27307 22565
rect 27249 22525 27261 22559
rect 27295 22556 27307 22559
rect 27338 22556 27344 22568
rect 27295 22528 27344 22556
rect 27295 22525 27307 22528
rect 27249 22519 27307 22525
rect 27338 22516 27344 22528
rect 27396 22556 27402 22568
rect 27614 22556 27620 22568
rect 27396 22528 27620 22556
rect 27396 22516 27402 22528
rect 27614 22516 27620 22528
rect 27672 22556 27678 22568
rect 28718 22556 28724 22568
rect 27672 22528 28580 22556
rect 28679 22528 28724 22556
rect 27672 22516 27678 22528
rect 26206 22460 27016 22488
rect 1486 22420 1492 22432
rect 1447 22392 1492 22420
rect 1486 22380 1492 22392
rect 1544 22380 1550 22432
rect 3418 22420 3424 22432
rect 3379 22392 3424 22420
rect 3418 22380 3424 22392
rect 3476 22380 3482 22432
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 22741 22423 22799 22429
rect 22741 22420 22753 22423
rect 22152 22392 22753 22420
rect 22152 22380 22158 22392
rect 22741 22389 22753 22392
rect 22787 22389 22799 22423
rect 24026 22420 24032 22432
rect 23987 22392 24032 22420
rect 22741 22383 22799 22389
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 24302 22380 24308 22432
rect 24360 22420 24366 22432
rect 25314 22420 25320 22432
rect 24360 22392 25320 22420
rect 24360 22380 24366 22392
rect 25314 22380 25320 22392
rect 25372 22420 25378 22432
rect 25685 22423 25743 22429
rect 25685 22420 25697 22423
rect 25372 22392 25697 22420
rect 25372 22380 25378 22392
rect 25685 22389 25697 22392
rect 25731 22420 25743 22423
rect 26206 22420 26234 22460
rect 27062 22448 27068 22500
rect 27120 22488 27126 22500
rect 28261 22491 28319 22497
rect 28261 22488 28273 22491
rect 27120 22460 28273 22488
rect 27120 22448 27126 22460
rect 28261 22457 28273 22460
rect 28307 22457 28319 22491
rect 28552 22488 28580 22528
rect 28718 22516 28724 22528
rect 28776 22516 28782 22568
rect 28813 22559 28871 22565
rect 28813 22525 28825 22559
rect 28859 22525 28871 22559
rect 31312 22556 31340 22587
rect 34514 22584 34520 22636
rect 34572 22624 34578 22636
rect 34977 22627 35035 22633
rect 34977 22624 34989 22627
rect 34572 22596 34989 22624
rect 34572 22584 34578 22596
rect 34977 22593 34989 22596
rect 35023 22593 35035 22627
rect 35802 22624 35808 22636
rect 35763 22596 35808 22624
rect 34977 22587 35035 22593
rect 35802 22584 35808 22596
rect 35860 22584 35866 22636
rect 37458 22633 37464 22636
rect 37456 22624 37464 22633
rect 37419 22596 37464 22624
rect 37456 22587 37464 22596
rect 37458 22584 37464 22587
rect 37516 22584 37522 22636
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22593 37611 22627
rect 37553 22587 37611 22593
rect 32125 22559 32183 22565
rect 32125 22556 32137 22559
rect 31312 22528 32137 22556
rect 28813 22519 28871 22525
rect 32125 22525 32137 22528
rect 32171 22525 32183 22559
rect 32125 22519 32183 22525
rect 28828 22488 28856 22519
rect 32490 22516 32496 22568
rect 32548 22556 32554 22568
rect 32585 22559 32643 22565
rect 32585 22556 32597 22559
rect 32548 22528 32597 22556
rect 32548 22516 32554 22528
rect 32585 22525 32597 22528
rect 32631 22556 32643 22559
rect 33689 22559 33747 22565
rect 33689 22556 33701 22559
rect 32631 22528 33701 22556
rect 32631 22525 32643 22528
rect 32585 22519 32643 22525
rect 33689 22525 33701 22528
rect 33735 22556 33747 22559
rect 34606 22556 34612 22568
rect 33735 22528 34612 22556
rect 33735 22525 33747 22528
rect 33689 22519 33747 22525
rect 34606 22516 34612 22528
rect 34664 22516 34670 22568
rect 34790 22556 34796 22568
rect 34751 22528 34796 22556
rect 34790 22516 34796 22528
rect 34848 22516 34854 22568
rect 37182 22516 37188 22568
rect 37240 22556 37246 22568
rect 37568 22556 37596 22587
rect 37734 22584 37740 22636
rect 37792 22633 37798 22636
rect 37792 22627 37831 22633
rect 37819 22593 37831 22627
rect 37792 22587 37831 22593
rect 37921 22627 37979 22633
rect 37921 22593 37933 22627
rect 37967 22624 37979 22627
rect 38102 22624 38108 22636
rect 37967 22596 38108 22624
rect 37967 22593 37979 22596
rect 37921 22587 37979 22593
rect 37792 22584 37798 22587
rect 38102 22584 38108 22596
rect 38160 22584 38166 22636
rect 38194 22556 38200 22568
rect 37240 22528 38200 22556
rect 37240 22516 37246 22528
rect 38194 22516 38200 22528
rect 38252 22516 38258 22568
rect 32214 22488 32220 22500
rect 28552 22460 28856 22488
rect 32175 22460 32220 22488
rect 28261 22451 28319 22457
rect 32214 22448 32220 22460
rect 32272 22448 32278 22500
rect 34054 22488 34060 22500
rect 34015 22460 34060 22488
rect 34054 22448 34060 22460
rect 34112 22448 34118 22500
rect 35066 22448 35072 22500
rect 35124 22488 35130 22500
rect 35345 22491 35403 22497
rect 35345 22488 35357 22491
rect 35124 22460 35357 22488
rect 35124 22448 35130 22460
rect 35345 22457 35357 22460
rect 35391 22457 35403 22491
rect 37277 22491 37335 22497
rect 37277 22488 37289 22491
rect 35345 22451 35403 22457
rect 35866 22460 37289 22488
rect 27798 22420 27804 22432
rect 25731 22392 26234 22420
rect 27759 22392 27804 22420
rect 25731 22389 25743 22392
rect 25685 22383 25743 22389
rect 27798 22380 27804 22392
rect 27856 22380 27862 22432
rect 31018 22380 31024 22432
rect 31076 22420 31082 22432
rect 35866 22420 35894 22460
rect 37277 22457 37289 22460
rect 37323 22457 37335 22491
rect 37277 22451 37335 22457
rect 31076 22392 35894 22420
rect 35989 22423 36047 22429
rect 31076 22380 31082 22392
rect 35989 22389 36001 22423
rect 36035 22420 36047 22423
rect 36078 22420 36084 22432
rect 36035 22392 36084 22420
rect 36035 22389 36047 22392
rect 35989 22383 36047 22389
rect 36078 22380 36084 22392
rect 36136 22380 36142 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 28902 22176 28908 22228
rect 28960 22216 28966 22228
rect 34057 22219 34115 22225
rect 34057 22216 34069 22219
rect 28960 22188 34069 22216
rect 28960 22176 28966 22188
rect 34057 22185 34069 22188
rect 34103 22216 34115 22219
rect 34514 22216 34520 22228
rect 34103 22188 34520 22216
rect 34103 22185 34115 22188
rect 34057 22179 34115 22185
rect 34514 22176 34520 22188
rect 34572 22176 34578 22228
rect 35161 22219 35219 22225
rect 35161 22185 35173 22219
rect 35207 22216 35219 22219
rect 35802 22216 35808 22228
rect 35207 22188 35808 22216
rect 35207 22185 35219 22188
rect 35161 22179 35219 22185
rect 35802 22176 35808 22188
rect 35860 22176 35866 22228
rect 35986 22176 35992 22228
rect 36044 22216 36050 22228
rect 37182 22216 37188 22228
rect 36044 22188 37188 22216
rect 36044 22176 36050 22188
rect 37182 22176 37188 22188
rect 37240 22176 37246 22228
rect 25869 22151 25927 22157
rect 25869 22117 25881 22151
rect 25915 22148 25927 22151
rect 26326 22148 26332 22160
rect 25915 22120 26332 22148
rect 25915 22117 25927 22120
rect 25869 22111 25927 22117
rect 26326 22108 26332 22120
rect 26384 22108 26390 22160
rect 27798 22108 27804 22160
rect 27856 22148 27862 22160
rect 28353 22151 28411 22157
rect 28353 22148 28365 22151
rect 27856 22120 28365 22148
rect 27856 22108 27862 22120
rect 28353 22117 28365 22120
rect 28399 22117 28411 22151
rect 28353 22111 28411 22117
rect 34698 22108 34704 22160
rect 34756 22148 34762 22160
rect 34977 22151 35035 22157
rect 34977 22148 34989 22151
rect 34756 22120 34989 22148
rect 34756 22108 34762 22120
rect 34977 22117 34989 22120
rect 35023 22117 35035 22151
rect 34977 22111 35035 22117
rect 2133 22083 2191 22089
rect 2133 22049 2145 22083
rect 2179 22080 2191 22083
rect 17218 22080 17224 22092
rect 2179 22052 17224 22080
rect 2179 22049 2191 22052
rect 2133 22043 2191 22049
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 22646 22040 22652 22092
rect 22704 22080 22710 22092
rect 23290 22080 23296 22092
rect 22704 22052 23296 22080
rect 22704 22040 22710 22052
rect 22554 22012 22560 22024
rect 22515 21984 22560 22012
rect 22554 21972 22560 21984
rect 22612 21972 22618 22024
rect 22848 22021 22876 22052
rect 23290 22040 23296 22052
rect 23348 22040 23354 22092
rect 25501 22083 25559 22089
rect 25501 22049 25513 22083
rect 25547 22080 25559 22083
rect 26142 22080 26148 22092
rect 25547 22052 26148 22080
rect 25547 22049 25559 22052
rect 25501 22043 25559 22049
rect 26142 22040 26148 22052
rect 26200 22040 26206 22092
rect 27430 22040 27436 22092
rect 27488 22080 27494 22092
rect 28074 22080 28080 22092
rect 27488 22052 28080 22080
rect 27488 22040 27494 22052
rect 28074 22040 28080 22052
rect 28132 22040 28138 22092
rect 28258 22080 28264 22092
rect 28219 22052 28264 22080
rect 28258 22040 28264 22052
rect 28316 22040 28322 22092
rect 28442 22040 28448 22092
rect 28500 22080 28506 22092
rect 28902 22080 28908 22092
rect 28500 22052 28908 22080
rect 28500 22040 28506 22052
rect 28902 22040 28908 22052
rect 28960 22040 28966 22092
rect 35342 22080 35348 22092
rect 32876 22052 35348 22080
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 24026 22012 24032 22024
rect 23063 21984 24032 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 24026 21972 24032 21984
rect 24084 21972 24090 22024
rect 24394 22012 24400 22024
rect 24355 21984 24400 22012
rect 24394 21972 24400 21984
rect 24452 21972 24458 22024
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 22012 24639 22015
rect 24946 22012 24952 22024
rect 24627 21984 24952 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 26234 21972 26240 22024
rect 26292 22012 26298 22024
rect 26421 22015 26479 22021
rect 26421 22012 26433 22015
rect 26292 21984 26433 22012
rect 26292 21972 26298 21984
rect 26421 21981 26433 21984
rect 26467 22012 26479 22015
rect 27522 22012 27528 22024
rect 26467 21984 27528 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 27522 21972 27528 21984
rect 27580 21972 27586 22024
rect 28626 22012 28632 22024
rect 27632 21984 28632 22012
rect 1854 21944 1860 21956
rect 1815 21916 1860 21944
rect 1854 21904 1860 21916
rect 1912 21944 1918 21956
rect 22738 21953 22744 21956
rect 2685 21947 2743 21953
rect 2685 21944 2697 21947
rect 1912 21916 2697 21944
rect 1912 21904 1918 21916
rect 2685 21913 2697 21916
rect 2731 21913 2743 21947
rect 2685 21907 2743 21913
rect 22715 21947 22744 21953
rect 22715 21913 22727 21947
rect 22715 21907 22744 21913
rect 22738 21904 22744 21907
rect 22796 21904 22802 21956
rect 22925 21947 22983 21953
rect 22925 21913 22937 21947
rect 22971 21944 22983 21947
rect 23661 21947 23719 21953
rect 23661 21944 23673 21947
rect 22971 21916 23673 21944
rect 22971 21913 22983 21916
rect 22925 21907 22983 21913
rect 23661 21913 23673 21916
rect 23707 21944 23719 21947
rect 23707 21916 26096 21944
rect 23707 21913 23719 21916
rect 23661 21907 23719 21913
rect 3418 21836 3424 21888
rect 3476 21876 3482 21888
rect 23201 21879 23259 21885
rect 23201 21876 23213 21879
rect 3476 21848 23213 21876
rect 3476 21836 3482 21848
rect 23201 21845 23213 21848
rect 23247 21845 23259 21879
rect 23201 21839 23259 21845
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 24765 21879 24823 21885
rect 24765 21876 24777 21879
rect 23808 21848 24777 21876
rect 23808 21836 23814 21848
rect 24765 21845 24777 21848
rect 24811 21845 24823 21879
rect 25958 21876 25964 21888
rect 25919 21848 25964 21876
rect 24765 21839 24823 21845
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 26068 21876 26096 21916
rect 26510 21904 26516 21956
rect 26568 21944 26574 21956
rect 26666 21947 26724 21953
rect 26666 21944 26678 21947
rect 26568 21916 26678 21944
rect 26568 21904 26574 21916
rect 26666 21913 26678 21916
rect 26712 21913 26724 21947
rect 26666 21907 26724 21913
rect 27632 21876 27660 21984
rect 28626 21972 28632 21984
rect 28684 21972 28690 22024
rect 31386 22012 31392 22024
rect 30944 21984 31392 22012
rect 28074 21904 28080 21956
rect 28132 21944 28138 21956
rect 28721 21947 28779 21953
rect 28721 21944 28733 21947
rect 28132 21916 28733 21944
rect 28132 21904 28138 21916
rect 28721 21913 28733 21916
rect 28767 21913 28779 21947
rect 28721 21907 28779 21913
rect 29822 21904 29828 21956
rect 29880 21944 29886 21956
rect 30837 21947 30895 21953
rect 30837 21944 30849 21947
rect 29880 21916 30849 21944
rect 29880 21904 29886 21916
rect 30837 21913 30849 21916
rect 30883 21913 30895 21947
rect 30837 21907 30895 21913
rect 30944 21888 30972 21984
rect 31386 21972 31392 21984
rect 31444 22012 31450 22024
rect 32876 22021 32904 22052
rect 35342 22040 35348 22052
rect 35400 22080 35406 22092
rect 35805 22083 35863 22089
rect 35805 22080 35817 22083
rect 35400 22052 35817 22080
rect 35400 22040 35406 22052
rect 35805 22049 35817 22052
rect 35851 22049 35863 22083
rect 35805 22043 35863 22049
rect 37642 22040 37648 22092
rect 37700 22080 37706 22092
rect 38010 22080 38016 22092
rect 37700 22052 38016 22080
rect 37700 22040 37706 22052
rect 38010 22040 38016 22052
rect 38068 22040 38074 22092
rect 32861 22015 32919 22021
rect 32861 22012 32873 22015
rect 31444 21984 32873 22012
rect 31444 21972 31450 21984
rect 32861 21981 32873 21984
rect 32907 21981 32919 22015
rect 33502 22012 33508 22024
rect 33463 21984 33508 22012
rect 32861 21975 32919 21981
rect 33502 21972 33508 21984
rect 33560 21972 33566 22024
rect 34606 21972 34612 22024
rect 34664 22012 34670 22024
rect 36078 22021 36084 22024
rect 34701 22015 34759 22021
rect 34701 22012 34713 22015
rect 34664 21984 34713 22012
rect 34664 21972 34670 21984
rect 34701 21981 34713 21984
rect 34747 21981 34759 22015
rect 34701 21975 34759 21981
rect 36072 21975 36084 22021
rect 36136 22012 36142 22024
rect 37829 22015 37887 22021
rect 36136 21984 36172 22012
rect 36078 21972 36084 21975
rect 36136 21972 36142 21984
rect 37829 21981 37841 22015
rect 37875 22012 37887 22015
rect 37918 22012 37924 22024
rect 37875 21984 37924 22012
rect 37875 21981 37887 21984
rect 37829 21975 37887 21981
rect 37918 21972 37924 21984
rect 37976 21972 37982 22024
rect 32616 21947 32674 21953
rect 32616 21913 32628 21947
rect 32662 21944 32674 21947
rect 32662 21916 33364 21944
rect 32662 21913 32674 21916
rect 32616 21907 32674 21913
rect 26068 21848 27660 21876
rect 27798 21836 27804 21888
rect 27856 21876 27862 21888
rect 28994 21876 29000 21888
rect 27856 21848 29000 21876
rect 27856 21836 27862 21848
rect 28994 21836 29000 21848
rect 29052 21836 29058 21888
rect 30926 21876 30932 21888
rect 30887 21848 30932 21876
rect 30926 21836 30932 21848
rect 30984 21836 30990 21888
rect 31481 21879 31539 21885
rect 31481 21845 31493 21879
rect 31527 21876 31539 21879
rect 32398 21876 32404 21888
rect 31527 21848 32404 21876
rect 31527 21845 31539 21848
rect 31481 21839 31539 21845
rect 32398 21836 32404 21848
rect 32456 21836 32462 21888
rect 33336 21885 33364 21916
rect 33321 21879 33379 21885
rect 33321 21845 33333 21879
rect 33367 21845 33379 21879
rect 38010 21876 38016 21888
rect 37971 21848 38016 21876
rect 33321 21839 33379 21845
rect 38010 21836 38016 21848
rect 38068 21836 38074 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 17218 21632 17224 21684
rect 17276 21672 17282 21684
rect 22646 21672 22652 21684
rect 17276 21644 22652 21672
rect 17276 21632 17282 21644
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 24118 21672 24124 21684
rect 22796 21644 24124 21672
rect 22796 21632 22802 21644
rect 24118 21632 24124 21644
rect 24176 21632 24182 21684
rect 26421 21675 26479 21681
rect 26421 21641 26433 21675
rect 26467 21672 26479 21675
rect 26510 21672 26516 21684
rect 26467 21644 26516 21672
rect 26467 21641 26479 21644
rect 26421 21635 26479 21641
rect 26510 21632 26516 21644
rect 26568 21632 26574 21684
rect 28258 21672 28264 21684
rect 26620 21644 28264 21672
rect 13814 21604 13820 21616
rect 13727 21576 13820 21604
rect 13814 21564 13820 21576
rect 13872 21604 13878 21616
rect 24302 21604 24308 21616
rect 13872 21576 24308 21604
rect 13872 21564 13878 21576
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21536 1458 21548
rect 2041 21539 2099 21545
rect 2041 21536 2053 21539
rect 1452 21508 2053 21536
rect 1452 21496 1458 21508
rect 2041 21505 2053 21508
rect 2087 21505 2099 21539
rect 14458 21536 14464 21548
rect 14419 21508 14464 21536
rect 2041 21499 2099 21505
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 14752 21545 14780 21576
rect 24302 21564 24308 21576
rect 24360 21564 24366 21616
rect 24394 21564 24400 21616
rect 24452 21604 24458 21616
rect 24673 21607 24731 21613
rect 24673 21604 24685 21607
rect 24452 21576 24685 21604
rect 24452 21564 24458 21576
rect 24673 21573 24685 21576
rect 24719 21573 24731 21607
rect 24673 21567 24731 21573
rect 14737 21539 14795 21545
rect 14737 21505 14749 21539
rect 14783 21505 14795 21539
rect 14737 21499 14795 21505
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 18121 21539 18179 21545
rect 18121 21536 18133 21539
rect 17460 21508 18133 21536
rect 17460 21496 17466 21508
rect 18121 21505 18133 21508
rect 18167 21505 18179 21539
rect 24486 21536 24492 21548
rect 24447 21508 24492 21536
rect 18121 21499 18179 21505
rect 24486 21496 24492 21508
rect 24544 21496 24550 21548
rect 25958 21496 25964 21548
rect 26016 21536 26022 21548
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 26016 21508 26249 21536
rect 26016 21496 26022 21508
rect 26237 21505 26249 21508
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 17865 21471 17923 21477
rect 17865 21468 17877 21471
rect 17328 21440 17877 21468
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 3050 21332 3056 21344
rect 1627 21304 3056 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 14274 21332 14280 21344
rect 14235 21304 14280 21332
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14550 21292 14556 21344
rect 14608 21332 14614 21344
rect 14645 21335 14703 21341
rect 14645 21332 14657 21335
rect 14608 21304 14657 21332
rect 14608 21292 14614 21304
rect 14645 21301 14657 21304
rect 14691 21301 14703 21335
rect 14645 21295 14703 21301
rect 16482 21292 16488 21344
rect 16540 21332 16546 21344
rect 17328 21341 17356 21440
rect 17865 21437 17877 21440
rect 17911 21437 17923 21471
rect 17865 21431 17923 21437
rect 23566 21428 23572 21480
rect 23624 21468 23630 21480
rect 26620 21468 26648 21644
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 29822 21672 29828 21684
rect 28368 21644 29828 21672
rect 27522 21564 27528 21616
rect 27580 21604 27586 21616
rect 28368 21613 28396 21644
rect 29822 21632 29828 21644
rect 29880 21632 29886 21684
rect 32125 21675 32183 21681
rect 32125 21641 32137 21675
rect 32171 21672 32183 21675
rect 32214 21672 32220 21684
rect 32171 21644 32220 21672
rect 32171 21641 32183 21644
rect 32125 21635 32183 21641
rect 32214 21632 32220 21644
rect 32272 21632 32278 21684
rect 32585 21675 32643 21681
rect 32585 21641 32597 21675
rect 32631 21672 32643 21675
rect 32766 21672 32772 21684
rect 32631 21644 32772 21672
rect 32631 21641 32643 21644
rect 32585 21635 32643 21641
rect 32766 21632 32772 21644
rect 32824 21632 32830 21684
rect 34054 21632 34060 21684
rect 34112 21672 34118 21684
rect 34609 21675 34667 21681
rect 34609 21672 34621 21675
rect 34112 21644 34621 21672
rect 34112 21632 34118 21644
rect 34609 21641 34621 21644
rect 34655 21641 34667 21675
rect 34609 21635 34667 21641
rect 37366 21632 37372 21684
rect 37424 21632 37430 21684
rect 28169 21607 28227 21613
rect 28169 21604 28181 21607
rect 27580 21576 28181 21604
rect 27580 21564 27586 21576
rect 28169 21573 28181 21576
rect 28215 21573 28227 21607
rect 28169 21567 28227 21573
rect 28353 21607 28411 21613
rect 28353 21573 28365 21607
rect 28399 21573 28411 21607
rect 35069 21607 35127 21613
rect 28353 21567 28411 21573
rect 29288 21576 31754 21604
rect 27338 21536 27344 21548
rect 27299 21508 27344 21536
rect 27338 21496 27344 21508
rect 27396 21536 27402 21548
rect 29288 21536 29316 21576
rect 27396 21508 29316 21536
rect 27396 21496 27402 21508
rect 29454 21496 29460 21548
rect 29512 21536 29518 21548
rect 29917 21539 29975 21545
rect 29917 21536 29929 21539
rect 29512 21508 29929 21536
rect 29512 21496 29518 21508
rect 29917 21505 29929 21508
rect 29963 21505 29975 21539
rect 31726 21536 31754 21576
rect 35069 21573 35081 21607
rect 35115 21604 35127 21607
rect 35894 21604 35900 21616
rect 35115 21576 35900 21604
rect 35115 21573 35127 21576
rect 35069 21567 35127 21573
rect 35894 21564 35900 21576
rect 35952 21604 35958 21616
rect 36357 21607 36415 21613
rect 36357 21604 36369 21607
rect 35952 21576 36369 21604
rect 35952 21564 35958 21576
rect 36357 21573 36369 21576
rect 36403 21573 36415 21607
rect 37384 21604 37412 21632
rect 37645 21607 37703 21613
rect 37645 21604 37657 21607
rect 36357 21567 36415 21573
rect 36464 21576 37657 21604
rect 36464 21548 36492 21576
rect 37645 21573 37657 21576
rect 37691 21573 37703 21607
rect 37645 21567 37703 21573
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 31726 21508 32505 21536
rect 29917 21499 29975 21505
rect 32493 21505 32505 21508
rect 32539 21536 32551 21539
rect 33321 21539 33379 21545
rect 33321 21536 33333 21539
rect 32539 21508 33333 21536
rect 32539 21505 32551 21508
rect 32493 21499 32551 21505
rect 33321 21505 33333 21508
rect 33367 21505 33379 21539
rect 33321 21499 33379 21505
rect 33962 21496 33968 21548
rect 34020 21536 34026 21548
rect 34057 21539 34115 21545
rect 34057 21536 34069 21539
rect 34020 21508 34069 21536
rect 34020 21496 34026 21508
rect 34057 21505 34069 21508
rect 34103 21536 34115 21539
rect 34977 21539 35035 21545
rect 34977 21536 34989 21539
rect 34103 21508 34989 21536
rect 34103 21505 34115 21508
rect 34057 21499 34115 21505
rect 34977 21505 34989 21508
rect 35023 21505 35035 21539
rect 34977 21499 35035 21505
rect 36260 21539 36318 21545
rect 36260 21505 36272 21539
rect 36306 21536 36318 21539
rect 36306 21508 36400 21536
rect 36306 21505 36318 21508
rect 36260 21499 36318 21505
rect 23624 21440 26648 21468
rect 23624 21428 23630 21440
rect 27154 21428 27160 21480
rect 27212 21468 27218 21480
rect 27433 21471 27491 21477
rect 27433 21468 27445 21471
rect 27212 21440 27445 21468
rect 27212 21428 27218 21440
rect 27433 21437 27445 21440
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 27525 21471 27583 21477
rect 27525 21437 27537 21471
rect 27571 21468 27583 21471
rect 27614 21468 27620 21480
rect 27571 21440 27620 21468
rect 27571 21437 27583 21440
rect 27525 21431 27583 21437
rect 22646 21360 22652 21412
rect 22704 21400 22710 21412
rect 24762 21400 24768 21412
rect 22704 21372 24768 21400
rect 22704 21360 22710 21372
rect 24762 21360 24768 21372
rect 24820 21360 24826 21412
rect 26326 21360 26332 21412
rect 26384 21400 26390 21412
rect 26973 21403 27031 21409
rect 26973 21400 26985 21403
rect 26384 21372 26985 21400
rect 26384 21360 26390 21372
rect 26973 21369 26985 21372
rect 27019 21369 27031 21403
rect 27448 21400 27476 21431
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 31113 21471 31171 21477
rect 31113 21437 31125 21471
rect 31159 21468 31171 21471
rect 32306 21468 32312 21480
rect 31159 21440 32312 21468
rect 31159 21437 31171 21440
rect 31113 21431 31171 21437
rect 32306 21428 32312 21440
rect 32364 21428 32370 21480
rect 32769 21471 32827 21477
rect 32769 21437 32781 21471
rect 32815 21468 32827 21471
rect 32950 21468 32956 21480
rect 32815 21440 32956 21468
rect 32815 21437 32827 21440
rect 32769 21431 32827 21437
rect 32950 21428 32956 21440
rect 33008 21468 33014 21480
rect 34790 21468 34796 21480
rect 33008 21440 34796 21468
rect 33008 21428 33014 21440
rect 34790 21428 34796 21440
rect 34848 21468 34854 21480
rect 35161 21471 35219 21477
rect 35161 21468 35173 21471
rect 34848 21440 35173 21468
rect 34848 21428 34854 21440
rect 35161 21437 35173 21440
rect 35207 21468 35219 21471
rect 35342 21468 35348 21480
rect 35207 21440 35348 21468
rect 35207 21437 35219 21440
rect 35161 21431 35219 21437
rect 35342 21428 35348 21440
rect 35400 21428 35406 21480
rect 27798 21400 27804 21412
rect 27448 21372 27804 21400
rect 26973 21363 27031 21369
rect 27798 21360 27804 21372
rect 27856 21360 27862 21412
rect 31481 21403 31539 21409
rect 31481 21369 31493 21403
rect 31527 21400 31539 21403
rect 31938 21400 31944 21412
rect 31527 21372 31944 21400
rect 31527 21369 31539 21372
rect 31481 21363 31539 21369
rect 31938 21360 31944 21372
rect 31996 21360 32002 21412
rect 36372 21400 36400 21508
rect 36446 21496 36452 21548
rect 36504 21536 36510 21548
rect 36630 21536 36636 21548
rect 36504 21508 36549 21536
rect 36591 21508 36636 21536
rect 36504 21496 36510 21508
rect 36630 21496 36636 21508
rect 36688 21496 36694 21548
rect 36725 21539 36783 21545
rect 36725 21505 36737 21539
rect 36771 21536 36783 21539
rect 36906 21536 36912 21548
rect 36771 21508 36912 21536
rect 36771 21505 36783 21508
rect 36725 21499 36783 21505
rect 36906 21496 36912 21508
rect 36964 21496 36970 21548
rect 36998 21496 37004 21548
rect 37056 21536 37062 21548
rect 37458 21545 37464 21548
rect 37415 21539 37464 21545
rect 37415 21536 37427 21539
rect 37056 21508 37427 21536
rect 37056 21496 37062 21508
rect 37415 21505 37427 21508
rect 37461 21505 37464 21539
rect 37415 21499 37464 21505
rect 37458 21496 37464 21499
rect 37516 21496 37522 21548
rect 37550 21496 37556 21548
rect 37608 21536 37614 21548
rect 37826 21536 37832 21548
rect 37608 21508 37653 21536
rect 37787 21508 37832 21536
rect 37608 21496 37614 21508
rect 37826 21496 37832 21508
rect 37884 21496 37890 21548
rect 37918 21496 37924 21548
rect 37976 21536 37982 21548
rect 38102 21536 38108 21548
rect 37976 21508 38108 21536
rect 37976 21496 37982 21508
rect 38102 21496 38108 21508
rect 38160 21496 38166 21548
rect 36998 21400 37004 21412
rect 36372 21372 37004 21400
rect 36998 21360 37004 21372
rect 37056 21360 37062 21412
rect 17313 21335 17371 21341
rect 17313 21332 17325 21335
rect 16540 21304 17325 21332
rect 16540 21292 16546 21304
rect 17313 21301 17325 21304
rect 17359 21301 17371 21335
rect 17313 21295 17371 21301
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 19245 21335 19303 21341
rect 19245 21332 19257 21335
rect 18840 21304 19257 21332
rect 18840 21292 18846 21304
rect 19245 21301 19257 21304
rect 19291 21301 19303 21335
rect 24302 21332 24308 21344
rect 24263 21304 24308 21332
rect 19245 21295 19303 21301
rect 24302 21292 24308 21304
rect 24360 21292 24366 21344
rect 24486 21292 24492 21344
rect 24544 21332 24550 21344
rect 25225 21335 25283 21341
rect 25225 21332 25237 21335
rect 24544 21304 25237 21332
rect 24544 21292 24550 21304
rect 25225 21301 25237 21304
rect 25271 21332 25283 21335
rect 28718 21332 28724 21344
rect 25271 21304 28724 21332
rect 25271 21301 25283 21304
rect 25225 21295 25283 21301
rect 28718 21292 28724 21304
rect 28776 21292 28782 21344
rect 31573 21335 31631 21341
rect 31573 21301 31585 21335
rect 31619 21332 31631 21335
rect 33502 21332 33508 21344
rect 31619 21304 33508 21332
rect 31619 21301 31631 21304
rect 31573 21295 31631 21301
rect 33502 21292 33508 21304
rect 33560 21292 33566 21344
rect 36078 21332 36084 21344
rect 36039 21304 36084 21332
rect 36078 21292 36084 21304
rect 36136 21292 36142 21344
rect 37277 21335 37335 21341
rect 37277 21301 37289 21335
rect 37323 21332 37335 21335
rect 37366 21332 37372 21344
rect 37323 21304 37372 21332
rect 37323 21301 37335 21304
rect 37277 21295 37335 21301
rect 37366 21292 37372 21304
rect 37424 21292 37430 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 13814 21128 13820 21140
rect 2280 21100 13820 21128
rect 2280 21088 2286 21100
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 23566 21128 23572 21140
rect 17972 21100 23572 21128
rect 14550 21020 14556 21072
rect 14608 21060 14614 21072
rect 16666 21060 16672 21072
rect 14608 21032 16672 21060
rect 14608 21020 14614 21032
rect 16666 21020 16672 21032
rect 16724 21060 16730 21072
rect 17865 21063 17923 21069
rect 17865 21060 17877 21063
rect 16724 21032 17877 21060
rect 16724 21020 16730 21032
rect 17865 21029 17877 21032
rect 17911 21029 17923 21063
rect 17865 21023 17923 21029
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 15010 20992 15016 21004
rect 2823 20964 2857 20992
rect 14660 20964 15016 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 2792 20924 2820 20955
rect 14660 20933 14688 20964
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 17972 20992 18000 21100
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 31018 21128 31024 21140
rect 23716 21100 31024 21128
rect 23716 21088 23722 21100
rect 31018 21088 31024 21100
rect 31076 21088 31082 21140
rect 31938 21128 31944 21140
rect 31899 21100 31944 21128
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 34146 21128 34152 21140
rect 34107 21100 34152 21128
rect 34146 21088 34152 21100
rect 34204 21088 34210 21140
rect 34716 21100 36860 21128
rect 21358 21020 21364 21072
rect 21416 21060 21422 21072
rect 26789 21063 26847 21069
rect 26789 21060 26801 21063
rect 21416 21032 26801 21060
rect 21416 21020 21422 21032
rect 26789 21029 26801 21032
rect 26835 21060 26847 21063
rect 27338 21060 27344 21072
rect 26835 21032 27344 21060
rect 26835 21029 26847 21032
rect 26789 21023 26847 21029
rect 27338 21020 27344 21032
rect 27396 21020 27402 21072
rect 34716 21060 34744 21100
rect 36832 21069 36860 21100
rect 36906 21088 36912 21140
rect 36964 21128 36970 21140
rect 37826 21128 37832 21140
rect 36964 21100 37832 21128
rect 36964 21088 36970 21100
rect 37826 21088 37832 21100
rect 37884 21088 37890 21140
rect 31726 21032 34744 21060
rect 36817 21063 36875 21069
rect 17788 20964 18000 20992
rect 14645 20927 14703 20933
rect 1719 20896 12434 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 12406 20856 12434 20896
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14918 20924 14924 20936
rect 14879 20896 14924 20924
rect 14645 20887 14703 20893
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 15105 20927 15163 20933
rect 15105 20893 15117 20927
rect 15151 20924 15163 20927
rect 15654 20924 15660 20936
rect 15151 20896 15660 20924
rect 15151 20893 15163 20896
rect 15105 20887 15163 20893
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 17126 20884 17132 20936
rect 17184 20924 17190 20936
rect 17788 20933 17816 20964
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 31726 20992 31754 21032
rect 36817 21029 36829 21063
rect 36863 21029 36875 21063
rect 36817 21023 36875 21029
rect 20128 20964 31754 20992
rect 32585 20995 32643 21001
rect 20128 20952 20134 20964
rect 32585 20961 32597 20995
rect 32631 20992 32643 20995
rect 32950 20992 32956 21004
rect 32631 20964 32956 20992
rect 32631 20961 32643 20964
rect 32585 20955 32643 20961
rect 32950 20952 32956 20964
rect 33008 20952 33014 21004
rect 35342 20992 35348 21004
rect 34072 20964 35204 20992
rect 35303 20964 35348 20992
rect 17773 20927 17831 20933
rect 17773 20924 17785 20927
rect 17184 20896 17785 20924
rect 17184 20884 17190 20896
rect 17773 20893 17785 20896
rect 17819 20893 17831 20927
rect 18046 20924 18052 20936
rect 18007 20896 18052 20924
rect 17773 20887 17831 20893
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 24394 20884 24400 20936
rect 24452 20924 24458 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24452 20896 24777 20924
rect 24452 20884 24458 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 32398 20924 32404 20936
rect 32311 20896 32404 20924
rect 24765 20887 24823 20893
rect 32398 20884 32404 20896
rect 32456 20924 32462 20936
rect 34072 20924 34100 20964
rect 32456 20896 34100 20924
rect 32456 20884 32462 20896
rect 34146 20884 34152 20936
rect 34204 20924 34210 20936
rect 35069 20927 35127 20933
rect 35069 20924 35081 20927
rect 34204 20896 35081 20924
rect 34204 20884 34210 20896
rect 35069 20893 35081 20896
rect 35115 20893 35127 20927
rect 35176 20924 35204 20964
rect 35342 20952 35348 20964
rect 35400 20952 35406 21004
rect 37642 20992 37648 21004
rect 35452 20964 37648 20992
rect 35452 20924 35480 20964
rect 35176 20896 35480 20924
rect 35989 20927 36047 20933
rect 35069 20887 35127 20893
rect 35989 20893 36001 20927
rect 36035 20924 36047 20927
rect 36814 20924 36820 20936
rect 36035 20896 36820 20924
rect 36035 20893 36047 20896
rect 35989 20887 36047 20893
rect 36814 20884 36820 20896
rect 36872 20884 36878 20936
rect 36998 20933 37004 20936
rect 36996 20924 37004 20933
rect 36959 20896 37004 20924
rect 36996 20887 37004 20896
rect 36998 20884 37004 20887
rect 37056 20884 37062 20936
rect 37093 20927 37151 20933
rect 37093 20893 37105 20927
rect 37139 20924 37151 20927
rect 37200 20924 37228 20964
rect 37642 20952 37648 20964
rect 37700 20952 37706 21004
rect 37139 20896 37228 20924
rect 37368 20927 37426 20933
rect 37139 20893 37151 20896
rect 37093 20887 37151 20893
rect 37368 20893 37380 20927
rect 37414 20893 37426 20927
rect 37368 20887 37426 20893
rect 37461 20927 37519 20933
rect 37461 20893 37473 20927
rect 37507 20924 37519 20927
rect 37826 20924 37832 20936
rect 37507 20896 37832 20924
rect 37507 20893 37519 20896
rect 37461 20887 37519 20893
rect 22922 20856 22928 20868
rect 12406 20828 22928 20856
rect 22922 20816 22928 20828
rect 22980 20816 22986 20868
rect 24581 20859 24639 20865
rect 24581 20825 24593 20859
rect 24627 20856 24639 20859
rect 27154 20856 27160 20868
rect 24627 20828 27160 20856
rect 24627 20825 24639 20828
rect 24581 20819 24639 20825
rect 27154 20816 27160 20828
rect 27212 20816 27218 20868
rect 32309 20859 32367 20865
rect 32309 20856 32321 20859
rect 31726 20828 32321 20856
rect 1486 20788 1492 20800
rect 1447 20760 1492 20788
rect 1486 20748 1492 20760
rect 1544 20748 1550 20800
rect 1854 20748 1860 20800
rect 1912 20788 1918 20800
rect 2133 20791 2191 20797
rect 2133 20788 2145 20791
rect 1912 20760 2145 20788
rect 1912 20748 1918 20760
rect 2133 20757 2145 20760
rect 2179 20757 2191 20791
rect 2133 20751 2191 20757
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 14461 20791 14519 20797
rect 14461 20788 14473 20791
rect 14424 20760 14473 20788
rect 14424 20748 14430 20760
rect 14461 20757 14473 20760
rect 14507 20757 14519 20791
rect 15654 20788 15660 20800
rect 15615 20760 15660 20788
rect 14461 20751 14519 20757
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17221 20791 17279 20797
rect 17221 20788 17233 20791
rect 17184 20760 17233 20788
rect 17184 20748 17190 20760
rect 17221 20757 17233 20760
rect 17267 20757 17279 20791
rect 18230 20788 18236 20800
rect 18191 20760 18236 20788
rect 17221 20751 17279 20757
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 24397 20791 24455 20797
rect 24397 20788 24409 20791
rect 23624 20760 24409 20788
rect 23624 20748 23630 20760
rect 24397 20757 24409 20760
rect 24443 20757 24455 20791
rect 24397 20751 24455 20757
rect 24670 20748 24676 20800
rect 24728 20788 24734 20800
rect 25130 20788 25136 20800
rect 24728 20760 25136 20788
rect 24728 20748 24734 20760
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 31386 20788 31392 20800
rect 31347 20760 31392 20788
rect 31386 20748 31392 20760
rect 31444 20788 31450 20800
rect 31726 20788 31754 20828
rect 32309 20825 32321 20828
rect 32355 20825 32367 20859
rect 32309 20819 32367 20825
rect 37185 20859 37243 20865
rect 37185 20825 37197 20859
rect 37231 20825 37243 20859
rect 37384 20856 37412 20887
rect 37826 20884 37832 20896
rect 37884 20884 37890 20936
rect 38102 20924 38108 20936
rect 38063 20896 38108 20924
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 37384 20828 37964 20856
rect 37185 20819 37243 20825
rect 34698 20788 34704 20800
rect 31444 20760 31754 20788
rect 34659 20760 34704 20788
rect 31444 20748 31450 20760
rect 34698 20748 34704 20760
rect 34756 20748 34762 20800
rect 35161 20791 35219 20797
rect 35161 20757 35173 20791
rect 35207 20788 35219 20791
rect 35986 20788 35992 20800
rect 35207 20760 35992 20788
rect 35207 20757 35219 20760
rect 35161 20751 35219 20757
rect 35986 20748 35992 20760
rect 36044 20748 36050 20800
rect 36170 20788 36176 20800
rect 36131 20760 36176 20788
rect 36170 20748 36176 20760
rect 36228 20748 36234 20800
rect 36446 20748 36452 20800
rect 36504 20788 36510 20800
rect 37200 20788 37228 20819
rect 37642 20788 37648 20800
rect 36504 20760 37648 20788
rect 36504 20748 36510 20760
rect 37642 20748 37648 20760
rect 37700 20748 37706 20800
rect 37936 20797 37964 20828
rect 37921 20791 37979 20797
rect 37921 20757 37933 20791
rect 37967 20757 37979 20791
rect 37921 20751 37979 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 13538 20584 13544 20596
rect 13451 20556 13544 20584
rect 13538 20544 13544 20556
rect 13596 20584 13602 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 13596 20556 15393 20584
rect 13596 20544 13602 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 17402 20584 17408 20596
rect 17363 20556 17408 20584
rect 15381 20547 15439 20553
rect 14274 20525 14280 20528
rect 14268 20516 14280 20525
rect 14235 20488 14280 20516
rect 14268 20479 14280 20488
rect 14274 20476 14280 20479
rect 14332 20476 14338 20528
rect 15396 20516 15424 20547
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 18046 20544 18052 20596
rect 18104 20584 18110 20596
rect 19797 20587 19855 20593
rect 19797 20584 19809 20587
rect 18104 20556 19809 20584
rect 18104 20544 18110 20556
rect 19797 20553 19809 20556
rect 19843 20553 19855 20587
rect 23474 20584 23480 20596
rect 23435 20556 23480 20584
rect 19797 20547 19855 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 23569 20587 23627 20593
rect 23569 20553 23581 20587
rect 23615 20584 23627 20587
rect 23658 20584 23664 20596
rect 23615 20556 23664 20584
rect 23615 20553 23627 20556
rect 23569 20547 23627 20553
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 25222 20584 25228 20596
rect 25183 20556 25228 20584
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 27157 20587 27215 20593
rect 27157 20553 27169 20587
rect 27203 20584 27215 20587
rect 27430 20584 27436 20596
rect 27203 20556 27436 20584
rect 27203 20553 27215 20556
rect 27157 20547 27215 20553
rect 27430 20544 27436 20556
rect 27488 20544 27494 20596
rect 36722 20584 36728 20596
rect 36683 20556 36728 20584
rect 36722 20544 36728 20556
rect 36780 20544 36786 20596
rect 37366 20544 37372 20596
rect 37424 20544 37430 20596
rect 18132 20519 18190 20525
rect 15396 20488 17356 20516
rect 1854 20448 1860 20460
rect 1815 20420 1860 20448
rect 1854 20408 1860 20420
rect 1912 20408 1918 20460
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20448 2743 20451
rect 2774 20448 2780 20460
rect 2731 20420 2780 20448
rect 2731 20417 2743 20420
rect 2685 20411 2743 20417
rect 2774 20408 2780 20420
rect 2832 20448 2838 20460
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 2832 20420 3341 20448
rect 2832 20408 2838 20420
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 17218 20448 17224 20460
rect 3329 20411 3387 20417
rect 12406 20420 16160 20448
rect 17179 20420 17224 20448
rect 2133 20315 2191 20321
rect 2133 20281 2145 20315
rect 2179 20312 2191 20315
rect 12406 20312 12434 20420
rect 13906 20340 13912 20392
rect 13964 20380 13970 20392
rect 16132 20389 16160 20420
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 17328 20448 17356 20488
rect 18132 20485 18144 20519
rect 18178 20516 18190 20519
rect 18230 20516 18236 20528
rect 18178 20488 18236 20516
rect 18178 20485 18190 20488
rect 18132 20479 18190 20485
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 20530 20516 20536 20528
rect 18340 20488 20536 20516
rect 18340 20448 18368 20488
rect 20530 20476 20536 20488
rect 20588 20476 20594 20528
rect 22922 20516 22928 20528
rect 22883 20488 22928 20516
rect 22922 20476 22928 20488
rect 22980 20476 22986 20528
rect 24394 20476 24400 20528
rect 24452 20516 24458 20528
rect 24673 20519 24731 20525
rect 24673 20516 24685 20519
rect 24452 20488 24685 20516
rect 24452 20476 24458 20488
rect 24673 20485 24685 20488
rect 24719 20485 24731 20519
rect 24673 20479 24731 20485
rect 17328 20420 18368 20448
rect 18598 20408 18604 20460
rect 18656 20448 18662 20460
rect 19981 20451 20039 20457
rect 19981 20448 19993 20451
rect 18656 20420 19993 20448
rect 18656 20408 18662 20420
rect 19981 20417 19993 20420
rect 20027 20417 20039 20451
rect 20254 20448 20260 20460
rect 20215 20420 20260 20448
rect 19981 20411 20039 20417
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 20441 20451 20499 20457
rect 20441 20417 20453 20451
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 14001 20383 14059 20389
rect 14001 20380 14013 20383
rect 13964 20352 14013 20380
rect 13964 20340 13970 20352
rect 14001 20349 14013 20352
rect 14047 20349 14059 20383
rect 14001 20343 14059 20349
rect 16117 20383 16175 20389
rect 16117 20349 16129 20383
rect 16163 20380 16175 20383
rect 16942 20380 16948 20392
rect 16163 20352 16948 20380
rect 16163 20349 16175 20352
rect 16117 20343 16175 20349
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 17865 20383 17923 20389
rect 17865 20349 17877 20383
rect 17911 20349 17923 20383
rect 20456 20380 20484 20411
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 22244 20420 23121 20448
rect 22244 20408 22250 20420
rect 23109 20417 23121 20420
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20448 23719 20451
rect 23750 20448 23756 20460
rect 23707 20420 23756 20448
rect 23707 20417 23719 20420
rect 23661 20411 23719 20417
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20448 24547 20451
rect 25240 20448 25268 20544
rect 37384 20516 37412 20544
rect 24535 20420 25268 20448
rect 25700 20488 37412 20516
rect 37553 20519 37611 20525
rect 24535 20417 24547 20420
rect 24489 20411 24547 20417
rect 23382 20389 23388 20392
rect 17865 20343 17923 20349
rect 19996 20352 20484 20380
rect 23368 20383 23388 20389
rect 2179 20284 12434 20312
rect 2179 20281 2191 20284
rect 2133 20275 2191 20281
rect 16482 20272 16488 20324
rect 16540 20312 16546 20324
rect 17880 20312 17908 20343
rect 16540 20284 17908 20312
rect 16540 20272 16546 20284
rect 19996 20256 20024 20352
rect 23368 20349 23380 20383
rect 23368 20343 23388 20349
rect 23382 20340 23388 20343
rect 23440 20340 23446 20392
rect 22646 20272 22652 20324
rect 22704 20312 22710 20324
rect 25700 20312 25728 20488
rect 37553 20485 37565 20519
rect 37599 20516 37611 20519
rect 38378 20516 38384 20528
rect 37599 20488 38384 20516
rect 37599 20485 37611 20488
rect 37553 20479 37611 20485
rect 38378 20476 38384 20488
rect 38436 20476 38442 20528
rect 26973 20451 27031 20457
rect 26973 20417 26985 20451
rect 27019 20448 27031 20451
rect 27706 20448 27712 20460
rect 27019 20420 27712 20448
rect 27019 20417 27031 20420
rect 26973 20411 27031 20417
rect 27706 20408 27712 20420
rect 27764 20408 27770 20460
rect 29730 20408 29736 20460
rect 29788 20448 29794 20460
rect 30662 20451 30720 20457
rect 30662 20448 30674 20451
rect 29788 20420 30674 20448
rect 29788 20408 29794 20420
rect 30662 20417 30674 20420
rect 30708 20417 30720 20451
rect 30662 20411 30720 20417
rect 32306 20408 32312 20460
rect 32364 20448 32370 20460
rect 32769 20451 32827 20457
rect 32769 20448 32781 20451
rect 32364 20420 32781 20448
rect 32364 20408 32370 20420
rect 32769 20417 32781 20420
rect 32815 20417 32827 20451
rect 32769 20411 32827 20417
rect 37366 20408 37372 20460
rect 37424 20457 37430 20460
rect 37424 20451 37473 20457
rect 37424 20417 37427 20451
rect 37461 20417 37473 20451
rect 37642 20448 37648 20460
rect 37603 20420 37648 20448
rect 37424 20411 37473 20417
rect 37424 20408 37430 20411
rect 37642 20408 37648 20420
rect 37700 20408 37706 20460
rect 37734 20408 37740 20460
rect 37792 20457 37798 20460
rect 37792 20451 37831 20457
rect 37819 20417 37831 20451
rect 37792 20411 37831 20417
rect 37792 20408 37798 20411
rect 37918 20408 37924 20460
rect 37976 20448 37982 20460
rect 37976 20420 38021 20448
rect 37976 20408 37982 20420
rect 30926 20380 30932 20392
rect 30887 20352 30932 20380
rect 30926 20340 30932 20352
rect 30984 20340 30990 20392
rect 33042 20380 33048 20392
rect 33003 20352 33048 20380
rect 33042 20340 33048 20352
rect 33100 20340 33106 20392
rect 22704 20284 25728 20312
rect 22704 20272 22710 20284
rect 27522 20272 27528 20324
rect 27580 20312 27586 20324
rect 29549 20315 29607 20321
rect 29549 20312 29561 20315
rect 27580 20284 29561 20312
rect 27580 20272 27586 20284
rect 29549 20281 29561 20284
rect 29595 20281 29607 20315
rect 38010 20312 38016 20324
rect 29549 20275 29607 20281
rect 31726 20284 38016 20312
rect 2866 20244 2872 20256
rect 2827 20216 2872 20244
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 16666 20204 16672 20256
rect 16724 20244 16730 20256
rect 17037 20247 17095 20253
rect 17037 20244 17049 20247
rect 16724 20216 17049 20244
rect 16724 20204 16730 20216
rect 17037 20213 17049 20216
rect 17083 20213 17095 20247
rect 17037 20207 17095 20213
rect 19245 20247 19303 20253
rect 19245 20213 19257 20247
rect 19291 20244 19303 20247
rect 19978 20244 19984 20256
rect 19291 20216 19984 20244
rect 19291 20213 19303 20216
rect 19245 20207 19303 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 24305 20247 24363 20253
rect 24305 20244 24317 20247
rect 23808 20216 24317 20244
rect 23808 20204 23814 20216
rect 24305 20213 24317 20216
rect 24351 20213 24363 20247
rect 27706 20244 27712 20256
rect 27667 20216 27712 20244
rect 24305 20207 24363 20213
rect 27706 20204 27712 20216
rect 27764 20204 27770 20256
rect 29564 20244 29592 20275
rect 31726 20244 31754 20284
rect 38010 20272 38016 20284
rect 38068 20272 38074 20324
rect 37274 20244 37280 20256
rect 29564 20216 31754 20244
rect 37235 20216 37280 20244
rect 37274 20204 37280 20216
rect 37332 20204 37338 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 12897 20043 12955 20049
rect 12897 20009 12909 20043
rect 12943 20040 12955 20043
rect 14458 20040 14464 20052
rect 12943 20012 14464 20040
rect 12943 20009 12955 20012
rect 12897 20003 12955 20009
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 14918 20000 14924 20052
rect 14976 20040 14982 20052
rect 16666 20040 16672 20052
rect 14976 20012 15884 20040
rect 16627 20012 16672 20040
rect 14976 20000 14982 20012
rect 14936 19972 14964 20000
rect 13372 19944 14964 19972
rect 15856 19972 15884 20012
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 18049 20043 18107 20049
rect 18049 20040 18061 20043
rect 17276 20012 18061 20040
rect 17276 20000 17282 20012
rect 18049 20009 18061 20012
rect 18095 20009 18107 20043
rect 18049 20003 18107 20009
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 23017 20043 23075 20049
rect 23017 20040 23029 20043
rect 19484 20012 23029 20040
rect 19484 20000 19490 20012
rect 23017 20009 23029 20012
rect 23063 20009 23075 20043
rect 23017 20003 23075 20009
rect 24394 20000 24400 20052
rect 24452 20040 24458 20052
rect 24581 20043 24639 20049
rect 24581 20040 24593 20043
rect 24452 20012 24593 20040
rect 24452 20000 24458 20012
rect 24581 20009 24593 20012
rect 24627 20009 24639 20043
rect 24581 20003 24639 20009
rect 24670 20000 24676 20052
rect 24728 20040 24734 20052
rect 29730 20040 29736 20052
rect 24728 20012 28994 20040
rect 29691 20012 29736 20040
rect 24728 20000 24734 20012
rect 22646 19972 22652 19984
rect 15856 19944 18552 19972
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1719 19808 3924 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 1854 19728 1860 19780
rect 1912 19768 1918 19780
rect 2685 19771 2743 19777
rect 2685 19768 2697 19771
rect 1912 19740 2697 19768
rect 1912 19728 1918 19740
rect 2685 19737 2697 19740
rect 2731 19737 2743 19771
rect 2685 19731 2743 19737
rect 3896 19712 3924 19808
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 13372 19845 13400 19944
rect 18524 19904 18552 19944
rect 22480 19944 22652 19972
rect 20254 19904 20260 19916
rect 18524 19876 20260 19904
rect 13081 19839 13139 19845
rect 13081 19836 13093 19839
rect 10376 19808 13093 19836
rect 10376 19796 10382 19808
rect 13081 19805 13093 19808
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13446 19836 13452 19848
rect 13403 19808 13452 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13096 19768 13124 19799
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 15841 19839 15899 19845
rect 13596 19808 13641 19836
rect 13596 19796 13602 19808
rect 15841 19805 15853 19839
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 15194 19768 15200 19780
rect 13096 19740 15200 19768
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 15596 19771 15654 19777
rect 15596 19737 15608 19771
rect 15642 19768 15654 19771
rect 15856 19768 15884 19799
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 15988 19808 16497 19836
rect 15988 19796 15994 19808
rect 16485 19805 16497 19808
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 16666 19796 16672 19848
rect 16724 19836 16730 19848
rect 18524 19845 18552 19876
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 22480 19913 22508 19944
rect 22646 19932 22652 19944
rect 22704 19932 22710 19984
rect 22922 19932 22928 19984
rect 22980 19972 22986 19984
rect 27525 19975 27583 19981
rect 27525 19972 27537 19975
rect 22980 19944 27537 19972
rect 22980 19932 22986 19944
rect 27525 19941 27537 19944
rect 27571 19972 27583 19975
rect 28966 19972 28994 20012
rect 29730 20000 29736 20012
rect 29788 20000 29794 20052
rect 32950 20040 32956 20052
rect 32911 20012 32956 20040
rect 32950 20000 32956 20012
rect 33008 20000 33014 20052
rect 37274 19972 37280 19984
rect 27571 19944 28488 19972
rect 28966 19944 37280 19972
rect 27571 19941 27583 19944
rect 27525 19935 27583 19941
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19873 22523 19907
rect 22465 19867 22523 19873
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19904 22615 19907
rect 23566 19904 23572 19916
rect 22603 19876 23572 19904
rect 22603 19873 22615 19876
rect 22557 19867 22615 19873
rect 23566 19864 23572 19876
rect 23624 19864 23630 19916
rect 23750 19904 23756 19916
rect 23711 19876 23756 19904
rect 23750 19864 23756 19876
rect 23808 19864 23814 19916
rect 27614 19864 27620 19916
rect 27672 19904 27678 19916
rect 28169 19907 28227 19913
rect 28169 19904 28181 19907
rect 27672 19876 28181 19904
rect 27672 19864 27678 19876
rect 28169 19873 28181 19876
rect 28215 19873 28227 19907
rect 28169 19867 28227 19873
rect 28460 19904 28488 19944
rect 37274 19932 37280 19944
rect 37332 19932 37338 19984
rect 38010 19972 38016 19984
rect 37971 19944 38016 19972
rect 38010 19932 38016 19944
rect 38068 19932 38074 19984
rect 28810 19904 28816 19916
rect 28460 19876 28816 19904
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16724 19808 16773 19836
rect 16724 19796 16730 19808
rect 16761 19805 16773 19808
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19805 18567 19839
rect 18690 19836 18696 19848
rect 18651 19808 18696 19836
rect 18509 19799 18567 19805
rect 18248 19768 18276 19799
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 22261 19839 22319 19845
rect 22261 19805 22273 19839
rect 22307 19836 22319 19839
rect 22738 19836 22744 19848
rect 22307 19808 22744 19836
rect 22307 19805 22319 19808
rect 22261 19799 22319 19805
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23457 19839 23515 19845
rect 23457 19805 23469 19839
rect 23503 19836 23515 19839
rect 24210 19836 24216 19848
rect 23503 19808 24216 19836
rect 23503 19805 23515 19808
rect 23457 19799 23515 19805
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19836 24455 19839
rect 24854 19836 24860 19848
rect 24443 19808 24860 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 28460 19845 28488 19876
rect 28810 19864 28816 19876
rect 28868 19864 28874 19916
rect 28948 19864 28954 19916
rect 29006 19904 29012 19916
rect 31386 19904 31392 19916
rect 29006 19876 31392 19904
rect 29006 19864 29012 19876
rect 31386 19864 31392 19876
rect 31444 19864 31450 19916
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 27580 19808 28365 19836
rect 27580 19796 27586 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19805 28503 19839
rect 28920 19832 29040 19836
rect 28445 19799 28503 19805
rect 28828 19808 29040 19832
rect 28828 19804 28948 19808
rect 18598 19768 18604 19780
rect 15642 19740 15792 19768
rect 15856 19740 16528 19768
rect 18248 19740 18604 19768
rect 15642 19737 15654 19740
rect 15596 19731 15654 19737
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 2133 19703 2191 19709
rect 2133 19700 2145 19703
rect 2004 19672 2145 19700
rect 2004 19660 2010 19672
rect 2133 19669 2145 19672
rect 2179 19669 2191 19703
rect 3878 19700 3884 19712
rect 3839 19672 3884 19700
rect 2133 19663 2191 19669
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 14458 19700 14464 19712
rect 14419 19672 14464 19700
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 15764 19700 15792 19740
rect 16500 19712 16528 19740
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 21821 19771 21879 19777
rect 21821 19768 21833 19771
rect 19392 19740 21833 19768
rect 19392 19728 19398 19740
rect 21821 19737 21833 19740
rect 21867 19737 21879 19771
rect 22002 19768 22008 19780
rect 21963 19740 22008 19768
rect 21821 19731 21879 19737
rect 22002 19728 22008 19740
rect 22060 19728 22066 19780
rect 23201 19771 23259 19777
rect 23201 19768 23213 19771
rect 22296 19740 23213 19768
rect 16301 19703 16359 19709
rect 16301 19700 16313 19703
rect 15764 19672 16313 19700
rect 16301 19669 16313 19672
rect 16347 19669 16359 19703
rect 16301 19663 16359 19669
rect 16482 19660 16488 19712
rect 16540 19700 16546 19712
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 16540 19672 17509 19700
rect 16540 19660 16546 19672
rect 17497 19669 17509 19672
rect 17543 19669 17555 19703
rect 17497 19663 17555 19669
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19978 19700 19984 19712
rect 19751 19672 19984 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 22296 19700 22324 19740
rect 23201 19737 23213 19740
rect 23247 19737 23259 19771
rect 23201 19731 23259 19737
rect 23661 19771 23719 19777
rect 23661 19737 23673 19771
rect 23707 19737 23719 19771
rect 28828 19768 28856 19804
rect 23661 19731 23719 19737
rect 28736 19740 28856 19768
rect 29012 19768 29040 19808
rect 29086 19796 29092 19848
rect 29144 19836 29150 19848
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29144 19808 29561 19836
rect 29144 19796 29150 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 36078 19836 36084 19848
rect 29549 19799 29607 19805
rect 31726 19808 36084 19836
rect 31726 19768 31754 19808
rect 36078 19796 36084 19808
rect 36136 19796 36142 19848
rect 36170 19796 36176 19848
rect 36228 19836 36234 19848
rect 37829 19839 37887 19845
rect 37829 19836 37841 19839
rect 36228 19808 37841 19836
rect 36228 19796 36234 19808
rect 37829 19805 37841 19808
rect 37875 19805 37887 19839
rect 37829 19799 37887 19805
rect 33045 19771 33103 19777
rect 33045 19768 33057 19771
rect 29012 19740 31754 19768
rect 32416 19740 33057 19768
rect 21324 19672 22324 19700
rect 21324 19660 21330 19672
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 23566 19700 23572 19712
rect 22428 19672 22473 19700
rect 23527 19672 23572 19700
rect 22428 19660 22434 19672
rect 23566 19660 23572 19672
rect 23624 19660 23630 19712
rect 23676 19700 23704 19731
rect 28736 19700 28764 19740
rect 32416 19712 32444 19740
rect 33045 19737 33057 19740
rect 33091 19737 33103 19771
rect 33045 19731 33103 19737
rect 23676 19672 28764 19700
rect 28813 19703 28871 19709
rect 28813 19669 28825 19703
rect 28859 19700 28871 19703
rect 28902 19700 28908 19712
rect 28859 19672 28908 19700
rect 28859 19669 28871 19672
rect 28813 19663 28871 19669
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 32398 19700 32404 19712
rect 32359 19672 32404 19700
rect 32398 19660 32404 19672
rect 32456 19660 32462 19712
rect 36265 19703 36323 19709
rect 36265 19669 36277 19703
rect 36311 19700 36323 19703
rect 36354 19700 36360 19712
rect 36311 19672 36360 19700
rect 36311 19669 36323 19672
rect 36265 19663 36323 19669
rect 36354 19660 36360 19672
rect 36412 19660 36418 19712
rect 37369 19703 37427 19709
rect 37369 19669 37381 19703
rect 37415 19700 37427 19703
rect 38102 19700 38108 19712
rect 37415 19672 38108 19700
rect 37415 19669 37427 19672
rect 37369 19663 37427 19669
rect 38102 19660 38108 19672
rect 38160 19660 38166 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3053 19499 3111 19505
rect 3053 19465 3065 19499
rect 3099 19496 3111 19499
rect 3694 19496 3700 19508
rect 3099 19468 3700 19496
rect 3099 19465 3111 19468
rect 3053 19459 3111 19465
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 15654 19496 15660 19508
rect 15335 19468 15660 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 15654 19456 15660 19468
rect 15712 19496 15718 19508
rect 19242 19496 19248 19508
rect 15712 19468 19248 19496
rect 15712 19456 15718 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20254 19456 20260 19508
rect 20312 19496 20318 19508
rect 22370 19496 22376 19508
rect 20312 19468 22376 19496
rect 20312 19456 20318 19468
rect 22370 19456 22376 19468
rect 22428 19496 22434 19508
rect 23477 19499 23535 19505
rect 23477 19496 23489 19499
rect 22428 19468 23489 19496
rect 22428 19456 22434 19468
rect 23477 19465 23489 19468
rect 23523 19496 23535 19499
rect 23566 19496 23572 19508
rect 23523 19468 23572 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 29086 19496 29092 19508
rect 29047 19468 29092 19496
rect 29086 19456 29092 19468
rect 29144 19456 29150 19508
rect 3878 19388 3884 19440
rect 3936 19428 3942 19440
rect 13722 19428 13728 19440
rect 3936 19400 13728 19428
rect 3936 19388 3942 19400
rect 13722 19388 13728 19400
rect 13780 19388 13786 19440
rect 16666 19388 16672 19440
rect 16724 19428 16730 19440
rect 18874 19428 18880 19440
rect 16724 19400 18880 19428
rect 16724 19388 16730 19400
rect 18874 19388 18880 19400
rect 18932 19428 18938 19440
rect 22922 19428 22928 19440
rect 18932 19400 22928 19428
rect 18932 19388 18938 19400
rect 22922 19388 22928 19400
rect 22980 19388 22986 19440
rect 24670 19428 24676 19440
rect 23584 19400 24676 19428
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2866 19360 2872 19372
rect 2731 19332 2872 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2866 19320 2872 19332
rect 2924 19360 2930 19372
rect 3513 19363 3571 19369
rect 3513 19360 3525 19363
rect 2924 19332 3525 19360
rect 2924 19320 2930 19332
rect 3513 19329 3525 19332
rect 3559 19329 3571 19363
rect 3513 19323 3571 19329
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 13906 19360 13912 19372
rect 13867 19332 13912 19360
rect 3697 19323 3755 19329
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 2958 19292 2964 19304
rect 2823 19264 2964 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3712 19292 3740 19323
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 14182 19369 14188 19372
rect 14176 19323 14188 19369
rect 14240 19360 14246 19372
rect 14240 19332 14276 19360
rect 14182 19320 14188 19323
rect 14240 19320 14246 19332
rect 20162 19320 20168 19372
rect 20220 19360 20226 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20220 19332 20729 19360
rect 20220 19320 20226 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 21082 19360 21088 19372
rect 21039 19332 21088 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 23584 19369 23612 19400
rect 24670 19388 24676 19400
rect 24728 19388 24734 19440
rect 27614 19428 27620 19440
rect 27575 19400 27620 19428
rect 27614 19388 27620 19400
rect 27672 19388 27678 19440
rect 36078 19388 36084 19440
rect 36136 19428 36142 19440
rect 36136 19400 37872 19428
rect 36136 19388 36142 19400
rect 21177 19363 21235 19369
rect 21177 19329 21189 19363
rect 21223 19360 21235 19363
rect 23109 19363 23167 19369
rect 23109 19360 23121 19363
rect 21223 19332 23121 19360
rect 21223 19329 21235 19332
rect 21177 19323 21235 19329
rect 23109 19329 23121 19332
rect 23155 19329 23167 19363
rect 23109 19323 23167 19329
rect 23569 19363 23627 19369
rect 23569 19329 23581 19363
rect 23615 19329 23627 19363
rect 23569 19323 23627 19329
rect 23661 19363 23719 19369
rect 23661 19329 23673 19363
rect 23707 19360 23719 19363
rect 24302 19360 24308 19372
rect 23707 19332 24308 19360
rect 23707 19329 23719 19332
rect 23661 19323 23719 19329
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 27801 19363 27859 19369
rect 27801 19360 27813 19363
rect 27632 19332 27813 19360
rect 3108 19264 3740 19292
rect 19613 19295 19671 19301
rect 3108 19252 3114 19264
rect 19613 19261 19625 19295
rect 19659 19292 19671 19295
rect 19978 19292 19984 19304
rect 19659 19264 19984 19292
rect 19659 19261 19671 19264
rect 19613 19255 19671 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 20901 19295 20959 19301
rect 20901 19292 20913 19295
rect 20680 19264 20913 19292
rect 20680 19252 20686 19264
rect 20901 19261 20913 19264
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 23368 19295 23426 19301
rect 23368 19261 23380 19295
rect 23414 19292 23426 19295
rect 23414 19264 23520 19292
rect 23414 19261 23426 19264
rect 23368 19255 23426 19261
rect 2133 19227 2191 19233
rect 2133 19193 2145 19227
rect 2179 19224 2191 19227
rect 9306 19224 9312 19236
rect 2179 19196 9312 19224
rect 2179 19193 2191 19196
rect 2133 19187 2191 19193
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 18690 19184 18696 19236
rect 18748 19224 18754 19236
rect 18877 19227 18935 19233
rect 18877 19224 18889 19227
rect 18748 19196 18889 19224
rect 18748 19184 18754 19196
rect 18877 19193 18889 19196
rect 18923 19224 18935 19227
rect 20806 19224 20812 19236
rect 18923 19196 19748 19224
rect 20767 19196 20812 19224
rect 18923 19193 18935 19196
rect 18877 19187 18935 19193
rect 2869 19159 2927 19165
rect 2869 19125 2881 19159
rect 2915 19156 2927 19159
rect 3050 19156 3056 19168
rect 2915 19128 3056 19156
rect 2915 19125 2927 19128
rect 2869 19119 2927 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3786 19116 3792 19168
rect 3844 19156 3850 19168
rect 3881 19159 3939 19165
rect 3881 19156 3893 19159
rect 3844 19128 3893 19156
rect 3844 19116 3850 19128
rect 3881 19125 3893 19128
rect 3927 19125 3939 19159
rect 3881 19119 3939 19125
rect 16025 19159 16083 19165
rect 16025 19125 16037 19159
rect 16071 19156 16083 19159
rect 16482 19156 16488 19168
rect 16071 19128 16488 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 16666 19156 16672 19168
rect 16627 19128 16672 19156
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 19720 19156 19748 19196
rect 20806 19184 20812 19196
rect 20864 19184 20870 19236
rect 22922 19224 22928 19236
rect 22883 19196 22928 19224
rect 22922 19184 22928 19196
rect 22980 19184 22986 19236
rect 23492 19224 23520 19264
rect 23842 19224 23848 19236
rect 23492 19196 23848 19224
rect 23842 19184 23848 19196
rect 23900 19184 23906 19236
rect 27632 19168 27660 19332
rect 27801 19329 27813 19332
rect 27847 19329 27859 19363
rect 36446 19360 36452 19372
rect 36407 19332 36452 19360
rect 27801 19323 27859 19329
rect 36446 19320 36452 19332
rect 36504 19320 36510 19372
rect 37844 19369 37872 19400
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 28626 19292 28632 19304
rect 28587 19264 28632 19292
rect 28626 19252 28632 19264
rect 28684 19252 28690 19304
rect 36725 19295 36783 19301
rect 36725 19292 36737 19295
rect 36372 19264 36737 19292
rect 28902 19224 28908 19236
rect 28863 19196 28908 19224
rect 28902 19184 28908 19196
rect 28960 19184 28966 19236
rect 36372 19168 36400 19264
rect 36725 19261 36737 19264
rect 36771 19261 36783 19295
rect 36725 19255 36783 19261
rect 22278 19156 22284 19168
rect 19720 19128 22284 19156
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 23382 19116 23388 19168
rect 23440 19156 23446 19168
rect 23934 19156 23940 19168
rect 23440 19128 23940 19156
rect 23440 19116 23446 19128
rect 23934 19116 23940 19128
rect 23992 19116 23998 19168
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19156 27215 19159
rect 27614 19156 27620 19168
rect 27203 19128 27620 19156
rect 27203 19125 27215 19128
rect 27157 19119 27215 19125
rect 27614 19116 27620 19128
rect 27672 19116 27678 19168
rect 34790 19156 34796 19168
rect 34751 19128 34796 19156
rect 34790 19116 34796 19128
rect 34848 19116 34854 19168
rect 35437 19159 35495 19165
rect 35437 19125 35449 19159
rect 35483 19156 35495 19159
rect 36354 19156 36360 19168
rect 35483 19128 36360 19156
rect 35483 19125 35495 19128
rect 35437 19119 35495 19125
rect 36354 19116 36360 19128
rect 36412 19116 36418 19168
rect 37274 19156 37280 19168
rect 37235 19128 37280 19156
rect 37274 19116 37280 19128
rect 37332 19116 37338 19168
rect 38010 19156 38016 19168
rect 37971 19128 38016 19156
rect 38010 19116 38016 19128
rect 38068 19116 38074 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 2777 18955 2835 18961
rect 2777 18921 2789 18955
rect 2823 18952 2835 18955
rect 3050 18952 3056 18964
rect 2823 18924 3056 18952
rect 2823 18921 2835 18924
rect 2777 18915 2835 18921
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 3510 18912 3516 18964
rect 3568 18952 3574 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3568 18924 3801 18952
rect 3568 18912 3574 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 15381 18955 15439 18961
rect 15381 18921 15393 18955
rect 15427 18952 15439 18955
rect 15930 18952 15936 18964
rect 15427 18924 15936 18952
rect 15427 18921 15439 18924
rect 15381 18915 15439 18921
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18921 20039 18955
rect 20162 18952 20168 18964
rect 20123 18924 20168 18952
rect 19981 18915 20039 18921
rect 2866 18884 2872 18896
rect 2792 18856 2872 18884
rect 2792 18825 2820 18856
rect 2866 18844 2872 18856
rect 2924 18844 2930 18896
rect 4062 18844 4068 18896
rect 4120 18884 4126 18896
rect 19334 18884 19340 18896
rect 4120 18856 19340 18884
rect 4120 18844 4126 18856
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 19996 18884 20024 18915
rect 20162 18912 20168 18924
rect 20220 18912 20226 18964
rect 21177 18955 21235 18961
rect 21177 18921 21189 18955
rect 21223 18952 21235 18955
rect 22002 18952 22008 18964
rect 21223 18924 22008 18952
rect 21223 18921 21235 18924
rect 21177 18915 21235 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22186 18952 22192 18964
rect 22147 18924 22192 18952
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 20714 18884 20720 18896
rect 19996 18856 20720 18884
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 20809 18887 20867 18893
rect 20809 18853 20821 18887
rect 20855 18884 20867 18887
rect 20898 18884 20904 18896
rect 20855 18856 20904 18884
rect 20855 18853 20867 18856
rect 20809 18847 20867 18853
rect 20898 18844 20904 18856
rect 20956 18884 20962 18896
rect 21821 18887 21879 18893
rect 21821 18884 21833 18887
rect 20956 18856 21833 18884
rect 20956 18844 20962 18856
rect 21821 18853 21833 18856
rect 21867 18853 21879 18887
rect 37826 18884 37832 18896
rect 21821 18847 21879 18853
rect 35912 18856 37832 18884
rect 2777 18819 2835 18825
rect 2777 18785 2789 18819
rect 2823 18785 2835 18819
rect 2777 18779 2835 18785
rect 3326 18776 3332 18828
rect 3384 18816 3390 18828
rect 3881 18819 3939 18825
rect 3881 18816 3893 18819
rect 3384 18788 3893 18816
rect 3384 18776 3390 18788
rect 3881 18785 3893 18788
rect 3927 18785 3939 18819
rect 3881 18779 3939 18785
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 19426 18816 19432 18828
rect 4028 18788 19432 18816
rect 4028 18776 4034 18788
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 20438 18816 20444 18828
rect 19904 18788 20444 18816
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18748 2927 18751
rect 3050 18748 3056 18760
rect 2915 18720 3056 18748
rect 2915 18717 2927 18720
rect 2869 18711 2927 18717
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 3786 18748 3792 18760
rect 3747 18720 3792 18748
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14458 18748 14464 18760
rect 14323 18720 14464 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 2409 18683 2467 18689
rect 2409 18680 2421 18683
rect 1596 18652 2421 18680
rect 1596 18621 1624 18652
rect 2409 18649 2421 18652
rect 2455 18680 2467 18683
rect 2958 18680 2964 18692
rect 2455 18652 2964 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 2958 18640 2964 18652
rect 3016 18680 3022 18692
rect 4080 18680 4108 18711
rect 14458 18708 14464 18720
rect 14516 18748 14522 18760
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14516 18720 14749 18748
rect 14516 18708 14522 18720
rect 14737 18717 14749 18720
rect 14783 18717 14795 18751
rect 14918 18748 14924 18760
rect 14879 18720 14924 18748
rect 14737 18711 14795 18717
rect 3016 18652 4108 18680
rect 3016 18640 3022 18652
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 13354 18680 13360 18692
rect 7524 18652 12434 18680
rect 13315 18652 13360 18680
rect 7524 18640 7530 18652
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 3053 18615 3111 18621
rect 3053 18581 3065 18615
rect 3099 18612 3111 18615
rect 3234 18612 3240 18624
rect 3099 18584 3240 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 5442 18612 5448 18624
rect 4295 18584 5448 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11848 18584 11989 18612
rect 11848 18572 11854 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 12406 18612 12434 18652
rect 13354 18640 13360 18652
rect 13412 18640 13418 18692
rect 13541 18683 13599 18689
rect 13541 18649 13553 18683
rect 13587 18680 13599 18683
rect 14550 18680 14556 18692
rect 13587 18652 14556 18680
rect 13587 18649 13599 18652
rect 13541 18643 13599 18649
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 14752 18680 14780 18711
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 15194 18748 15200 18760
rect 15155 18720 15200 18748
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 18230 18708 18236 18760
rect 18288 18748 18294 18760
rect 19904 18757 19932 18788
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 35912 18825 35940 18856
rect 37826 18844 37832 18856
rect 37884 18844 37890 18896
rect 35897 18819 35955 18825
rect 35897 18785 35909 18819
rect 35943 18785 35955 18819
rect 35897 18779 35955 18785
rect 37185 18819 37243 18825
rect 37185 18785 37197 18819
rect 37231 18816 37243 18819
rect 37366 18816 37372 18828
rect 37231 18788 37372 18816
rect 37231 18785 37243 18788
rect 37185 18779 37243 18785
rect 37366 18776 37372 18788
rect 37424 18776 37430 18828
rect 19889 18751 19947 18757
rect 18288 18720 19840 18748
rect 18288 18708 18294 18720
rect 16298 18680 16304 18692
rect 14752 18652 16304 18680
rect 16298 18640 16304 18652
rect 16356 18640 16362 18692
rect 19702 18680 19708 18692
rect 19663 18652 19708 18680
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 19812 18680 19840 18720
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 20021 18751 20079 18757
rect 20021 18717 20033 18751
rect 20067 18748 20079 18751
rect 20162 18748 20168 18760
rect 20067 18720 20168 18748
rect 20067 18717 20079 18720
rect 20021 18711 20079 18717
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18717 21051 18751
rect 21726 18748 21732 18760
rect 21687 18720 21732 18748
rect 20993 18711 21051 18717
rect 20622 18680 20628 18692
rect 19812 18652 20628 18680
rect 20622 18640 20628 18652
rect 20680 18680 20686 18692
rect 20916 18680 20944 18711
rect 20680 18652 20944 18680
rect 21008 18680 21036 18711
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 21910 18748 21916 18760
rect 21871 18720 21916 18748
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18717 22063 18751
rect 27706 18748 27712 18760
rect 27619 18720 27712 18748
rect 22005 18711 22063 18717
rect 22020 18680 22048 18711
rect 27706 18708 27712 18720
rect 27764 18748 27770 18760
rect 28074 18748 28080 18760
rect 27764 18720 28080 18748
rect 27764 18708 27770 18720
rect 28074 18708 28080 18720
rect 28132 18748 28138 18760
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 28132 18720 28181 18748
rect 28132 18708 28138 18720
rect 28169 18717 28181 18720
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 28445 18751 28503 18757
rect 28445 18717 28457 18751
rect 28491 18748 28503 18751
rect 28626 18748 28632 18760
rect 28491 18720 28632 18748
rect 28491 18717 28503 18720
rect 28445 18711 28503 18717
rect 28626 18708 28632 18720
rect 28684 18748 28690 18760
rect 30098 18748 30104 18760
rect 28684 18720 30104 18748
rect 28684 18708 28690 18720
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 32398 18748 32404 18760
rect 31864 18720 32404 18748
rect 24854 18680 24860 18692
rect 21008 18652 22048 18680
rect 24815 18652 24860 18680
rect 20680 18640 20686 18652
rect 16666 18612 16672 18624
rect 12406 18584 16672 18612
rect 11977 18575 12035 18581
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 21008 18612 21036 18652
rect 24854 18640 24860 18652
rect 24912 18640 24918 18692
rect 25038 18640 25044 18692
rect 25096 18680 25102 18692
rect 25774 18680 25780 18692
rect 25096 18652 25780 18680
rect 25096 18640 25102 18652
rect 25774 18640 25780 18652
rect 25832 18640 25838 18692
rect 31864 18624 31892 18720
rect 32398 18708 32404 18720
rect 32456 18708 32462 18760
rect 36173 18751 36231 18757
rect 36173 18717 36185 18751
rect 36219 18717 36231 18751
rect 36173 18711 36231 18717
rect 21082 18612 21088 18624
rect 17552 18584 21088 18612
rect 17552 18572 17558 18584
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 26881 18615 26939 18621
rect 26881 18581 26893 18615
rect 26927 18612 26939 18615
rect 27614 18612 27620 18624
rect 26927 18584 27620 18612
rect 26927 18581 26939 18584
rect 26881 18575 26939 18581
rect 27614 18572 27620 18584
rect 27672 18572 27678 18624
rect 31846 18612 31852 18624
rect 31807 18584 31852 18612
rect 31846 18572 31852 18584
rect 31904 18572 31910 18624
rect 32582 18612 32588 18624
rect 32543 18584 32588 18612
rect 32582 18572 32588 18584
rect 32640 18572 32646 18624
rect 34790 18572 34796 18624
rect 34848 18612 34854 18624
rect 34885 18615 34943 18621
rect 34885 18612 34897 18615
rect 34848 18584 34897 18612
rect 34848 18572 34854 18584
rect 34885 18581 34897 18584
rect 34931 18612 34943 18615
rect 35710 18612 35716 18624
rect 34931 18584 35716 18612
rect 34931 18581 34943 18584
rect 34885 18575 34943 18581
rect 35710 18572 35716 18584
rect 35768 18612 35774 18624
rect 36188 18612 36216 18711
rect 37274 18708 37280 18760
rect 37332 18748 37338 18760
rect 37461 18751 37519 18757
rect 37461 18748 37473 18751
rect 37332 18720 37473 18748
rect 37332 18708 37338 18720
rect 37461 18717 37473 18720
rect 37507 18717 37519 18751
rect 38102 18748 38108 18760
rect 38063 18720 38108 18748
rect 37461 18711 37519 18717
rect 38102 18708 38108 18720
rect 38160 18708 38166 18760
rect 35768 18584 36216 18612
rect 35768 18572 35774 18584
rect 37366 18572 37372 18624
rect 37424 18612 37430 18624
rect 37921 18615 37979 18621
rect 37921 18612 37933 18615
rect 37424 18584 37933 18612
rect 37424 18572 37430 18584
rect 37921 18581 37933 18584
rect 37967 18581 37979 18615
rect 37921 18575 37979 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1394 18368 1400 18420
rect 1452 18408 1458 18420
rect 2685 18411 2743 18417
rect 2685 18408 2697 18411
rect 1452 18380 2697 18408
rect 1452 18368 1458 18380
rect 2685 18377 2697 18380
rect 2731 18377 2743 18411
rect 10318 18408 10324 18420
rect 2685 18371 2743 18377
rect 9232 18380 10324 18408
rect 2222 18340 2228 18352
rect 2183 18312 2228 18340
rect 2222 18300 2228 18312
rect 2280 18300 2286 18352
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 3234 18272 3240 18284
rect 3195 18244 3240 18272
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 3326 18232 3332 18284
rect 3384 18272 3390 18284
rect 3510 18272 3516 18284
rect 3384 18244 3429 18272
rect 3471 18244 3516 18272
rect 3384 18232 3390 18244
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 9232 18281 9260 18380
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 13446 18408 13452 18420
rect 13407 18380 13452 18408
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 14182 18408 14188 18420
rect 14143 18380 14188 18408
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 19978 18408 19984 18420
rect 17000 18380 19984 18408
rect 17000 18368 17006 18380
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20257 18411 20315 18417
rect 20257 18377 20269 18411
rect 20303 18408 20315 18411
rect 21266 18408 21272 18420
rect 20303 18380 20852 18408
rect 21227 18380 21272 18408
rect 20303 18377 20315 18380
rect 20257 18371 20315 18377
rect 9306 18300 9312 18352
rect 9364 18340 9370 18352
rect 17126 18340 17132 18352
rect 9364 18312 17132 18340
rect 9364 18300 9370 18312
rect 17126 18300 17132 18312
rect 17184 18300 17190 18352
rect 18785 18343 18843 18349
rect 18785 18309 18797 18343
rect 18831 18340 18843 18343
rect 19426 18340 19432 18352
rect 18831 18312 19432 18340
rect 18831 18309 18843 18312
rect 18785 18303 18843 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 20530 18340 20536 18352
rect 20171 18312 20536 18340
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18241 9275 18275
rect 9490 18272 9496 18284
rect 9451 18244 9496 18272
rect 9217 18235 9275 18241
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 10042 18272 10048 18284
rect 9723 18244 10048 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 12342 18272 12348 18284
rect 12303 18244 12348 18272
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 13170 18272 13176 18284
rect 12544 18244 13176 18272
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18173 4031 18207
rect 12544 18204 12572 18244
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18241 13415 18275
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 13357 18235 13415 18241
rect 3973 18167 4031 18173
rect 9416 18176 12572 18204
rect 3988 18136 4016 18167
rect 3988 18108 9260 18136
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9122 18068 9128 18080
rect 9079 18040 9128 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 9232 18068 9260 18108
rect 9416 18068 9444 18176
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12676 18176 12721 18204
rect 12676 18164 12682 18176
rect 12437 18139 12495 18145
rect 12437 18105 12449 18139
rect 12483 18136 12495 18139
rect 13262 18136 13268 18148
rect 12483 18108 13268 18136
rect 12483 18105 12495 18108
rect 12437 18099 12495 18105
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 9232 18040 9444 18068
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10137 18071 10195 18077
rect 10137 18068 10149 18071
rect 10100 18040 10149 18068
rect 10100 18028 10106 18040
rect 10137 18037 10149 18040
rect 10183 18037 10195 18071
rect 10137 18031 10195 18037
rect 10226 18028 10232 18080
rect 10284 18068 10290 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10284 18040 10701 18068
rect 10284 18028 10290 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 10689 18031 10747 18037
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18068 11759 18071
rect 11790 18068 11796 18080
rect 11747 18040 11796 18068
rect 11747 18037 11759 18040
rect 11701 18031 11759 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12250 18028 12256 18080
rect 12308 18068 12314 18080
rect 12529 18071 12587 18077
rect 12529 18068 12541 18071
rect 12308 18040 12541 18068
rect 12308 18028 12314 18040
rect 12529 18037 12541 18040
rect 12575 18068 12587 18071
rect 13372 18068 13400 18235
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 19794 18232 19800 18284
rect 19852 18272 19858 18284
rect 20171 18281 20199 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 20824 18281 20852 18380
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 21726 18368 21732 18420
rect 21784 18408 21790 18420
rect 22281 18411 22339 18417
rect 22281 18408 22293 18411
rect 21784 18380 22293 18408
rect 21784 18368 21790 18380
rect 22281 18377 22293 18380
rect 22327 18377 22339 18411
rect 22281 18371 22339 18377
rect 20990 18300 20996 18352
rect 21048 18340 21054 18352
rect 25685 18343 25743 18349
rect 25685 18340 25697 18343
rect 21048 18312 25697 18340
rect 21048 18300 21054 18312
rect 25685 18309 25697 18312
rect 25731 18309 25743 18343
rect 25685 18303 25743 18309
rect 25869 18343 25927 18349
rect 25869 18309 25881 18343
rect 25915 18340 25927 18343
rect 27522 18340 27528 18352
rect 25915 18312 27528 18340
rect 25915 18309 25927 18312
rect 25869 18303 25927 18309
rect 27522 18300 27528 18312
rect 27580 18300 27586 18352
rect 20113 18275 20199 18281
rect 19852 18244 19897 18272
rect 19852 18232 19858 18244
rect 20113 18241 20125 18275
rect 20159 18244 20199 18275
rect 20809 18275 20867 18281
rect 20159 18241 20171 18244
rect 20113 18235 20171 18241
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 20956 18244 21001 18272
rect 20956 18232 20962 18244
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 21140 18244 21185 18272
rect 21140 18232 21146 18244
rect 21450 18232 21456 18284
rect 21508 18272 21514 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21508 18244 21833 18272
rect 21508 18232 21514 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18272 22155 18275
rect 22186 18272 22192 18284
rect 22143 18244 22192 18272
rect 22143 18241 22155 18244
rect 22097 18235 22155 18241
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 25958 18232 25964 18284
rect 26016 18272 26022 18284
rect 26053 18275 26111 18281
rect 26053 18272 26065 18275
rect 26016 18244 26065 18272
rect 26016 18232 26022 18244
rect 26053 18241 26065 18244
rect 26099 18241 26111 18275
rect 26053 18235 26111 18241
rect 26973 18275 27031 18281
rect 26973 18241 26985 18275
rect 27019 18272 27031 18275
rect 27614 18272 27620 18284
rect 27019 18244 27620 18272
rect 27019 18241 27031 18244
rect 26973 18235 27031 18241
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 30929 18275 30987 18281
rect 30929 18272 30941 18275
rect 30484 18244 30941 18272
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 14240 18176 14657 18204
rect 14240 18164 14246 18176
rect 14645 18173 14657 18176
rect 14691 18204 14703 18207
rect 19610 18204 19616 18216
rect 14691 18176 19616 18204
rect 14691 18173 14703 18176
rect 14645 18167 14703 18173
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 19886 18204 19892 18216
rect 19847 18176 19892 18204
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 20438 18164 20444 18216
rect 20496 18204 20502 18216
rect 21910 18204 21916 18216
rect 20496 18176 21916 18204
rect 20496 18164 20502 18176
rect 21910 18164 21916 18176
rect 21968 18164 21974 18216
rect 24489 18207 24547 18213
rect 24489 18204 24501 18207
rect 22066 18176 24501 18204
rect 13538 18096 13544 18148
rect 13596 18136 13602 18148
rect 13596 18108 19932 18136
rect 13596 18096 13602 18108
rect 12575 18040 13400 18068
rect 12575 18037 12587 18040
rect 12529 18031 12587 18037
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19794 18068 19800 18080
rect 19392 18040 19437 18068
rect 19755 18040 19800 18068
rect 19392 18028 19398 18040
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 19904 18068 19932 18108
rect 20622 18096 20628 18148
rect 20680 18136 20686 18148
rect 20993 18139 21051 18145
rect 20993 18136 21005 18139
rect 20680 18108 21005 18136
rect 20680 18096 20686 18108
rect 20993 18105 21005 18108
rect 21039 18105 21051 18139
rect 22066 18136 22094 18176
rect 24489 18173 24501 18176
rect 24535 18204 24547 18207
rect 24946 18204 24952 18216
rect 24535 18176 24952 18204
rect 24535 18173 24547 18176
rect 24489 18167 24547 18173
rect 24946 18164 24952 18176
rect 25004 18164 25010 18216
rect 27154 18164 27160 18216
rect 27212 18204 27218 18216
rect 28258 18204 28264 18216
rect 27212 18176 28264 18204
rect 27212 18164 27218 18176
rect 28258 18164 28264 18176
rect 28316 18164 28322 18216
rect 30009 18207 30067 18213
rect 30009 18173 30021 18207
rect 30055 18204 30067 18207
rect 30098 18204 30104 18216
rect 30055 18176 30104 18204
rect 30055 18173 30067 18176
rect 30009 18167 30067 18173
rect 30098 18164 30104 18176
rect 30156 18164 30162 18216
rect 30484 18213 30512 18244
rect 30929 18241 30941 18244
rect 30975 18241 30987 18275
rect 34514 18272 34520 18284
rect 34475 18244 34520 18272
rect 30929 18235 30987 18241
rect 34514 18232 34520 18244
rect 34572 18232 34578 18284
rect 35710 18272 35716 18284
rect 35671 18244 35716 18272
rect 35710 18232 35716 18244
rect 35768 18232 35774 18284
rect 36354 18232 36360 18284
rect 36412 18272 36418 18284
rect 36449 18275 36507 18281
rect 36449 18272 36461 18275
rect 36412 18244 36461 18272
rect 36412 18232 36418 18244
rect 36449 18241 36461 18244
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 37829 18275 37887 18281
rect 37829 18241 37841 18275
rect 37875 18241 37887 18275
rect 37829 18235 37887 18241
rect 30469 18207 30527 18213
rect 30469 18173 30481 18207
rect 30515 18173 30527 18207
rect 30469 18167 30527 18173
rect 32306 18164 32312 18216
rect 32364 18204 32370 18216
rect 37844 18204 37872 18235
rect 32364 18176 37872 18204
rect 32364 18164 32370 18176
rect 20993 18099 21051 18105
rect 21100 18108 22094 18136
rect 21100 18068 21128 18108
rect 24210 18096 24216 18148
rect 24268 18136 24274 18148
rect 25038 18136 25044 18148
rect 24268 18108 25044 18136
rect 24268 18096 24274 18108
rect 25038 18096 25044 18108
rect 25096 18096 25102 18148
rect 29270 18136 29276 18148
rect 25148 18108 29276 18136
rect 19904 18040 21128 18068
rect 21726 18028 21732 18080
rect 21784 18068 21790 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 21784 18040 21833 18068
rect 21784 18028 21790 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 21821 18031 21879 18037
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 22833 18071 22891 18077
rect 22833 18068 22845 18071
rect 22244 18040 22845 18068
rect 22244 18028 22250 18040
rect 22833 18037 22845 18040
rect 22879 18068 22891 18071
rect 25148 18068 25176 18108
rect 29270 18096 29276 18108
rect 29328 18096 29334 18148
rect 30282 18136 30288 18148
rect 30243 18108 30288 18136
rect 30282 18096 30288 18108
rect 30340 18096 30346 18148
rect 35802 18096 35808 18148
rect 35860 18136 35866 18148
rect 35897 18139 35955 18145
rect 35897 18136 35909 18139
rect 35860 18108 35909 18136
rect 35860 18096 35866 18108
rect 35897 18105 35909 18108
rect 35943 18136 35955 18139
rect 36262 18136 36268 18148
rect 35943 18108 36268 18136
rect 35943 18105 35955 18108
rect 35897 18099 35955 18105
rect 36262 18096 36268 18108
rect 36320 18096 36326 18148
rect 36630 18136 36636 18148
rect 36591 18108 36636 18136
rect 36630 18096 36636 18108
rect 36688 18096 36694 18148
rect 22879 18040 25176 18068
rect 27157 18071 27215 18077
rect 22879 18037 22891 18040
rect 22833 18031 22891 18037
rect 27157 18037 27169 18071
rect 27203 18068 27215 18071
rect 27246 18068 27252 18080
rect 27203 18040 27252 18068
rect 27203 18037 27215 18040
rect 27157 18031 27215 18037
rect 27246 18028 27252 18040
rect 27304 18028 27310 18080
rect 31110 18068 31116 18080
rect 31071 18040 31116 18068
rect 31110 18028 31116 18040
rect 31168 18028 31174 18080
rect 34701 18071 34759 18077
rect 34701 18037 34713 18071
rect 34747 18068 34759 18071
rect 34790 18068 34796 18080
rect 34747 18040 34796 18068
rect 34747 18037 34759 18040
rect 34701 18031 34759 18037
rect 34790 18028 34796 18040
rect 34848 18028 34854 18080
rect 37274 18068 37280 18080
rect 37235 18040 37280 18068
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 38010 18068 38016 18080
rect 37971 18040 38016 18068
rect 38010 18028 38016 18040
rect 38068 18028 38074 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1486 17864 1492 17876
rect 1447 17836 1492 17864
rect 1486 17824 1492 17836
rect 1544 17824 1550 17876
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 3050 17864 3056 17876
rect 2363 17836 3056 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3568 17836 4077 17864
rect 3568 17824 3574 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 9640 17836 11468 17864
rect 9640 17824 9646 17836
rect 3326 17756 3332 17808
rect 3384 17796 3390 17808
rect 3927 17799 3985 17805
rect 3927 17796 3939 17799
rect 3384 17768 3939 17796
rect 3384 17756 3390 17768
rect 3927 17765 3939 17768
rect 3973 17765 3985 17799
rect 3927 17759 3985 17765
rect 6362 17756 6368 17808
rect 6420 17796 6426 17808
rect 7101 17799 7159 17805
rect 7101 17796 7113 17799
rect 6420 17768 7113 17796
rect 6420 17756 6426 17768
rect 7101 17765 7113 17768
rect 7147 17796 7159 17799
rect 11054 17796 11060 17808
rect 7147 17768 11060 17796
rect 7147 17765 7159 17768
rect 7101 17759 7159 17765
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 11440 17805 11468 17836
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12161 17867 12219 17873
rect 12161 17864 12173 17867
rect 12124 17836 12173 17864
rect 12124 17824 12130 17836
rect 12161 17833 12173 17836
rect 12207 17864 12219 17867
rect 12434 17864 12440 17876
rect 12207 17836 12440 17864
rect 12207 17833 12219 17836
rect 12161 17827 12219 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 13446 17864 13452 17876
rect 12676 17836 13452 17864
rect 12676 17824 12682 17836
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 14182 17864 14188 17876
rect 14143 17836 14188 17864
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 19794 17824 19800 17876
rect 19852 17864 19858 17876
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 19852 17836 20637 17864
rect 19852 17824 19858 17836
rect 20625 17833 20637 17836
rect 20671 17833 20683 17867
rect 20625 17827 20683 17833
rect 11425 17799 11483 17805
rect 11425 17765 11437 17799
rect 11471 17796 11483 17799
rect 12529 17799 12587 17805
rect 11471 17768 12480 17796
rect 11471 17765 11483 17768
rect 11425 17759 11483 17765
rect 3145 17731 3203 17737
rect 3145 17697 3157 17731
rect 3191 17728 3203 17731
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 3191 17700 4169 17728
rect 3191 17697 3203 17700
rect 3145 17691 3203 17697
rect 4157 17697 4169 17700
rect 4203 17728 4215 17731
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 4203 17700 7205 17728
rect 4203 17697 4215 17700
rect 4157 17691 4215 17697
rect 7193 17697 7205 17700
rect 7239 17728 7251 17731
rect 7374 17728 7380 17740
rect 7239 17700 7380 17728
rect 7239 17697 7251 17700
rect 7193 17691 7251 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17728 9827 17731
rect 10134 17728 10140 17740
rect 9815 17700 10140 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 12452 17728 12480 17768
rect 12529 17765 12541 17799
rect 12575 17796 12587 17799
rect 20640 17796 20668 17827
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 20809 17867 20867 17873
rect 20809 17864 20821 17867
rect 20772 17836 20821 17864
rect 20772 17824 20778 17836
rect 20809 17833 20821 17836
rect 20855 17833 20867 17867
rect 20809 17827 20867 17833
rect 22005 17867 22063 17873
rect 22005 17833 22017 17867
rect 22051 17864 22063 17867
rect 22554 17864 22560 17876
rect 22051 17836 22560 17864
rect 22051 17833 22063 17836
rect 22005 17827 22063 17833
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 28169 17867 28227 17873
rect 28169 17864 28181 17867
rect 27672 17836 28181 17864
rect 27672 17824 27678 17836
rect 28169 17833 28181 17836
rect 28215 17833 28227 17867
rect 28169 17827 28227 17833
rect 12575 17768 20576 17796
rect 20640 17768 20760 17796
rect 12575 17765 12587 17768
rect 12529 17759 12587 17765
rect 13538 17728 13544 17740
rect 12452 17700 13544 17728
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17728 17187 17731
rect 19886 17728 19892 17740
rect 17175 17700 19892 17728
rect 17175 17697 17187 17700
rect 17129 17691 17187 17697
rect 19886 17688 19892 17700
rect 19944 17728 19950 17740
rect 20438 17728 20444 17740
rect 19944 17700 20444 17728
rect 19944 17688 19950 17700
rect 20438 17688 20444 17700
rect 20496 17688 20502 17740
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 1673 17623 1731 17629
rect 1688 17592 1716 17623
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3694 17620 3700 17672
rect 3752 17660 3758 17672
rect 3789 17663 3847 17669
rect 3789 17660 3801 17663
rect 3752 17632 3801 17660
rect 3752 17620 3758 17632
rect 3789 17629 3801 17632
rect 3835 17629 3847 17663
rect 3789 17623 3847 17629
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 6822 17660 6828 17672
rect 5500 17632 6828 17660
rect 5500 17620 5506 17632
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 6972 17663 7030 17669
rect 6972 17629 6984 17663
rect 7018 17660 7030 17663
rect 7282 17660 7288 17672
rect 7018 17632 7288 17660
rect 7018 17629 7030 17632
rect 6972 17623 7030 17629
rect 7282 17620 7288 17632
rect 7340 17620 7346 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10318 17660 10324 17672
rect 10091 17632 10324 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11146 17660 11152 17672
rect 11020 17632 11152 17660
rect 11020 17620 11026 17632
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 3326 17592 3332 17604
rect 1688 17564 3332 17592
rect 3326 17552 3332 17564
rect 3384 17552 3390 17604
rect 4525 17595 4583 17601
rect 4525 17561 4537 17595
rect 4571 17592 4583 17595
rect 7558 17592 7564 17604
rect 4571 17564 7420 17592
rect 7519 17564 7564 17592
rect 4571 17561 4583 17564
rect 4525 17555 4583 17561
rect 6362 17524 6368 17536
rect 6323 17496 6368 17524
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 7392 17524 7420 17564
rect 7558 17552 7564 17564
rect 7616 17552 7622 17604
rect 12176 17592 12204 17623
rect 10796 17564 12204 17592
rect 10796 17536 10824 17564
rect 10778 17524 10784 17536
rect 7392 17496 10784 17524
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 12268 17524 12296 17623
rect 15930 17620 15936 17672
rect 15988 17660 15994 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 15988 17632 16865 17660
rect 15988 17620 15994 17632
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 18782 17620 18788 17672
rect 18840 17660 18846 17672
rect 19337 17663 19395 17669
rect 19337 17660 19349 17663
rect 18840 17632 19349 17660
rect 18840 17620 18846 17632
rect 19337 17629 19349 17632
rect 19383 17660 19395 17663
rect 20070 17660 20076 17672
rect 19383 17632 20076 17660
rect 19383 17629 19395 17632
rect 19337 17623 19395 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20346 17660 20352 17672
rect 20307 17632 20352 17660
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 13170 17552 13176 17604
rect 13228 17592 13234 17604
rect 13357 17595 13415 17601
rect 13228 17564 13273 17592
rect 13228 17552 13234 17564
rect 13357 17561 13369 17595
rect 13403 17592 13415 17595
rect 13446 17592 13452 17604
rect 13403 17564 13452 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 16390 17552 16396 17604
rect 16448 17592 16454 17604
rect 19702 17592 19708 17604
rect 16448 17564 19708 17592
rect 16448 17552 16454 17564
rect 19702 17552 19708 17564
rect 19760 17592 19766 17604
rect 20364 17592 20392 17620
rect 19760 17564 20392 17592
rect 19760 17552 19766 17564
rect 11848 17496 12296 17524
rect 16117 17527 16175 17533
rect 11848 17484 11854 17496
rect 16117 17493 16129 17527
rect 16163 17524 16175 17527
rect 16298 17524 16304 17536
rect 16163 17496 16304 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 19889 17527 19947 17533
rect 19889 17524 19901 17527
rect 16632 17496 19901 17524
rect 16632 17484 16638 17496
rect 19889 17493 19901 17496
rect 19935 17524 19947 17527
rect 20438 17524 20444 17536
rect 19935 17496 20444 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20548 17524 20576 17768
rect 20732 17728 20760 17768
rect 20898 17756 20904 17808
rect 20956 17796 20962 17808
rect 21637 17799 21695 17805
rect 21637 17796 21649 17799
rect 20956 17768 21649 17796
rect 20956 17756 20962 17768
rect 21637 17765 21649 17768
rect 21683 17765 21695 17799
rect 21637 17759 21695 17765
rect 21910 17756 21916 17808
rect 21968 17796 21974 17808
rect 23014 17796 23020 17808
rect 21968 17768 23020 17796
rect 21968 17756 21974 17768
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 24673 17799 24731 17805
rect 24673 17765 24685 17799
rect 24719 17796 24731 17799
rect 25958 17796 25964 17808
rect 24719 17768 25964 17796
rect 24719 17765 24731 17768
rect 24673 17759 24731 17765
rect 25958 17756 25964 17768
rect 26016 17756 26022 17808
rect 20806 17728 20812 17740
rect 20719 17700 20812 17728
rect 20806 17688 20812 17700
rect 20864 17728 20870 17740
rect 21082 17728 21088 17740
rect 20864 17700 21088 17728
rect 20864 17688 20870 17700
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 22002 17728 22008 17740
rect 21744 17700 22008 17728
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 20680 17632 20725 17660
rect 20680 17620 20686 17632
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21744 17669 21772 17700
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 21324 17632 21557 17660
rect 21324 17620 21330 17632
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 21729 17663 21787 17669
rect 21729 17629 21741 17663
rect 21775 17629 21787 17663
rect 21729 17623 21787 17629
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 24489 17663 24547 17669
rect 24489 17660 24501 17663
rect 21821 17623 21879 17629
rect 22296 17632 24501 17660
rect 21450 17552 21456 17604
rect 21508 17592 21514 17604
rect 21846 17592 21874 17623
rect 21508 17564 21874 17592
rect 21508 17552 21514 17564
rect 22296 17524 22324 17632
rect 24489 17629 24501 17632
rect 24535 17660 24547 17663
rect 24854 17660 24860 17672
rect 24535 17632 24860 17660
rect 24535 17629 24547 17632
rect 24489 17623 24547 17629
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 26053 17663 26111 17669
rect 26053 17629 26065 17663
rect 26099 17660 26111 17663
rect 26142 17660 26148 17672
rect 26099 17632 26148 17660
rect 26099 17629 26111 17632
rect 26053 17623 26111 17629
rect 26142 17620 26148 17632
rect 26200 17620 26206 17672
rect 28184 17660 28212 17827
rect 30650 17824 30656 17876
rect 30708 17864 30714 17876
rect 32401 17867 32459 17873
rect 32401 17864 32413 17867
rect 30708 17836 32413 17864
rect 30708 17824 30714 17836
rect 32401 17833 32413 17836
rect 32447 17864 32459 17867
rect 36170 17864 36176 17876
rect 32447 17836 36176 17864
rect 32447 17833 32459 17836
rect 32401 17827 32459 17833
rect 36170 17824 36176 17836
rect 36228 17824 36234 17876
rect 36814 17824 36820 17876
rect 36872 17864 36878 17876
rect 37921 17867 37979 17873
rect 37921 17864 37933 17867
rect 36872 17836 37933 17864
rect 36872 17824 36878 17836
rect 37921 17833 37933 17836
rect 37967 17833 37979 17867
rect 37921 17827 37979 17833
rect 30466 17796 30472 17808
rect 30427 17768 30472 17796
rect 30466 17756 30472 17768
rect 30524 17756 30530 17808
rect 36078 17796 36084 17808
rect 36039 17768 36084 17796
rect 36078 17756 36084 17768
rect 36136 17756 36142 17808
rect 28813 17663 28871 17669
rect 28813 17660 28825 17663
rect 28184 17632 28825 17660
rect 28813 17629 28825 17632
rect 28859 17629 28871 17663
rect 28813 17623 28871 17629
rect 28997 17663 29055 17669
rect 28997 17629 29009 17663
rect 29043 17660 29055 17663
rect 30374 17660 30380 17672
rect 29043 17632 30380 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 30926 17620 30932 17672
rect 30984 17660 30990 17672
rect 31021 17663 31079 17669
rect 31021 17660 31033 17663
rect 30984 17632 31033 17660
rect 30984 17620 30990 17632
rect 31021 17629 31033 17632
rect 31067 17660 31079 17663
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 31067 17632 34713 17660
rect 31067 17629 31079 17632
rect 31021 17623 31079 17629
rect 34701 17629 34713 17632
rect 34747 17660 34759 17663
rect 36541 17663 36599 17669
rect 36541 17660 36553 17663
rect 34747 17632 36553 17660
rect 34747 17629 34759 17632
rect 34701 17623 34759 17629
rect 36541 17629 36553 17632
rect 36587 17629 36599 17663
rect 36541 17623 36599 17629
rect 26320 17595 26378 17601
rect 26320 17561 26332 17595
rect 26366 17592 26378 17595
rect 26418 17592 26424 17604
rect 26366 17564 26424 17592
rect 26366 17561 26378 17564
rect 26320 17555 26378 17561
rect 26418 17552 26424 17564
rect 26476 17552 26482 17604
rect 29638 17592 29644 17604
rect 26988 17564 29644 17592
rect 20548 17496 22324 17524
rect 22370 17484 22376 17536
rect 22428 17524 22434 17536
rect 22465 17527 22523 17533
rect 22465 17524 22477 17527
rect 22428 17496 22477 17524
rect 22428 17484 22434 17496
rect 22465 17493 22477 17496
rect 22511 17493 22523 17527
rect 25130 17524 25136 17536
rect 25091 17496 25136 17524
rect 22465 17487 22523 17493
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 25590 17484 25596 17536
rect 25648 17524 25654 17536
rect 26988 17524 27016 17564
rect 29638 17552 29644 17564
rect 29696 17552 29702 17604
rect 30098 17592 30104 17604
rect 30059 17564 30104 17592
rect 30098 17552 30104 17564
rect 30156 17552 30162 17604
rect 31110 17552 31116 17604
rect 31168 17592 31174 17604
rect 31266 17595 31324 17601
rect 31266 17592 31278 17595
rect 31168 17564 31278 17592
rect 31168 17552 31174 17564
rect 31266 17561 31278 17564
rect 31312 17561 31324 17595
rect 31266 17555 31324 17561
rect 31846 17552 31852 17604
rect 31904 17592 31910 17604
rect 32953 17595 33011 17601
rect 32953 17592 32965 17595
rect 31904 17564 32965 17592
rect 31904 17552 31910 17564
rect 32953 17561 32965 17564
rect 32999 17592 33011 17595
rect 33597 17595 33655 17601
rect 33597 17592 33609 17595
rect 32999 17564 33609 17592
rect 32999 17561 33011 17564
rect 32953 17555 33011 17561
rect 33597 17561 33609 17564
rect 33643 17561 33655 17595
rect 33597 17555 33655 17561
rect 33781 17595 33839 17601
rect 33781 17561 33793 17595
rect 33827 17592 33839 17595
rect 34422 17592 34428 17604
rect 33827 17564 34428 17592
rect 33827 17561 33839 17564
rect 33781 17555 33839 17561
rect 34422 17552 34428 17564
rect 34480 17552 34486 17604
rect 34790 17552 34796 17604
rect 34848 17592 34854 17604
rect 34946 17595 35004 17601
rect 34946 17592 34958 17595
rect 34848 17564 34958 17592
rect 34848 17552 34854 17564
rect 34946 17561 34958 17564
rect 34992 17561 35004 17595
rect 34946 17555 35004 17561
rect 35894 17552 35900 17604
rect 35952 17592 35958 17604
rect 36786 17595 36844 17601
rect 36786 17592 36798 17595
rect 35952 17564 36798 17592
rect 35952 17552 35958 17564
rect 36786 17561 36798 17564
rect 36832 17561 36844 17595
rect 36786 17555 36844 17561
rect 25648 17496 27016 17524
rect 25648 17484 25654 17496
rect 27062 17484 27068 17536
rect 27120 17524 27126 17536
rect 27433 17527 27491 17533
rect 27433 17524 27445 17527
rect 27120 17496 27445 17524
rect 27120 17484 27126 17496
rect 27433 17493 27445 17496
rect 27479 17493 27491 17527
rect 27433 17487 27491 17493
rect 30561 17527 30619 17533
rect 30561 17493 30573 17527
rect 30607 17524 30619 17527
rect 31570 17524 31576 17536
rect 30607 17496 31576 17524
rect 30607 17493 30619 17496
rect 30561 17487 30619 17493
rect 31570 17484 31576 17496
rect 31628 17484 31634 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 2130 17320 2136 17332
rect 2091 17292 2136 17320
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 3326 17320 3332 17332
rect 3239 17292 3332 17320
rect 3326 17280 3332 17292
rect 3384 17320 3390 17332
rect 3970 17320 3976 17332
rect 3384 17292 3976 17320
rect 3384 17280 3390 17292
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 12066 17320 12072 17332
rect 6604 17292 12072 17320
rect 6604 17280 6610 17292
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 13354 17320 13360 17332
rect 13315 17292 13360 17320
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 14461 17323 14519 17329
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 14550 17320 14556 17332
rect 14507 17292 14556 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 14550 17280 14556 17292
rect 14608 17320 14614 17332
rect 16574 17320 16580 17332
rect 14608 17292 16580 17320
rect 14608 17280 14614 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 18472 17292 19012 17320
rect 18472 17280 18478 17292
rect 12342 17252 12348 17264
rect 7024 17224 12348 17252
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 2777 17187 2835 17193
rect 2777 17184 2789 17187
rect 1719 17156 2789 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 2777 17153 2789 17156
rect 2823 17184 2835 17187
rect 4062 17184 4068 17196
rect 2823 17156 4068 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7024 17193 7052 17224
rect 12342 17212 12348 17224
rect 12400 17252 12406 17264
rect 18322 17252 18328 17264
rect 12400 17224 18328 17252
rect 12400 17212 12406 17224
rect 7009 17187 7067 17193
rect 7009 17184 7021 17187
rect 6972 17156 7021 17184
rect 6972 17144 6978 17156
rect 7009 17153 7021 17156
rect 7055 17153 7067 17187
rect 7009 17147 7067 17153
rect 8472 17187 8530 17193
rect 8472 17153 8484 17187
rect 8518 17184 8530 17187
rect 8938 17184 8944 17196
rect 8518 17156 8944 17184
rect 8518 17153 8530 17156
rect 8472 17147 8530 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11790 17184 11796 17196
rect 11112 17156 11796 17184
rect 11112 17144 11118 17156
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12584 17156 12633 17184
rect 12584 17144 12590 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12710 17144 12716 17196
rect 12768 17184 12774 17196
rect 13740 17193 13768 17224
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 18506 17252 18512 17264
rect 18467 17224 18512 17252
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 18782 17252 18788 17264
rect 18743 17224 18788 17252
rect 18782 17212 18788 17224
rect 18840 17212 18846 17264
rect 18984 17261 19012 17292
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 20346 17320 20352 17332
rect 19484 17292 20352 17320
rect 19484 17280 19490 17292
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 21818 17320 21824 17332
rect 20496 17292 21128 17320
rect 21779 17292 21824 17320
rect 20496 17280 20502 17292
rect 18984 17255 19053 17261
rect 18984 17224 19007 17255
rect 18995 17221 19007 17224
rect 19041 17221 19053 17255
rect 18995 17215 19053 17221
rect 19242 17212 19248 17264
rect 19300 17252 19306 17264
rect 20254 17252 20260 17264
rect 19300 17224 20260 17252
rect 19300 17212 19306 17224
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12768 17156 12817 17184
rect 12768 17144 12774 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17153 13783 17187
rect 13725 17147 13783 17153
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 14424 17156 17141 17184
rect 14424 17144 14430 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17153 18751 17187
rect 18693 17147 18751 17153
rect 18878 17187 18936 17193
rect 18878 17153 18890 17187
rect 18924 17174 18936 17187
rect 19889 17187 19947 17193
rect 19058 17174 19064 17186
rect 18924 17153 19064 17174
rect 18878 17147 19064 17153
rect 6822 17076 6828 17128
rect 6880 17116 6886 17128
rect 7156 17119 7214 17125
rect 7156 17116 7168 17119
rect 6880 17088 7168 17116
rect 6880 17076 6886 17088
rect 7156 17085 7168 17088
rect 7202 17085 7214 17119
rect 7374 17116 7380 17128
rect 7335 17088 7380 17116
rect 7156 17079 7214 17085
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8110 17076 8116 17128
rect 8168 17116 8174 17128
rect 8205 17119 8263 17125
rect 8205 17116 8217 17119
rect 8168 17088 8217 17116
rect 8168 17076 8174 17088
rect 8205 17085 8217 17088
rect 8251 17085 8263 17119
rect 10686 17116 10692 17128
rect 10647 17088 10692 17116
rect 8205 17079 8263 17085
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 13633 17119 13691 17125
rect 10796 17088 12434 17116
rect 9585 17051 9643 17057
rect 9585 17017 9597 17051
rect 9631 17048 9643 17051
rect 10042 17048 10048 17060
rect 9631 17020 10048 17048
rect 9631 17017 9643 17020
rect 9585 17011 9643 17017
rect 10042 17008 10048 17020
rect 10100 17048 10106 17060
rect 10796 17048 10824 17088
rect 10100 17020 10824 17048
rect 12406 17048 12434 17088
rect 12728 17088 13584 17116
rect 12728 17048 12756 17088
rect 12406 17020 12756 17048
rect 13556 17048 13584 17088
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 14918 17116 14924 17128
rect 13679 17088 14924 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 18708 17116 18736 17147
rect 18892 17146 19064 17147
rect 19058 17134 19064 17146
rect 19116 17134 19122 17186
rect 19889 17153 19901 17187
rect 19935 17184 19947 17187
rect 20898 17184 20904 17196
rect 19935 17156 20904 17184
rect 19935 17153 19947 17156
rect 19889 17147 19947 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 21100 17193 21128 17292
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 23293 17323 23351 17329
rect 23293 17320 23305 17323
rect 21928 17292 23305 17320
rect 21266 17212 21272 17264
rect 21324 17252 21330 17264
rect 21928 17252 21956 17292
rect 23293 17289 23305 17292
rect 23339 17289 23351 17323
rect 23293 17283 23351 17289
rect 23753 17323 23811 17329
rect 23753 17289 23765 17323
rect 23799 17320 23811 17323
rect 26970 17320 26976 17332
rect 23799 17292 26976 17320
rect 23799 17289 23811 17292
rect 23753 17283 23811 17289
rect 21324 17224 21956 17252
rect 21324 17212 21330 17224
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 21450 17144 21456 17196
rect 21508 17184 21514 17196
rect 21818 17184 21824 17196
rect 21508 17156 21824 17184
rect 21508 17144 21514 17156
rect 21818 17144 21824 17156
rect 21876 17184 21882 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21876 17156 22017 17184
rect 21876 17144 21882 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22278 17184 22284 17196
rect 22239 17156 22284 17184
rect 22005 17147 22063 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 22646 17144 22652 17196
rect 22704 17184 22710 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22704 17156 22845 17184
rect 22704 17144 22710 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 23014 17184 23020 17196
rect 22975 17156 23020 17184
rect 22833 17147 22891 17153
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 23109 17187 23167 17193
rect 23109 17153 23121 17187
rect 23155 17184 23167 17187
rect 23768 17184 23796 17283
rect 26970 17280 26976 17292
rect 27028 17280 27034 17332
rect 30193 17323 30251 17329
rect 30193 17289 30205 17323
rect 30239 17320 30251 17323
rect 30282 17320 30288 17332
rect 30239 17292 30288 17320
rect 30239 17289 30251 17292
rect 30193 17283 30251 17289
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 33689 17323 33747 17329
rect 33689 17289 33701 17323
rect 33735 17320 33747 17323
rect 34514 17320 34520 17332
rect 33735 17292 34520 17320
rect 33735 17289 33747 17292
rect 33689 17283 33747 17289
rect 34514 17280 34520 17292
rect 34572 17280 34578 17332
rect 35342 17320 35348 17332
rect 35303 17292 35348 17320
rect 35342 17280 35348 17292
rect 35400 17280 35406 17332
rect 25777 17255 25835 17261
rect 25777 17221 25789 17255
rect 25823 17252 25835 17255
rect 30650 17252 30656 17264
rect 25823 17224 30656 17252
rect 25823 17221 25835 17224
rect 25777 17215 25835 17221
rect 30650 17212 30656 17224
rect 30708 17212 30714 17264
rect 30742 17212 30748 17264
rect 30800 17252 30806 17264
rect 33962 17252 33968 17264
rect 30800 17224 33968 17252
rect 30800 17212 30806 17224
rect 33962 17212 33968 17224
rect 34020 17252 34026 17264
rect 34609 17255 34667 17261
rect 34020 17224 34560 17252
rect 34020 17212 34026 17224
rect 24854 17184 24860 17196
rect 23155 17156 23796 17184
rect 24815 17156 24860 17184
rect 23155 17153 23167 17156
rect 23109 17147 23167 17153
rect 24854 17144 24860 17156
rect 24912 17144 24918 17196
rect 25590 17184 25596 17196
rect 25056 17156 25596 17184
rect 19153 17119 19211 17125
rect 18708 17088 18920 17116
rect 17313 17051 17371 17057
rect 13556 17020 15884 17048
rect 10100 17008 10106 17020
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 7340 16952 7385 16980
rect 7340 16940 7346 16952
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13538 16980 13544 16992
rect 12952 16952 12997 16980
rect 13499 16952 13544 16980
rect 12952 16940 12958 16952
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 15856 16989 15884 17020
rect 17313 17017 17325 17051
rect 17359 17048 17371 17051
rect 17494 17048 17500 17060
rect 17359 17020 17500 17048
rect 17359 17017 17371 17020
rect 17313 17011 17371 17017
rect 17494 17008 17500 17020
rect 17552 17008 17558 17060
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 16114 16980 16120 16992
rect 15887 16952 16120 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 18892 16980 18920 17088
rect 19153 17085 19165 17119
rect 19199 17116 19211 17119
rect 19242 17116 19248 17128
rect 19199 17088 19248 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 19613 17119 19671 17125
rect 19613 17085 19625 17119
rect 19659 17085 19671 17119
rect 25056 17116 25084 17156
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 25958 17184 25964 17196
rect 25919 17156 25964 17184
rect 25958 17144 25964 17156
rect 26016 17144 26022 17196
rect 27706 17184 27712 17196
rect 27667 17156 27712 17184
rect 27706 17144 27712 17156
rect 27764 17144 27770 17196
rect 29638 17144 29644 17196
rect 29696 17184 29702 17196
rect 30561 17187 30619 17193
rect 30561 17184 30573 17187
rect 29696 17156 30573 17184
rect 29696 17144 29702 17156
rect 30561 17153 30573 17156
rect 30607 17184 30619 17187
rect 31570 17184 31576 17196
rect 30607 17156 30880 17184
rect 31531 17156 31576 17184
rect 30607 17153 30619 17156
rect 30561 17147 30619 17153
rect 19613 17079 19671 17085
rect 20732 17088 25084 17116
rect 18966 17008 18972 17060
rect 19024 17048 19030 17060
rect 19628 17048 19656 17079
rect 19024 17020 19656 17048
rect 19024 17008 19030 17020
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 20438 17048 20444 17060
rect 19760 17020 20444 17048
rect 19760 17008 19766 17020
rect 20438 17008 20444 17020
rect 20496 17048 20502 17060
rect 20732 17048 20760 17088
rect 25130 17076 25136 17128
rect 25188 17116 25194 17128
rect 25188 17088 25233 17116
rect 25188 17076 25194 17088
rect 27338 17076 27344 17128
rect 27396 17116 27402 17128
rect 27433 17119 27491 17125
rect 27433 17116 27445 17119
rect 27396 17088 27445 17116
rect 27396 17076 27402 17088
rect 27433 17085 27445 17088
rect 27479 17116 27491 17119
rect 27982 17116 27988 17128
rect 27479 17088 27988 17116
rect 27479 17085 27491 17088
rect 27433 17079 27491 17085
rect 27982 17076 27988 17088
rect 28040 17116 28046 17128
rect 28353 17119 28411 17125
rect 28353 17116 28365 17119
rect 28040 17088 28365 17116
rect 28040 17076 28046 17088
rect 28353 17085 28365 17088
rect 28399 17085 28411 17119
rect 28353 17079 28411 17085
rect 30374 17076 30380 17128
rect 30432 17116 30438 17128
rect 30745 17119 30803 17125
rect 30745 17116 30757 17119
rect 30432 17088 30757 17116
rect 30432 17076 30438 17088
rect 30745 17085 30757 17088
rect 30791 17085 30803 17119
rect 30852 17116 30880 17156
rect 31570 17144 31576 17156
rect 31628 17144 31634 17196
rect 34532 17193 34560 17224
rect 34609 17221 34621 17255
rect 34655 17252 34667 17255
rect 36078 17252 36084 17264
rect 34655 17224 36084 17252
rect 34655 17221 34667 17224
rect 34609 17215 34667 17221
rect 36078 17212 36084 17224
rect 36136 17252 36142 17264
rect 37090 17252 37096 17264
rect 36136 17224 37096 17252
rect 36136 17212 36142 17224
rect 37090 17212 37096 17224
rect 37148 17212 37154 17264
rect 37921 17255 37979 17261
rect 37921 17221 37933 17255
rect 37967 17252 37979 17255
rect 38286 17252 38292 17264
rect 37967 17224 38292 17252
rect 37967 17221 37979 17224
rect 37921 17215 37979 17221
rect 38286 17212 38292 17224
rect 38344 17212 38350 17264
rect 34517 17187 34575 17193
rect 34517 17153 34529 17187
rect 34563 17153 34575 17187
rect 34517 17147 34575 17153
rect 36449 17187 36507 17193
rect 36449 17153 36461 17187
rect 36495 17184 36507 17187
rect 37182 17184 37188 17196
rect 36495 17156 37188 17184
rect 36495 17153 36507 17156
rect 36449 17147 36507 17153
rect 37182 17144 37188 17156
rect 37240 17144 37246 17196
rect 37274 17144 37280 17196
rect 37332 17184 37338 17196
rect 37737 17187 37795 17193
rect 37737 17184 37749 17187
rect 37332 17156 37749 17184
rect 37332 17144 37338 17156
rect 37737 17153 37749 17156
rect 37783 17153 37795 17187
rect 37737 17147 37795 17153
rect 33134 17116 33140 17128
rect 30852 17088 33140 17116
rect 30745 17079 30803 17085
rect 33134 17076 33140 17088
rect 33192 17076 33198 17128
rect 33226 17076 33232 17128
rect 33284 17116 33290 17128
rect 34701 17119 34759 17125
rect 33284 17088 33329 17116
rect 33284 17076 33290 17088
rect 34701 17085 34713 17119
rect 34747 17085 34759 17119
rect 34701 17079 34759 17085
rect 20990 17048 20996 17060
rect 20496 17020 20760 17048
rect 20824 17020 20996 17048
rect 20496 17008 20502 17020
rect 20824 16980 20852 17020
rect 20990 17008 20996 17020
rect 21048 17008 21054 17060
rect 21910 17008 21916 17060
rect 21968 17048 21974 17060
rect 22097 17051 22155 17057
rect 22097 17048 22109 17051
rect 21968 17020 22109 17048
rect 21968 17008 21974 17020
rect 22097 17017 22109 17020
rect 22143 17017 22155 17051
rect 22097 17011 22155 17017
rect 22189 17051 22247 17057
rect 22189 17017 22201 17051
rect 22235 17048 22247 17051
rect 22370 17048 22376 17060
rect 22235 17020 22376 17048
rect 22235 17017 22247 17020
rect 22189 17011 22247 17017
rect 22370 17008 22376 17020
rect 22428 17008 22434 17060
rect 22462 17008 22468 17060
rect 22520 17048 22526 17060
rect 23014 17048 23020 17060
rect 22520 17020 23020 17048
rect 22520 17008 22526 17020
rect 23014 17008 23020 17020
rect 23072 17008 23078 17060
rect 23658 17008 23664 17060
rect 23716 17048 23722 17060
rect 25593 17051 25651 17057
rect 25593 17048 25605 17051
rect 23716 17020 25605 17048
rect 23716 17008 23722 17020
rect 25593 17017 25605 17020
rect 25639 17017 25651 17051
rect 28534 17048 28540 17060
rect 25593 17011 25651 17017
rect 27540 17020 28540 17048
rect 18892 16952 20852 16980
rect 20901 16983 20959 16989
rect 20901 16949 20913 16983
rect 20947 16980 20959 16983
rect 21082 16980 21088 16992
rect 20947 16952 21088 16980
rect 20947 16949 20959 16952
rect 20901 16943 20959 16949
rect 21082 16940 21088 16952
rect 21140 16980 21146 16992
rect 21726 16980 21732 16992
rect 21140 16952 21732 16980
rect 21140 16940 21146 16952
rect 21726 16940 21732 16952
rect 21784 16980 21790 16992
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 21784 16952 22845 16980
rect 21784 16940 21790 16952
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 24673 16983 24731 16989
rect 24673 16949 24685 16983
rect 24719 16980 24731 16983
rect 24762 16980 24768 16992
rect 24719 16952 24768 16980
rect 24719 16949 24731 16952
rect 24673 16943 24731 16949
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 24946 16940 24952 16992
rect 25004 16980 25010 16992
rect 25041 16983 25099 16989
rect 25041 16980 25053 16983
rect 25004 16952 25053 16980
rect 25004 16940 25010 16952
rect 25041 16949 25053 16952
rect 25087 16980 25099 16983
rect 25222 16980 25228 16992
rect 25087 16952 25228 16980
rect 25087 16949 25099 16952
rect 25041 16943 25099 16949
rect 25222 16940 25228 16952
rect 25280 16980 25286 16992
rect 27540 16989 27568 17020
rect 28534 17008 28540 17020
rect 28592 17048 28598 17060
rect 28997 17051 29055 17057
rect 28997 17048 29009 17051
rect 28592 17020 29009 17048
rect 28592 17008 28598 17020
rect 28997 17017 29009 17020
rect 29043 17017 29055 17051
rect 28997 17011 29055 17017
rect 33597 17051 33655 17057
rect 33597 17017 33609 17051
rect 33643 17048 33655 17051
rect 34149 17051 34207 17057
rect 34149 17048 34161 17051
rect 33643 17020 34161 17048
rect 33643 17017 33655 17020
rect 33597 17011 33655 17017
rect 34149 17017 34161 17020
rect 34195 17017 34207 17051
rect 34149 17011 34207 17017
rect 34422 17008 34428 17060
rect 34480 17048 34486 17060
rect 34716 17048 34744 17079
rect 35342 17076 35348 17128
rect 35400 17116 35406 17128
rect 36354 17116 36360 17128
rect 35400 17088 36360 17116
rect 35400 17076 35406 17088
rect 36354 17076 36360 17088
rect 36412 17116 36418 17128
rect 36725 17119 36783 17125
rect 36725 17116 36737 17119
rect 36412 17088 36737 17116
rect 36412 17076 36418 17088
rect 36725 17085 36737 17088
rect 36771 17085 36783 17119
rect 36725 17079 36783 17085
rect 34480 17020 34744 17048
rect 34480 17008 34486 17020
rect 27525 16983 27583 16989
rect 27525 16980 27537 16983
rect 25280 16952 27537 16980
rect 25280 16940 25286 16952
rect 27525 16949 27537 16952
rect 27571 16949 27583 16983
rect 27525 16943 27583 16949
rect 27798 16940 27804 16992
rect 27856 16980 27862 16992
rect 27893 16983 27951 16989
rect 27893 16980 27905 16983
rect 27856 16952 27905 16980
rect 27856 16940 27862 16952
rect 27893 16949 27905 16952
rect 27939 16949 27951 16983
rect 27893 16943 27951 16949
rect 29641 16983 29699 16989
rect 29641 16949 29653 16983
rect 29687 16980 29699 16983
rect 29730 16980 29736 16992
rect 29687 16952 29736 16980
rect 29687 16949 29699 16952
rect 29641 16943 29699 16949
rect 29730 16940 29736 16952
rect 29788 16980 29794 16992
rect 30742 16980 30748 16992
rect 29788 16952 30748 16980
rect 29788 16940 29794 16952
rect 30742 16940 30748 16952
rect 30800 16940 30806 16992
rect 31202 16940 31208 16992
rect 31260 16980 31266 16992
rect 31389 16983 31447 16989
rect 31389 16980 31401 16983
rect 31260 16952 31401 16980
rect 31260 16940 31266 16952
rect 31389 16949 31401 16952
rect 31435 16949 31447 16983
rect 31389 16943 31447 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2133 16779 2191 16785
rect 2133 16745 2145 16779
rect 2179 16776 2191 16779
rect 6270 16776 6276 16788
rect 2179 16748 6276 16776
rect 2179 16745 2191 16748
rect 2133 16739 2191 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6438 16779 6496 16785
rect 6438 16745 6450 16779
rect 6484 16776 6496 16779
rect 6822 16776 6828 16788
rect 6484 16748 6828 16776
rect 6484 16745 6496 16748
rect 6438 16739 6496 16745
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 16206 16776 16212 16788
rect 13136 16748 16068 16776
rect 16167 16748 16212 16776
rect 13136 16736 13142 16748
rect 6546 16708 6552 16720
rect 6507 16680 6552 16708
rect 6546 16668 6552 16680
rect 6604 16668 6610 16720
rect 12434 16708 12440 16720
rect 12360 16680 12440 16708
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 7374 16640 7380 16652
rect 6687 16612 7380 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 9508 16612 10977 16640
rect 9508 16584 9536 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 12250 16640 12256 16652
rect 11287 16612 12256 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 12360 16649 12388 16680
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 13354 16668 13360 16720
rect 13412 16708 13418 16720
rect 15930 16708 15936 16720
rect 13412 16680 15936 16708
rect 13412 16668 13418 16680
rect 15930 16668 15936 16680
rect 15988 16668 15994 16720
rect 16040 16708 16068 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 17681 16779 17739 16785
rect 17681 16745 17693 16779
rect 17727 16776 17739 16779
rect 19242 16776 19248 16788
rect 17727 16748 19248 16776
rect 17727 16745 17739 16748
rect 17681 16739 17739 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 22189 16779 22247 16785
rect 21836 16748 22094 16776
rect 19702 16708 19708 16720
rect 16040 16680 19708 16708
rect 19702 16668 19708 16680
rect 19760 16668 19766 16720
rect 21836 16717 21864 16748
rect 21821 16711 21879 16717
rect 21821 16677 21833 16711
rect 21867 16677 21879 16711
rect 22066 16708 22094 16748
rect 22189 16745 22201 16779
rect 22235 16776 22247 16779
rect 22830 16776 22836 16788
rect 22235 16748 22836 16776
rect 22235 16745 22247 16748
rect 22189 16739 22247 16745
rect 22830 16736 22836 16748
rect 22888 16736 22894 16788
rect 26234 16776 26240 16788
rect 24504 16748 26240 16776
rect 22370 16708 22376 16720
rect 22066 16680 22376 16708
rect 21821 16671 21879 16677
rect 22370 16668 22376 16680
rect 22428 16668 22434 16720
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 13320 16612 14565 16640
rect 13320 16600 13326 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 14875 16612 15976 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 7926 16572 7932 16584
rect 7887 16544 7932 16572
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16572 8263 16575
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8251 16544 8953 16572
rect 8251 16541 8263 16544
rect 8205 16535 8263 16541
rect 8941 16541 8953 16544
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16572 9459 16575
rect 9490 16572 9496 16584
rect 9447 16544 9496 16572
rect 9447 16541 9459 16544
rect 9401 16535 9459 16541
rect 1854 16504 1860 16516
rect 1815 16476 1860 16504
rect 1854 16464 1860 16476
rect 1912 16504 1918 16516
rect 2685 16507 2743 16513
rect 2685 16504 2697 16507
rect 1912 16476 2697 16504
rect 1912 16464 1918 16476
rect 2685 16473 2697 16476
rect 2731 16473 2743 16507
rect 6270 16504 6276 16516
rect 6231 16476 6276 16504
rect 2685 16467 2743 16473
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 7006 16504 7012 16516
rect 6967 16476 7012 16504
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 8036 16504 8064 16535
rect 9140 16504 9168 16535
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 9950 16572 9956 16584
rect 9631 16544 9956 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 10836 16544 12449 16572
rect 10836 16532 10842 16544
rect 12437 16541 12449 16544
rect 12483 16572 12495 16575
rect 12526 16572 12532 16584
rect 12483 16544 12532 16572
rect 12483 16541 12495 16544
rect 12437 16535 12495 16541
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 12986 16572 12992 16584
rect 12947 16544 12992 16572
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 15948 16572 15976 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 16080 16612 16313 16640
rect 16080 16600 16086 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 17000 16612 17325 16640
rect 17000 16600 17006 16612
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 18230 16640 18236 16652
rect 17451 16612 18236 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16640 19855 16643
rect 20254 16640 20260 16652
rect 19843 16612 20260 16640
rect 19843 16609 19855 16612
rect 19797 16603 19855 16609
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 20772 16612 20821 16640
rect 20772 16600 20778 16612
rect 20809 16609 20821 16612
rect 20855 16640 20867 16643
rect 23290 16640 23296 16652
rect 20855 16612 23296 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 23290 16600 23296 16612
rect 23348 16600 23354 16652
rect 24504 16649 24532 16748
rect 26234 16736 26240 16748
rect 26292 16736 26298 16788
rect 30466 16776 30472 16788
rect 30427 16748 30472 16776
rect 30466 16736 30472 16748
rect 30524 16736 30530 16788
rect 32769 16779 32827 16785
rect 32769 16776 32781 16779
rect 30944 16748 32781 16776
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16609 24547 16643
rect 26252 16640 26280 16736
rect 29656 16680 30512 16708
rect 27525 16643 27583 16649
rect 27525 16640 27537 16643
rect 26252 16612 27537 16640
rect 24489 16603 24547 16609
rect 27525 16609 27537 16612
rect 27571 16609 27583 16643
rect 27525 16603 27583 16609
rect 16209 16575 16267 16581
rect 16209 16572 16221 16575
rect 15948 16544 16221 16572
rect 16209 16541 16221 16544
rect 16255 16572 16267 16575
rect 16390 16572 16396 16584
rect 16255 16544 16396 16572
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 10318 16504 10324 16516
rect 8036 16476 8524 16504
rect 9140 16476 10324 16504
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8389 16439 8447 16445
rect 8389 16436 8401 16439
rect 8352 16408 8401 16436
rect 8352 16396 8358 16408
rect 8389 16405 8401 16408
rect 8435 16405 8447 16439
rect 8496 16436 8524 16476
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 16298 16464 16304 16516
rect 16356 16504 16362 16516
rect 16500 16504 16528 16535
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 17221 16575 17279 16581
rect 17221 16572 17233 16575
rect 16724 16544 17233 16572
rect 16724 16532 16730 16544
rect 17221 16541 17233 16544
rect 17267 16541 17279 16575
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 17221 16535 17279 16541
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 20073 16575 20131 16581
rect 20073 16572 20085 16575
rect 17644 16544 20085 16572
rect 17644 16532 17650 16544
rect 20073 16541 20085 16544
rect 20119 16572 20131 16575
rect 21726 16572 21732 16584
rect 20119 16544 20668 16572
rect 21687 16544 21732 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20640 16513 20668 16544
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 21910 16572 21916 16584
rect 21871 16544 21916 16572
rect 21910 16532 21916 16544
rect 21968 16532 21974 16584
rect 24762 16581 24768 16584
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16541 22063 16575
rect 24756 16572 24768 16581
rect 24723 16544 24768 16572
rect 22005 16535 22063 16541
rect 24756 16535 24768 16544
rect 16356 16476 16528 16504
rect 20625 16507 20683 16513
rect 16356 16464 16362 16476
rect 20625 16473 20637 16507
rect 20671 16473 20683 16507
rect 20625 16467 20683 16473
rect 21818 16464 21824 16516
rect 21876 16504 21882 16516
rect 22020 16504 22048 16535
rect 24762 16532 24768 16535
rect 24820 16532 24826 16584
rect 26605 16575 26663 16581
rect 26605 16541 26617 16575
rect 26651 16541 26663 16575
rect 26878 16572 26884 16584
rect 26839 16544 26884 16572
rect 26605 16535 26663 16541
rect 24946 16504 24952 16516
rect 21876 16476 22048 16504
rect 22112 16476 24952 16504
rect 21876 16464 21882 16476
rect 10686 16436 10692 16448
rect 8496 16408 10692 16436
rect 8389 16399 8447 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 12345 16439 12403 16445
rect 12345 16405 12357 16439
rect 12391 16436 12403 16439
rect 12802 16436 12808 16448
rect 12391 16408 12808 16436
rect 12391 16405 12403 16408
rect 12345 16399 12403 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18601 16439 18659 16445
rect 18601 16436 18613 16439
rect 18196 16408 18613 16436
rect 18196 16396 18202 16408
rect 18601 16405 18613 16408
rect 18647 16405 18659 16439
rect 18601 16399 18659 16405
rect 18782 16396 18788 16448
rect 18840 16436 18846 16448
rect 22112 16436 22140 16476
rect 24946 16464 24952 16476
rect 25004 16504 25010 16516
rect 26620 16504 26648 16535
rect 26878 16532 26884 16544
rect 26936 16532 26942 16584
rect 27062 16572 27068 16584
rect 27023 16544 27068 16572
rect 27062 16532 27068 16544
rect 27120 16532 27126 16584
rect 27798 16581 27804 16584
rect 27792 16572 27804 16581
rect 27759 16544 27804 16572
rect 27792 16535 27804 16544
rect 27798 16532 27804 16535
rect 27856 16532 27862 16584
rect 27430 16504 27436 16516
rect 25004 16476 27436 16504
rect 25004 16464 25010 16476
rect 27430 16464 27436 16476
rect 27488 16464 27494 16516
rect 18840 16408 22140 16436
rect 18840 16396 18846 16408
rect 22370 16396 22376 16448
rect 22428 16436 22434 16448
rect 22649 16439 22707 16445
rect 22649 16436 22661 16439
rect 22428 16408 22661 16436
rect 22428 16396 22434 16408
rect 22649 16405 22661 16408
rect 22695 16405 22707 16439
rect 23290 16436 23296 16448
rect 23251 16408 23296 16436
rect 22649 16399 22707 16405
rect 23290 16396 23296 16408
rect 23348 16396 23354 16448
rect 25406 16396 25412 16448
rect 25464 16436 25470 16448
rect 25869 16439 25927 16445
rect 25869 16436 25881 16439
rect 25464 16408 25881 16436
rect 25464 16396 25470 16408
rect 25869 16405 25881 16408
rect 25915 16405 25927 16439
rect 25869 16399 25927 16405
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 26421 16439 26479 16445
rect 26421 16436 26433 16439
rect 26292 16408 26433 16436
rect 26292 16396 26298 16408
rect 26421 16405 26433 16408
rect 26467 16405 26479 16439
rect 26421 16399 26479 16405
rect 28166 16396 28172 16448
rect 28224 16436 28230 16448
rect 28905 16439 28963 16445
rect 28905 16436 28917 16439
rect 28224 16408 28917 16436
rect 28224 16396 28230 16408
rect 28905 16405 28917 16408
rect 28951 16436 28963 16439
rect 29656 16436 29684 16680
rect 29917 16643 29975 16649
rect 29917 16609 29929 16643
rect 29963 16640 29975 16643
rect 30374 16640 30380 16652
rect 29963 16612 30380 16640
rect 29963 16609 29975 16612
rect 29917 16603 29975 16609
rect 30374 16600 30380 16612
rect 30432 16600 30438 16652
rect 29730 16532 29736 16584
rect 29788 16572 29794 16584
rect 30101 16575 30159 16581
rect 30101 16572 30113 16575
rect 29788 16544 30113 16572
rect 29788 16532 29794 16544
rect 30101 16541 30113 16544
rect 30147 16541 30159 16575
rect 30101 16535 30159 16541
rect 30484 16504 30512 16680
rect 30944 16649 30972 16748
rect 32769 16745 32781 16748
rect 32815 16776 32827 16779
rect 34054 16776 34060 16788
rect 32815 16748 34060 16776
rect 32815 16745 32827 16748
rect 32769 16739 32827 16745
rect 34054 16736 34060 16748
rect 34112 16736 34118 16788
rect 32306 16708 32312 16720
rect 32267 16680 32312 16708
rect 32306 16668 32312 16680
rect 32364 16668 32370 16720
rect 33134 16668 33140 16720
rect 33192 16708 33198 16720
rect 33413 16711 33471 16717
rect 33413 16708 33425 16711
rect 33192 16680 33425 16708
rect 33192 16668 33198 16680
rect 33413 16677 33425 16680
rect 33459 16677 33471 16711
rect 33962 16708 33968 16720
rect 33923 16680 33968 16708
rect 33413 16671 33471 16677
rect 30929 16643 30987 16649
rect 30929 16609 30941 16643
rect 30975 16609 30987 16643
rect 33428 16640 33456 16671
rect 33962 16668 33968 16680
rect 34020 16668 34026 16720
rect 34422 16668 34428 16720
rect 34480 16708 34486 16720
rect 34480 16680 35296 16708
rect 34480 16668 34486 16680
rect 35268 16649 35296 16680
rect 35161 16643 35219 16649
rect 33428 16612 35112 16640
rect 30929 16603 30987 16609
rect 31202 16581 31208 16584
rect 31196 16572 31208 16581
rect 31163 16544 31208 16572
rect 31196 16535 31208 16544
rect 31202 16532 31208 16535
rect 31260 16532 31266 16584
rect 35084 16581 35112 16612
rect 35161 16609 35173 16643
rect 35207 16609 35219 16643
rect 35161 16603 35219 16609
rect 35253 16643 35311 16649
rect 35253 16609 35265 16643
rect 35299 16609 35311 16643
rect 35253 16603 35311 16609
rect 35360 16612 36860 16640
rect 35069 16575 35127 16581
rect 35069 16541 35081 16575
rect 35115 16541 35127 16575
rect 35176 16572 35204 16603
rect 35360 16572 35388 16612
rect 36832 16584 36860 16612
rect 35176 16544 35388 16572
rect 35989 16575 36047 16581
rect 35069 16535 35127 16541
rect 35989 16541 36001 16575
rect 36035 16572 36047 16575
rect 36078 16572 36084 16584
rect 36035 16544 36084 16572
rect 36035 16541 36047 16544
rect 35989 16535 36047 16541
rect 36078 16532 36084 16544
rect 36136 16532 36142 16584
rect 36814 16532 36820 16584
rect 36872 16532 36878 16584
rect 36998 16581 37004 16584
rect 36996 16572 37004 16581
rect 36959 16544 37004 16572
rect 36996 16535 37004 16544
rect 36998 16532 37004 16535
rect 37056 16532 37062 16584
rect 37182 16572 37188 16584
rect 37143 16544 37188 16572
rect 37182 16532 37188 16544
rect 37240 16532 37246 16584
rect 37366 16572 37372 16584
rect 37327 16544 37372 16572
rect 37366 16532 37372 16544
rect 37424 16532 37430 16584
rect 37458 16532 37464 16584
rect 37516 16572 37522 16584
rect 37516 16544 37561 16572
rect 37516 16532 37522 16544
rect 37642 16532 37648 16584
rect 37700 16572 37706 16584
rect 38102 16572 38108 16584
rect 37700 16544 38108 16572
rect 37700 16532 37706 16544
rect 38102 16532 38108 16544
rect 38160 16532 38166 16584
rect 32214 16504 32220 16516
rect 30024 16476 30236 16504
rect 30484 16476 32220 16504
rect 30024 16448 30052 16476
rect 30006 16436 30012 16448
rect 28951 16408 29684 16436
rect 29967 16408 30012 16436
rect 28951 16405 28963 16408
rect 28905 16399 28963 16405
rect 30006 16396 30012 16408
rect 30064 16396 30070 16448
rect 30208 16436 30236 16476
rect 32214 16464 32220 16476
rect 32272 16464 32278 16516
rect 36832 16504 36860 16532
rect 37093 16507 37151 16513
rect 37093 16504 37105 16507
rect 36832 16476 37105 16504
rect 37093 16473 37105 16476
rect 37139 16473 37151 16507
rect 37093 16467 37151 16473
rect 32306 16436 32312 16448
rect 30208 16408 32312 16436
rect 32306 16396 32312 16408
rect 32364 16396 32370 16448
rect 34701 16439 34759 16445
rect 34701 16405 34713 16439
rect 34747 16436 34759 16439
rect 34790 16436 34796 16448
rect 34747 16408 34796 16436
rect 34747 16405 34759 16408
rect 34701 16399 34759 16405
rect 34790 16396 34796 16408
rect 34848 16396 34854 16448
rect 36170 16436 36176 16448
rect 36131 16408 36176 16436
rect 36170 16396 36176 16408
rect 36228 16396 36234 16448
rect 36814 16436 36820 16448
rect 36775 16408 36820 16436
rect 36814 16396 36820 16408
rect 36872 16396 36878 16448
rect 37366 16396 37372 16448
rect 37424 16436 37430 16448
rect 37921 16439 37979 16445
rect 37921 16436 37933 16439
rect 37424 16408 37933 16436
rect 37424 16396 37430 16408
rect 37921 16405 37933 16408
rect 37967 16405 37979 16439
rect 37921 16399 37979 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 6914 16232 6920 16244
rect 6875 16204 6920 16232
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 13906 16232 13912 16244
rect 12406 16204 13912 16232
rect 8110 16164 8116 16176
rect 8023 16136 8116 16164
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2130 16096 2136 16108
rect 2091 16068 2136 16096
rect 2130 16056 2136 16068
rect 2188 16096 2194 16108
rect 2777 16099 2835 16105
rect 2777 16096 2789 16099
rect 2188 16068 2789 16096
rect 2188 16056 2194 16068
rect 2777 16065 2789 16068
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 6270 16056 6276 16108
rect 6328 16096 6334 16108
rect 8036 16105 8064 16136
rect 8110 16124 8116 16136
rect 8168 16164 8174 16176
rect 12406 16164 12434 16204
rect 13906 16192 13912 16204
rect 13964 16232 13970 16244
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 13964 16204 15117 16232
rect 13964 16192 13970 16204
rect 15105 16201 15117 16204
rect 15151 16201 15163 16235
rect 15105 16195 15163 16201
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 18966 16232 18972 16244
rect 16816 16204 18972 16232
rect 16816 16192 16822 16204
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 21634 16192 21640 16244
rect 21692 16232 21698 16244
rect 21821 16235 21879 16241
rect 21821 16232 21833 16235
rect 21692 16204 21833 16232
rect 21692 16192 21698 16204
rect 21821 16201 21833 16204
rect 21867 16201 21879 16235
rect 21821 16195 21879 16201
rect 22830 16192 22836 16244
rect 22888 16232 22894 16244
rect 23293 16235 23351 16241
rect 23293 16232 23305 16235
rect 22888 16204 23305 16232
rect 22888 16192 22894 16204
rect 23293 16201 23305 16204
rect 23339 16201 23351 16235
rect 23293 16195 23351 16201
rect 24765 16235 24823 16241
rect 24765 16201 24777 16235
rect 24811 16232 24823 16235
rect 24854 16232 24860 16244
rect 24811 16204 24860 16232
rect 24811 16201 24823 16204
rect 24765 16195 24823 16201
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 26418 16232 26424 16244
rect 26379 16204 26424 16232
rect 26418 16192 26424 16204
rect 26476 16192 26482 16244
rect 27617 16235 27675 16241
rect 27617 16201 27629 16235
rect 27663 16232 27675 16235
rect 27706 16232 27712 16244
rect 27663 16204 27712 16232
rect 27663 16201 27675 16204
rect 27617 16195 27675 16201
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 28166 16232 28172 16244
rect 28127 16204 28172 16232
rect 28166 16192 28172 16204
rect 28224 16192 28230 16244
rect 14366 16164 14372 16176
rect 8168 16136 12434 16164
rect 14327 16136 14372 16164
rect 8168 16124 8174 16136
rect 14366 16124 14372 16136
rect 14424 16124 14430 16176
rect 21542 16164 21548 16176
rect 15028 16136 21548 16164
rect 8294 16105 8300 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6328 16068 6837 16096
rect 6328 16056 6334 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16065 8079 16099
rect 8288 16096 8300 16105
rect 8255 16068 8300 16096
rect 8021 16059 8079 16065
rect 8288 16059 8300 16068
rect 8294 16056 8300 16059
rect 8352 16056 8358 16108
rect 10778 16096 10784 16108
rect 10739 16068 10784 16096
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 12250 16096 12256 16108
rect 12211 16068 12256 16096
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13538 16096 13544 16108
rect 13219 16068 13544 16096
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 13538 16056 13544 16068
rect 13596 16096 13602 16108
rect 15028 16096 15056 16136
rect 21542 16124 21548 16136
rect 21600 16164 21606 16176
rect 22646 16164 22652 16176
rect 21600 16136 22652 16164
rect 21600 16124 21606 16136
rect 22646 16124 22652 16136
rect 22704 16124 22710 16176
rect 28184 16164 28212 16192
rect 29454 16164 29460 16176
rect 25240 16136 25544 16164
rect 15194 16096 15200 16108
rect 13596 16068 15056 16096
rect 15155 16068 15200 16096
rect 13596 16056 13602 16068
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15930 16096 15936 16108
rect 15891 16068 15936 16096
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 17586 16096 17592 16108
rect 16040 16068 17592 16096
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 6972 16000 7481 16028
rect 6972 15988 6978 16000
rect 7469 15997 7481 16000
rect 7515 16028 7527 16031
rect 7926 16028 7932 16040
rect 7515 16000 7932 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12492 16000 12909 16028
rect 12492 15988 12498 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 16040 16028 16068 16068
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 18138 16056 18144 16108
rect 18196 16096 18202 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18196 16068 19073 16096
rect 18196 16056 18202 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 21450 16096 21456 16108
rect 21315 16068 21456 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 21818 16056 21824 16108
rect 21876 16096 21882 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21876 16068 22017 16096
rect 21876 16056 21882 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22462 16096 22468 16108
rect 22327 16068 22468 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 22664 16096 22692 16124
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22664 16068 22845 16096
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 24946 16096 24952 16108
rect 23155 16068 23888 16096
rect 24907 16068 24952 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 16758 16028 16764 16040
rect 12897 15991 12955 15997
rect 13004 16000 16068 16028
rect 16719 16000 16764 16028
rect 11882 15920 11888 15972
rect 11940 15960 11946 15972
rect 12618 15960 12624 15972
rect 11940 15932 12624 15960
rect 11940 15920 11946 15932
rect 12618 15920 12624 15932
rect 12676 15960 12682 15972
rect 13004 15960 13032 16000
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17037 16031 17095 16037
rect 17037 16028 17049 16031
rect 17000 16000 17049 16028
rect 17000 15988 17006 16000
rect 17037 15997 17049 16000
rect 17083 15997 17095 16031
rect 18782 16028 18788 16040
rect 18743 16000 18788 16028
rect 17037 15991 17095 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19300 16000 19533 16028
rect 19300 15988 19306 16000
rect 19521 15997 19533 16000
rect 19567 16028 19579 16031
rect 19567 16000 22876 16028
rect 19567 15997 19579 16000
rect 19521 15991 19579 15997
rect 12676 15932 13032 15960
rect 14476 15932 19334 15960
rect 12676 15920 12682 15932
rect 14476 15904 14504 15932
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2317 15895 2375 15901
rect 2317 15861 2329 15895
rect 2363 15892 2375 15895
rect 2590 15892 2596 15904
rect 2363 15864 2596 15892
rect 2363 15861 2375 15864
rect 2317 15855 2375 15861
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 9401 15895 9459 15901
rect 9401 15861 9413 15895
rect 9447 15892 9459 15895
rect 9950 15892 9956 15904
rect 9447 15864 9956 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10870 15892 10876 15904
rect 10831 15864 10876 15892
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 10962 15852 10968 15904
rect 11020 15892 11026 15904
rect 11977 15895 12035 15901
rect 11977 15892 11989 15895
rect 11020 15864 11989 15892
rect 11020 15852 11026 15864
rect 11977 15861 11989 15864
rect 12023 15892 12035 15895
rect 14274 15892 14280 15904
rect 12023 15864 14280 15892
rect 12023 15861 12035 15864
rect 11977 15855 12035 15861
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14458 15892 14464 15904
rect 14419 15864 14464 15892
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15749 15895 15807 15901
rect 15749 15861 15761 15895
rect 15795 15892 15807 15895
rect 16022 15892 16028 15904
rect 15795 15864 16028 15892
rect 15795 15861 15807 15864
rect 15749 15855 15807 15861
rect 16022 15852 16028 15864
rect 16080 15852 16086 15904
rect 19306 15892 19334 15932
rect 20806 15920 20812 15972
rect 20864 15960 20870 15972
rect 21910 15960 21916 15972
rect 20864 15932 21916 15960
rect 20864 15920 20870 15932
rect 21910 15920 21916 15932
rect 21968 15960 21974 15972
rect 22097 15963 22155 15969
rect 22097 15960 22109 15963
rect 21968 15932 22109 15960
rect 21968 15920 21974 15932
rect 22097 15929 22109 15932
rect 22143 15929 22155 15963
rect 22097 15923 22155 15929
rect 22189 15963 22247 15969
rect 22189 15929 22201 15963
rect 22235 15960 22247 15963
rect 22370 15960 22376 15972
rect 22235 15932 22376 15960
rect 22235 15929 22247 15932
rect 22189 15923 22247 15929
rect 22370 15920 22376 15932
rect 22428 15920 22434 15972
rect 22848 15960 22876 16000
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 23860 16037 23888 16068
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 25240 16105 25268 16136
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16065 25283 16099
rect 25406 16096 25412 16108
rect 25367 16068 25412 16096
rect 25225 16059 25283 16065
rect 25406 16056 25412 16068
rect 25464 16056 25470 16108
rect 23845 16031 23903 16037
rect 22980 16000 23025 16028
rect 22980 15988 22986 16000
rect 23845 15997 23857 16031
rect 23891 16028 23903 16031
rect 25424 16028 25452 16056
rect 23891 16000 25452 16028
rect 25516 16028 25544 16136
rect 27080 16136 28212 16164
rect 29415 16136 29460 16164
rect 25866 16056 25872 16108
rect 25924 16096 25930 16108
rect 25961 16099 26019 16105
rect 25961 16096 25973 16099
rect 25924 16068 25973 16096
rect 25924 16056 25930 16068
rect 25961 16065 25973 16068
rect 26007 16065 26019 16099
rect 26234 16096 26240 16108
rect 26195 16068 26240 16096
rect 25961 16059 26019 16065
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 26970 16096 26976 16108
rect 26883 16068 26976 16096
rect 26970 16056 26976 16068
rect 27028 16096 27034 16108
rect 27080 16096 27108 16136
rect 29454 16124 29460 16136
rect 29512 16124 29518 16176
rect 27028 16068 27108 16096
rect 27157 16099 27215 16105
rect 27028 16056 27034 16068
rect 27157 16065 27169 16099
rect 27203 16065 27215 16099
rect 27430 16096 27436 16108
rect 27391 16068 27436 16096
rect 27157 16059 27215 16065
rect 26878 16028 26884 16040
rect 25516 16000 26884 16028
rect 23891 15997 23903 16000
rect 23845 15991 23903 15997
rect 26878 15988 26884 16000
rect 26936 16028 26942 16040
rect 27172 16028 27200 16059
rect 27430 16056 27436 16068
rect 27488 16056 27494 16108
rect 29273 16099 29331 16105
rect 29273 16096 29285 16099
rect 28644 16068 29285 16096
rect 26936 16000 27200 16028
rect 26936 15988 26942 16000
rect 28644 15969 28672 16068
rect 29273 16065 29285 16068
rect 29319 16065 29331 16099
rect 29273 16059 29331 16065
rect 33042 16056 33048 16108
rect 33100 16096 33106 16108
rect 33137 16099 33195 16105
rect 33137 16096 33149 16099
rect 33100 16068 33149 16096
rect 33100 16056 33106 16068
rect 33137 16065 33149 16068
rect 33183 16065 33195 16099
rect 33137 16059 33195 16065
rect 36998 16056 37004 16108
rect 37056 16096 37062 16108
rect 37553 16099 37611 16105
rect 37553 16096 37565 16099
rect 37056 16068 37565 16096
rect 37056 16056 37062 16068
rect 37553 16065 37565 16068
rect 37599 16065 37611 16099
rect 37553 16059 37611 16065
rect 33226 15988 33232 16040
rect 33284 16028 33290 16040
rect 33413 16031 33471 16037
rect 33413 16028 33425 16031
rect 33284 16000 33425 16028
rect 33284 15988 33290 16000
rect 33413 15997 33425 16000
rect 33459 16028 33471 16031
rect 34238 16028 34244 16040
rect 33459 16000 34244 16028
rect 33459 15997 33471 16000
rect 33413 15991 33471 15997
rect 34238 15988 34244 16000
rect 34296 16028 34302 16040
rect 34517 16031 34575 16037
rect 34517 16028 34529 16031
rect 34296 16000 34529 16028
rect 34296 15988 34302 16000
rect 34517 15997 34529 16000
rect 34563 15997 34575 16031
rect 34517 15991 34575 15997
rect 35710 15988 35716 16040
rect 35768 16028 35774 16040
rect 35897 16031 35955 16037
rect 35897 16028 35909 16031
rect 35768 16000 35909 16028
rect 35768 15988 35774 16000
rect 35897 15997 35909 16000
rect 35943 15997 35955 16031
rect 35897 15991 35955 15997
rect 36173 16031 36231 16037
rect 36173 15997 36185 16031
rect 36219 15997 36231 16031
rect 37274 16028 37280 16040
rect 37235 16000 37280 16028
rect 36173 15991 36231 15997
rect 28629 15963 28687 15969
rect 28629 15960 28641 15963
rect 22848 15932 28641 15960
rect 28629 15929 28641 15932
rect 28675 15929 28687 15963
rect 34790 15960 34796 15972
rect 34751 15932 34796 15960
rect 28629 15923 28687 15929
rect 34790 15920 34796 15932
rect 34848 15920 34854 15972
rect 36188 15960 36216 15991
rect 37274 15988 37280 16000
rect 37332 15988 37338 16040
rect 37458 15960 37464 15972
rect 36188 15932 37464 15960
rect 37458 15920 37464 15932
rect 37516 15920 37522 15972
rect 21818 15892 21824 15904
rect 19306 15864 21824 15892
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 22922 15892 22928 15904
rect 22520 15864 22928 15892
rect 22520 15852 22526 15864
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 23109 15895 23167 15901
rect 23109 15861 23121 15895
rect 23155 15892 23167 15895
rect 23290 15892 23296 15904
rect 23155 15864 23296 15892
rect 23155 15861 23167 15864
rect 23109 15855 23167 15861
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 25222 15852 25228 15904
rect 25280 15892 25286 15904
rect 26053 15895 26111 15901
rect 26053 15892 26065 15895
rect 25280 15864 26065 15892
rect 25280 15852 25286 15864
rect 26053 15861 26065 15864
rect 26099 15861 26111 15895
rect 26053 15855 26111 15861
rect 34977 15895 35035 15901
rect 34977 15861 34989 15895
rect 35023 15892 35035 15895
rect 35618 15892 35624 15904
rect 35023 15864 35624 15892
rect 35023 15861 35035 15864
rect 34977 15855 35035 15861
rect 35618 15852 35624 15864
rect 35676 15852 35682 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 2133 15691 2191 15697
rect 2133 15657 2145 15691
rect 2179 15688 2191 15691
rect 7466 15688 7472 15700
rect 2179 15660 7472 15688
rect 2179 15657 2191 15660
rect 2133 15651 2191 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8938 15688 8944 15700
rect 8899 15660 8944 15688
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 9309 15691 9367 15697
rect 9309 15657 9321 15691
rect 9355 15688 9367 15691
rect 9766 15688 9772 15700
rect 9355 15660 9772 15688
rect 9355 15657 9367 15660
rect 9309 15651 9367 15657
rect 9766 15648 9772 15660
rect 9824 15688 9830 15700
rect 10686 15688 10692 15700
rect 9824 15660 10692 15688
rect 9824 15648 9830 15660
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 11882 15688 11888 15700
rect 11843 15660 11888 15688
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 13078 15688 13084 15700
rect 13004 15660 13084 15688
rect 13004 15620 13032 15660
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 13265 15691 13323 15697
rect 13265 15657 13277 15691
rect 13311 15688 13323 15691
rect 14366 15688 14372 15700
rect 13311 15660 14372 15688
rect 13311 15657 13323 15660
rect 13265 15651 13323 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 16206 15688 16212 15700
rect 14783 15660 16212 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 21818 15688 21824 15700
rect 16316 15660 21036 15688
rect 21779 15660 21824 15688
rect 13170 15620 13176 15632
rect 9416 15592 13032 15620
rect 13131 15592 13176 15620
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9416 15493 9444 15592
rect 13170 15580 13176 15592
rect 13228 15580 13234 15632
rect 14274 15580 14280 15632
rect 14332 15620 14338 15632
rect 16316 15620 16344 15660
rect 14332 15592 16344 15620
rect 16393 15623 16451 15629
rect 14332 15580 14338 15592
rect 16393 15589 16405 15623
rect 16439 15620 16451 15623
rect 16850 15620 16856 15632
rect 16439 15592 16856 15620
rect 16439 15589 16451 15592
rect 16393 15583 16451 15589
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 17034 15580 17040 15632
rect 17092 15620 17098 15632
rect 18230 15620 18236 15632
rect 17092 15592 18236 15620
rect 17092 15580 17098 15592
rect 18230 15580 18236 15592
rect 18288 15620 18294 15632
rect 18693 15623 18751 15629
rect 18693 15620 18705 15623
rect 18288 15592 18705 15620
rect 18288 15580 18294 15592
rect 18693 15589 18705 15592
rect 18739 15589 18751 15623
rect 18693 15583 18751 15589
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 12802 15552 12808 15564
rect 10827 15524 12808 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 1854 15416 1860 15428
rect 1815 15388 1860 15416
rect 1854 15376 1860 15388
rect 1912 15416 1918 15428
rect 2685 15419 2743 15425
rect 2685 15416 2697 15419
rect 1912 15388 2697 15416
rect 1912 15376 1918 15388
rect 2685 15385 2697 15388
rect 2731 15385 2743 15419
rect 9416 15416 9444 15447
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 12544 15493 12572 15524
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 12986 15552 12992 15564
rect 12947 15524 12992 15552
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 16022 15552 16028 15564
rect 15983 15524 16028 15552
rect 16022 15512 16028 15524
rect 16080 15512 16086 15564
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 20714 15552 20720 15564
rect 20119 15524 20720 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20864 15524 20909 15552
rect 20864 15512 20870 15524
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 10928 15456 12081 15484
rect 10928 15444 10934 15456
rect 12069 15453 12081 15456
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 12575 15456 12609 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 2685 15379 2743 15385
rect 8312 15388 9444 15416
rect 12161 15419 12219 15425
rect 8312 15360 8340 15388
rect 12161 15385 12173 15419
rect 12207 15385 12219 15419
rect 12161 15379 12219 15385
rect 8294 15348 8300 15360
rect 8255 15320 8300 15348
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 11204 15320 11345 15348
rect 11204 15308 11210 15320
rect 11333 15317 11345 15320
rect 11379 15348 11391 15351
rect 12176 15348 12204 15379
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 12452 15416 12480 15447
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 14550 15484 14556 15496
rect 13320 15456 13365 15484
rect 14511 15456 14556 15484
rect 13320 15444 13326 15456
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15252 15456 15485 15484
rect 15252 15444 15258 15456
rect 15473 15453 15485 15456
rect 15519 15484 15531 15487
rect 15519 15456 16068 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 12894 15416 12900 15428
rect 12308 15388 12353 15416
rect 12452 15388 12900 15416
rect 12308 15376 12314 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 13446 15376 13452 15428
rect 13504 15416 13510 15428
rect 15289 15419 15347 15425
rect 15289 15416 15301 15419
rect 13504 15388 15301 15416
rect 13504 15376 13510 15388
rect 15289 15385 15301 15388
rect 15335 15385 15347 15419
rect 15289 15379 15347 15385
rect 15654 15376 15660 15428
rect 15712 15416 15718 15428
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 15712 15388 15945 15416
rect 15712 15376 15718 15388
rect 15933 15385 15945 15388
rect 15979 15385 15991 15419
rect 16040 15416 16068 15456
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 16172 15456 16221 15484
rect 16172 15444 16178 15456
rect 16209 15453 16221 15456
rect 16255 15484 16267 15487
rect 16390 15484 16396 15496
rect 16255 15456 16396 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 19058 15484 19064 15496
rect 18472 15456 19064 15484
rect 18472 15444 18478 15456
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 19392 15456 19809 15484
rect 19392 15444 19398 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 20533 15487 20591 15493
rect 20533 15453 20545 15487
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 17405 15419 17463 15425
rect 17405 15416 17417 15419
rect 16040 15388 17417 15416
rect 15933 15379 15991 15385
rect 17405 15385 17417 15388
rect 17451 15385 17463 15419
rect 18506 15416 18512 15428
rect 18419 15388 18512 15416
rect 17405 15379 17463 15385
rect 18506 15376 18512 15388
rect 18564 15416 18570 15428
rect 20548 15416 20576 15447
rect 18564 15388 20576 15416
rect 18564 15376 18570 15388
rect 11379 15320 12204 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 17494 15348 17500 15360
rect 16540 15320 17500 15348
rect 16540 15308 16546 15320
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 21008 15348 21036 15660
rect 21818 15648 21824 15660
rect 21876 15688 21882 15700
rect 23290 15688 23296 15700
rect 21876 15660 23296 15688
rect 21876 15648 21882 15660
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 25133 15691 25191 15697
rect 25133 15657 25145 15691
rect 25179 15688 25191 15691
rect 25222 15688 25228 15700
rect 25179 15660 25228 15688
rect 25179 15657 25191 15660
rect 25133 15651 25191 15657
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 35805 15691 35863 15697
rect 35805 15657 35817 15691
rect 35851 15688 35863 15691
rect 35894 15688 35900 15700
rect 35851 15660 35900 15688
rect 35851 15657 35863 15660
rect 35805 15651 35863 15657
rect 35894 15648 35900 15660
rect 35952 15648 35958 15700
rect 21726 15580 21732 15632
rect 21784 15620 21790 15632
rect 22281 15623 22339 15629
rect 22281 15620 22293 15623
rect 21784 15592 22293 15620
rect 21784 15580 21790 15592
rect 22281 15589 22293 15592
rect 22327 15589 22339 15623
rect 22281 15583 22339 15589
rect 22833 15623 22891 15629
rect 22833 15589 22845 15623
rect 22879 15620 22891 15623
rect 27062 15620 27068 15632
rect 22879 15592 27068 15620
rect 22879 15589 22891 15592
rect 22833 15583 22891 15589
rect 21913 15555 21971 15561
rect 21913 15521 21925 15555
rect 21959 15552 21971 15555
rect 22002 15552 22008 15564
rect 21959 15524 22008 15552
rect 21959 15521 21971 15524
rect 21913 15515 21971 15521
rect 22002 15512 22008 15524
rect 22060 15552 22066 15564
rect 22462 15552 22468 15564
rect 22060 15524 22468 15552
rect 22060 15512 22066 15524
rect 22462 15512 22468 15524
rect 22520 15512 22526 15564
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 21600 15456 21833 15484
rect 21600 15444 21606 15456
rect 21821 15453 21833 15456
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 22097 15487 22155 15493
rect 22097 15453 22109 15487
rect 22143 15484 22155 15487
rect 22848 15484 22876 15583
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 22143 15456 22876 15484
rect 25777 15487 25835 15493
rect 22143 15453 22155 15456
rect 22097 15447 22155 15453
rect 25777 15453 25789 15487
rect 25823 15484 25835 15487
rect 30006 15484 30012 15496
rect 25823 15456 30012 15484
rect 25823 15453 25835 15456
rect 25777 15447 25835 15453
rect 30006 15444 30012 15456
rect 30064 15444 30070 15496
rect 35618 15484 35624 15496
rect 35579 15456 35624 15484
rect 35618 15444 35624 15456
rect 35676 15444 35682 15496
rect 36998 15493 37004 15496
rect 36996 15484 37004 15493
rect 36959 15456 37004 15484
rect 36996 15447 37004 15456
rect 36998 15444 37004 15447
rect 37056 15444 37062 15496
rect 37182 15484 37188 15496
rect 37143 15456 37188 15484
rect 37182 15444 37188 15456
rect 37240 15444 37246 15496
rect 37366 15484 37372 15496
rect 37327 15456 37372 15484
rect 37366 15444 37372 15456
rect 37424 15444 37430 15496
rect 37458 15444 37464 15496
rect 37516 15484 37522 15496
rect 38102 15484 38108 15496
rect 37516 15456 37561 15484
rect 38063 15456 38108 15484
rect 37516 15444 37522 15456
rect 38102 15444 38108 15456
rect 38160 15444 38166 15496
rect 24581 15419 24639 15425
rect 24581 15385 24593 15419
rect 24627 15416 24639 15419
rect 25958 15416 25964 15428
rect 24627 15388 25728 15416
rect 25919 15388 25964 15416
rect 24627 15385 24639 15388
rect 24581 15379 24639 15385
rect 24596 15348 24624 15379
rect 25590 15348 25596 15360
rect 21008 15320 24624 15348
rect 25551 15320 25596 15348
rect 25590 15308 25596 15320
rect 25648 15308 25654 15360
rect 25700 15348 25728 15388
rect 25958 15376 25964 15388
rect 26016 15376 26022 15428
rect 27062 15376 27068 15428
rect 27120 15416 27126 15428
rect 27433 15419 27491 15425
rect 27433 15416 27445 15419
rect 27120 15388 27445 15416
rect 27120 15376 27126 15388
rect 27433 15385 27445 15388
rect 27479 15416 27491 15419
rect 33410 15416 33416 15428
rect 27479 15388 33416 15416
rect 27479 15385 27491 15388
rect 27433 15379 27491 15385
rect 33410 15376 33416 15388
rect 33468 15376 33474 15428
rect 37090 15416 37096 15428
rect 34256 15388 36860 15416
rect 37051 15388 37096 15416
rect 26878 15348 26884 15360
rect 25700 15320 26884 15348
rect 26878 15308 26884 15320
rect 26936 15308 26942 15360
rect 28994 15308 29000 15360
rect 29052 15348 29058 15360
rect 34256 15348 34284 15388
rect 36832 15357 36860 15388
rect 37090 15376 37096 15388
rect 37148 15376 37154 15428
rect 29052 15320 34284 15348
rect 36817 15351 36875 15357
rect 29052 15308 29058 15320
rect 36817 15317 36829 15351
rect 36863 15317 36875 15351
rect 36817 15311 36875 15317
rect 37366 15308 37372 15360
rect 37424 15348 37430 15360
rect 37921 15351 37979 15357
rect 37921 15348 37933 15351
rect 37424 15320 37933 15348
rect 37424 15308 37430 15320
rect 37921 15317 37933 15320
rect 37967 15317 37979 15351
rect 37921 15311 37979 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 6270 15144 6276 15156
rect 2280 15116 6276 15144
rect 2280 15104 2286 15116
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 17310 15144 17316 15156
rect 10008 15116 15792 15144
rect 17271 15116 17316 15144
rect 10008 15104 10014 15116
rect 10965 15079 11023 15085
rect 10965 15045 10977 15079
rect 11011 15076 11023 15079
rect 11054 15076 11060 15088
rect 11011 15048 11060 15076
rect 11011 15045 11023 15048
rect 10965 15039 11023 15045
rect 11054 15036 11060 15048
rect 11112 15076 11118 15088
rect 12069 15079 12127 15085
rect 12069 15076 12081 15079
rect 11112 15048 12081 15076
rect 11112 15036 11118 15048
rect 12069 15045 12081 15048
rect 12115 15045 12127 15079
rect 12069 15039 12127 15045
rect 14366 15036 14372 15088
rect 14424 15076 14430 15088
rect 14553 15079 14611 15085
rect 14553 15076 14565 15079
rect 14424 15048 14565 15076
rect 14424 15036 14430 15048
rect 14553 15045 14565 15048
rect 14599 15045 14611 15079
rect 14553 15039 14611 15045
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 15008 1458 15020
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 1452 14980 2053 15008
rect 1452 14968 1458 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 14458 15008 14464 15020
rect 13403 14980 14464 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15654 15008 15660 15020
rect 15344 14980 15660 15008
rect 15344 14968 15350 14980
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 15764 15008 15792 15116
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 35710 15144 35716 15156
rect 18748 15116 31754 15144
rect 35671 15116 35716 15144
rect 18748 15104 18754 15116
rect 17678 15076 17684 15088
rect 16684 15048 17684 15076
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15764 14980 15945 15008
rect 15933 14977 15945 14980
rect 15979 15008 15991 15011
rect 16684 15008 16712 15048
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18322 15085 18328 15088
rect 18050 15079 18108 15085
rect 18050 15076 18062 15079
rect 18012 15048 18062 15076
rect 18012 15036 18018 15048
rect 18050 15045 18062 15048
rect 18096 15045 18108 15079
rect 18050 15039 18108 15045
rect 18279 15079 18328 15085
rect 18279 15045 18291 15079
rect 18325 15045 18328 15079
rect 18279 15039 18328 15045
rect 18322 15036 18328 15039
rect 18380 15036 18386 15088
rect 20530 15036 20536 15088
rect 20588 15076 20594 15088
rect 22370 15076 22376 15088
rect 20588 15048 22376 15076
rect 20588 15036 20594 15048
rect 22370 15036 22376 15048
rect 22428 15036 22434 15088
rect 22646 15036 22652 15088
rect 22704 15076 22710 15088
rect 25130 15076 25136 15088
rect 22704 15048 25136 15076
rect 22704 15036 22710 15048
rect 25130 15036 25136 15048
rect 25188 15036 25194 15088
rect 25498 15036 25504 15088
rect 25556 15076 25562 15088
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 25556 15048 25697 15076
rect 25556 15036 25562 15048
rect 25685 15045 25697 15048
rect 25731 15076 25743 15079
rect 25866 15076 25872 15088
rect 25731 15048 25872 15076
rect 25731 15045 25743 15048
rect 25685 15039 25743 15045
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 26329 15079 26387 15085
rect 26329 15045 26341 15079
rect 26375 15076 26387 15079
rect 26878 15076 26884 15088
rect 26375 15048 26884 15076
rect 26375 15045 26387 15048
rect 26329 15039 26387 15045
rect 26878 15036 26884 15048
rect 26936 15036 26942 15088
rect 31726 15076 31754 15116
rect 35710 15104 35716 15116
rect 35768 15104 35774 15156
rect 36725 15147 36783 15153
rect 36725 15113 36737 15147
rect 36771 15144 36783 15147
rect 37642 15144 37648 15156
rect 36771 15116 37648 15144
rect 36771 15113 36783 15116
rect 36725 15107 36783 15113
rect 37642 15104 37648 15116
rect 37700 15104 37706 15156
rect 38010 15144 38016 15156
rect 37971 15116 38016 15144
rect 38010 15104 38016 15116
rect 38068 15104 38074 15156
rect 37274 15076 37280 15088
rect 31726 15048 37280 15076
rect 37274 15036 37280 15048
rect 37332 15036 37338 15088
rect 16850 15008 16856 15020
rect 15979 14980 16712 15008
rect 16811 14980 16856 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 17126 15008 17132 15020
rect 17087 14980 17132 15008
rect 17126 14968 17132 14980
rect 17184 14968 17190 15020
rect 18141 15011 18199 15017
rect 17958 15001 18016 15007
rect 17958 14998 17970 15001
rect 17880 14970 17970 14998
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 15749 14943 15807 14949
rect 15749 14940 15761 14943
rect 15436 14912 15761 14940
rect 15436 14900 15442 14912
rect 15749 14909 15761 14912
rect 15795 14940 15807 14943
rect 16022 14940 16028 14952
rect 15795 14912 16028 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 17034 14940 17040 14952
rect 16995 14912 17040 14940
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 12986 14872 12992 14884
rect 12299 14844 12992 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 13170 14872 13176 14884
rect 13131 14844 13176 14872
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 14734 14872 14740 14884
rect 14695 14844 14740 14872
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 16206 14872 16212 14884
rect 15948 14844 16212 14872
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 2498 14804 2504 14816
rect 1627 14776 2504 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 14001 14807 14059 14813
rect 14001 14804 14013 14807
rect 12952 14776 14013 14804
rect 12952 14764 12958 14776
rect 14001 14773 14013 14776
rect 14047 14804 14059 14807
rect 15654 14804 15660 14816
rect 14047 14776 15660 14804
rect 14047 14773 14059 14776
rect 14001 14767 14059 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 15948 14813 15976 14844
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 16850 14832 16856 14884
rect 16908 14872 16914 14884
rect 16945 14875 17003 14881
rect 16945 14872 16957 14875
rect 16908 14844 16957 14872
rect 16908 14832 16914 14844
rect 16945 14841 16957 14844
rect 16991 14841 17003 14875
rect 16945 14835 17003 14841
rect 15933 14807 15991 14813
rect 15933 14773 15945 14807
rect 15979 14773 15991 14807
rect 15933 14767 15991 14773
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 16080 14776 16129 14804
rect 16080 14764 16086 14776
rect 16117 14773 16129 14776
rect 16163 14773 16175 14807
rect 17770 14804 17776 14816
rect 17731 14776 17776 14804
rect 16117 14767 16175 14773
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 17880 14804 17908 14970
rect 17958 14967 17970 14970
rect 18004 14967 18016 15001
rect 18141 14977 18153 15011
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 17958 14961 18016 14967
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 18156 14872 18184 14971
rect 21542 14968 21548 15020
rect 21600 15008 21606 15020
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21600 14980 21833 15008
rect 21600 14968 21606 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 21821 14971 21879 14977
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 22143 14980 22845 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22833 14977 22845 14980
rect 22879 15008 22891 15011
rect 28902 15008 28908 15020
rect 22879 14980 28908 15008
rect 22879 14977 22891 14980
rect 22833 14971 22891 14977
rect 28902 14968 28908 14980
rect 28960 14968 28966 15020
rect 34698 15008 34704 15020
rect 34659 14980 34704 15008
rect 34698 14968 34704 14980
rect 34756 14968 34762 15020
rect 37829 15011 37887 15017
rect 37829 14977 37841 15011
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 18417 14943 18475 14949
rect 18417 14909 18429 14943
rect 18463 14940 18475 14943
rect 18598 14940 18604 14952
rect 18463 14912 18604 14940
rect 18463 14909 18475 14912
rect 18417 14903 18475 14909
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18892 14912 21588 14940
rect 18012 14844 18184 14872
rect 18012 14832 18018 14844
rect 18782 14832 18788 14884
rect 18840 14872 18846 14884
rect 18892 14881 18920 14912
rect 18877 14875 18935 14881
rect 18877 14872 18889 14875
rect 18840 14844 18889 14872
rect 18840 14832 18846 14844
rect 18877 14841 18889 14844
rect 18923 14841 18935 14875
rect 18877 14835 18935 14841
rect 18966 14832 18972 14884
rect 19024 14872 19030 14884
rect 19334 14872 19340 14884
rect 19024 14844 19340 14872
rect 19024 14832 19030 14844
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 20717 14875 20775 14881
rect 20717 14841 20729 14875
rect 20763 14872 20775 14875
rect 21450 14872 21456 14884
rect 20763 14844 21456 14872
rect 20763 14841 20775 14844
rect 20717 14835 20775 14841
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 21560 14872 21588 14912
rect 22940 14912 30052 14940
rect 22278 14872 22284 14884
rect 21560 14844 22094 14872
rect 22239 14844 22284 14872
rect 18046 14804 18052 14816
rect 17880 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 21177 14807 21235 14813
rect 21177 14804 21189 14807
rect 20588 14776 21189 14804
rect 20588 14764 20594 14776
rect 21177 14773 21189 14776
rect 21223 14773 21235 14807
rect 21818 14804 21824 14816
rect 21779 14776 21824 14804
rect 21177 14767 21235 14773
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 22066 14804 22094 14844
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 22940 14804 22968 14912
rect 29914 14872 29920 14884
rect 29875 14844 29920 14872
rect 29914 14832 29920 14844
rect 29972 14832 29978 14884
rect 30024 14872 30052 14912
rect 30098 14900 30104 14952
rect 30156 14940 30162 14952
rect 30285 14943 30343 14949
rect 30285 14940 30297 14943
rect 30156 14912 30297 14940
rect 30156 14900 30162 14912
rect 30285 14909 30297 14912
rect 30331 14909 30343 14943
rect 30285 14903 30343 14909
rect 31754 14900 31760 14952
rect 31812 14940 31818 14952
rect 37844 14940 37872 14971
rect 31812 14912 37872 14940
rect 31812 14900 31818 14912
rect 36814 14872 36820 14884
rect 30024 14844 36820 14872
rect 36814 14832 36820 14844
rect 36872 14832 36878 14884
rect 22066 14776 22968 14804
rect 25133 14807 25191 14813
rect 25133 14773 25145 14807
rect 25179 14804 25191 14807
rect 25222 14804 25228 14816
rect 25179 14776 25228 14804
rect 25179 14773 25191 14776
rect 25133 14767 25191 14773
rect 25222 14764 25228 14776
rect 25280 14804 25286 14816
rect 25406 14804 25412 14816
rect 25280 14776 25412 14804
rect 25280 14764 25286 14776
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 25774 14764 25780 14816
rect 25832 14804 25838 14816
rect 27338 14804 27344 14816
rect 25832 14776 27344 14804
rect 25832 14764 25838 14776
rect 27338 14764 27344 14776
rect 27396 14764 27402 14816
rect 29178 14764 29184 14816
rect 29236 14804 29242 14816
rect 29825 14807 29883 14813
rect 29825 14804 29837 14807
rect 29236 14776 29837 14804
rect 29236 14764 29242 14776
rect 29825 14773 29837 14776
rect 29871 14773 29883 14807
rect 29825 14767 29883 14773
rect 34790 14764 34796 14816
rect 34848 14804 34854 14816
rect 34885 14807 34943 14813
rect 34885 14804 34897 14807
rect 34848 14776 34897 14804
rect 34848 14764 34854 14776
rect 34885 14773 34897 14776
rect 34931 14773 34943 14807
rect 34885 14767 34943 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 14458 14600 14464 14612
rect 13372 14572 14464 14600
rect 11885 14535 11943 14541
rect 11885 14501 11897 14535
rect 11931 14532 11943 14535
rect 13372 14532 13400 14572
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 15562 14600 15568 14612
rect 15475 14572 15568 14600
rect 15562 14560 15568 14572
rect 15620 14600 15626 14612
rect 16206 14600 16212 14612
rect 15620 14572 16212 14600
rect 15620 14560 15626 14572
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 23658 14600 23664 14612
rect 18104 14572 23664 14600
rect 18104 14560 18110 14572
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 31754 14560 31760 14612
rect 31812 14600 31818 14612
rect 34054 14600 34060 14612
rect 31812 14572 31857 14600
rect 34015 14572 34060 14600
rect 31812 14560 31818 14572
rect 34054 14560 34060 14572
rect 34112 14560 34118 14612
rect 34698 14560 34704 14612
rect 34756 14600 34762 14612
rect 35161 14603 35219 14609
rect 35161 14600 35173 14603
rect 34756 14572 35173 14600
rect 34756 14560 34762 14572
rect 35161 14569 35173 14572
rect 35207 14569 35219 14603
rect 38102 14600 38108 14612
rect 38063 14572 38108 14600
rect 35161 14563 35219 14569
rect 38102 14560 38108 14572
rect 38160 14560 38166 14612
rect 11931 14504 13400 14532
rect 13449 14535 13507 14541
rect 11931 14501 11943 14504
rect 11885 14495 11943 14501
rect 13449 14501 13461 14535
rect 13495 14532 13507 14535
rect 13906 14532 13912 14544
rect 13495 14504 13912 14532
rect 13495 14501 13507 14504
rect 13449 14495 13507 14501
rect 13906 14492 13912 14504
rect 13964 14532 13970 14544
rect 14550 14532 14556 14544
rect 13964 14504 14556 14532
rect 13964 14492 13970 14504
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 15654 14492 15660 14544
rect 15712 14532 15718 14544
rect 18690 14532 18696 14544
rect 15712 14504 18696 14532
rect 15712 14492 15718 14504
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 34422 14492 34428 14544
rect 34480 14532 34486 14544
rect 34977 14535 35035 14541
rect 34977 14532 34989 14535
rect 34480 14504 34989 14532
rect 34480 14492 34486 14504
rect 34977 14501 34989 14504
rect 35023 14501 35035 14535
rect 34977 14495 35035 14501
rect 36817 14535 36875 14541
rect 36817 14501 36829 14535
rect 36863 14501 36875 14535
rect 36817 14495 36875 14501
rect 15378 14464 15384 14476
rect 15339 14436 15384 14464
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15580 14436 16221 14464
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12986 14396 12992 14408
rect 12115 14368 12992 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12986 14356 12992 14368
rect 13044 14396 13050 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13044 14368 13277 14396
rect 13044 14356 13050 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 15286 14396 15292 14408
rect 14700 14368 15292 14396
rect 14700 14356 14706 14368
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 15580 14405 15608 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 25590 14464 25596 14476
rect 16209 14427 16267 14433
rect 17236 14436 25596 14464
rect 17236 14405 17264 14436
rect 25590 14424 25596 14436
rect 25648 14424 25654 14476
rect 25958 14424 25964 14476
rect 26016 14464 26022 14476
rect 36832 14464 36860 14495
rect 26016 14436 30512 14464
rect 26016 14424 26022 14436
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 15528 14368 15577 14396
rect 15528 14356 15534 14368
rect 15565 14365 15577 14368
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14365 17279 14399
rect 17678 14396 17684 14408
rect 17639 14368 17684 14396
rect 17221 14359 17279 14365
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 17920 14368 18153 14396
rect 17920 14356 17926 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 30282 14356 30288 14408
rect 30340 14396 30346 14408
rect 30377 14399 30435 14405
rect 30377 14396 30389 14399
rect 30340 14368 30389 14396
rect 30340 14356 30346 14368
rect 30377 14365 30389 14368
rect 30423 14365 30435 14399
rect 30484 14396 30512 14436
rect 31726 14436 36860 14464
rect 31726 14396 31754 14436
rect 35986 14396 35992 14408
rect 30484 14368 31754 14396
rect 35947 14368 35992 14396
rect 30377 14359 30435 14365
rect 35986 14356 35992 14368
rect 36044 14356 36050 14408
rect 36998 14405 37004 14408
rect 36996 14396 37004 14405
rect 36959 14368 37004 14396
rect 36996 14359 37004 14368
rect 36998 14356 37004 14359
rect 37056 14356 37062 14408
rect 37182 14396 37188 14408
rect 37143 14368 37188 14396
rect 37182 14356 37188 14368
rect 37240 14356 37246 14408
rect 37366 14396 37372 14408
rect 37327 14368 37372 14396
rect 37366 14356 37372 14368
rect 37424 14356 37430 14408
rect 37458 14356 37464 14408
rect 37516 14396 37522 14408
rect 37516 14368 37609 14396
rect 37516 14356 37522 14368
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 2133 14331 2191 14337
rect 2133 14328 2145 14331
rect 1452 14300 2145 14328
rect 1452 14288 1458 14300
rect 2133 14297 2145 14300
rect 2179 14297 2191 14331
rect 2133 14291 2191 14297
rect 12342 14288 12348 14340
rect 12400 14328 12406 14340
rect 12529 14331 12587 14337
rect 12529 14328 12541 14331
rect 12400 14300 12541 14328
rect 12400 14288 12406 14300
rect 12529 14297 12541 14300
rect 12575 14297 12587 14331
rect 12529 14291 12587 14297
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 12713 14331 12771 14337
rect 12713 14328 12725 14331
rect 12676 14300 12725 14328
rect 12676 14288 12682 14300
rect 12713 14297 12725 14300
rect 12759 14297 12771 14331
rect 12713 14291 12771 14297
rect 13078 14288 13084 14340
rect 13136 14328 13142 14340
rect 14553 14331 14611 14337
rect 14553 14328 14565 14331
rect 13136 14300 14565 14328
rect 13136 14288 13142 14300
rect 14553 14297 14565 14300
rect 14599 14297 14611 14331
rect 14553 14291 14611 14297
rect 14737 14331 14795 14337
rect 14737 14297 14749 14331
rect 14783 14328 14795 14331
rect 14918 14328 14924 14340
rect 14783 14300 14924 14328
rect 14783 14297 14795 14300
rect 14737 14291 14795 14297
rect 14918 14288 14924 14300
rect 14976 14328 14982 14340
rect 17313 14331 17371 14337
rect 14976 14300 17264 14328
rect 14976 14288 14982 14300
rect 17236 14272 17264 14300
rect 17313 14297 17325 14331
rect 17359 14297 17371 14331
rect 17313 14291 17371 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 9217 14263 9275 14269
rect 9217 14260 9229 14263
rect 2372 14232 9229 14260
rect 2372 14220 2378 14232
rect 9217 14229 9229 14232
rect 9263 14260 9275 14263
rect 9858 14260 9864 14272
rect 9263 14232 9864 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 13354 14260 13360 14272
rect 12952 14232 13360 14260
rect 12952 14220 12958 14232
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14260 15807 14263
rect 16114 14260 16120 14272
rect 15795 14232 16120 14260
rect 15795 14229 15807 14232
rect 15749 14223 15807 14229
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17034 14260 17040 14272
rect 16995 14232 17040 14260
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 17218 14220 17224 14272
rect 17276 14220 17282 14272
rect 17328 14260 17356 14291
rect 17402 14288 17408 14340
rect 17460 14328 17466 14340
rect 17586 14337 17592 14340
rect 17543 14331 17592 14337
rect 17460 14300 17505 14328
rect 17460 14288 17466 14300
rect 17543 14297 17555 14331
rect 17589 14297 17592 14331
rect 17543 14291 17592 14297
rect 17586 14288 17592 14291
rect 17644 14288 17650 14340
rect 17770 14288 17776 14340
rect 17828 14328 17834 14340
rect 21637 14331 21695 14337
rect 21637 14328 21649 14331
rect 17828 14300 21649 14328
rect 17828 14288 17834 14300
rect 21637 14297 21649 14300
rect 21683 14328 21695 14331
rect 21818 14328 21824 14340
rect 21683 14300 21824 14328
rect 21683 14297 21695 14300
rect 21637 14291 21695 14297
rect 21818 14288 21824 14300
rect 21876 14288 21882 14340
rect 29362 14288 29368 14340
rect 29420 14328 29426 14340
rect 30622 14331 30680 14337
rect 30622 14328 30634 14331
rect 29420 14300 30634 14328
rect 29420 14288 29426 14300
rect 30622 14297 30634 14300
rect 30668 14297 30680 14331
rect 30622 14291 30680 14297
rect 34238 14288 34244 14340
rect 34296 14328 34302 14340
rect 34701 14331 34759 14337
rect 34701 14328 34713 14331
rect 34296 14300 34713 14328
rect 34296 14288 34302 14300
rect 34701 14297 34713 14300
rect 34747 14297 34759 14331
rect 37090 14328 37096 14340
rect 37051 14300 37096 14328
rect 34701 14291 34759 14297
rect 37090 14288 37096 14300
rect 37148 14288 37154 14340
rect 37274 14288 37280 14340
rect 37332 14328 37338 14340
rect 37476 14328 37504 14356
rect 37332 14300 37504 14328
rect 37332 14288 37338 14300
rect 17862 14260 17868 14272
rect 17328 14232 17868 14260
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 29086 14220 29092 14272
rect 29144 14260 29150 14272
rect 29641 14263 29699 14269
rect 29641 14260 29653 14263
rect 29144 14232 29653 14260
rect 29144 14220 29150 14232
rect 29641 14229 29653 14232
rect 29687 14260 29699 14263
rect 30190 14260 30196 14272
rect 29687 14232 30196 14260
rect 29687 14229 29699 14232
rect 29641 14223 29699 14229
rect 30190 14220 30196 14232
rect 30248 14220 30254 14272
rect 36170 14260 36176 14272
rect 36131 14232 36176 14260
rect 36170 14220 36176 14232
rect 36228 14220 36234 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 8294 14056 8300 14068
rect 1688 14028 8300 14056
rect 1688 13997 1716 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8938 14056 8944 14068
rect 8851 14028 8944 14056
rect 8938 14016 8944 14028
rect 8996 14056 9002 14068
rect 13722 14056 13728 14068
rect 8996 14028 13728 14056
rect 8996 14016 9002 14028
rect 13722 14016 13728 14028
rect 13780 14056 13786 14068
rect 15565 14059 15623 14065
rect 13780 14028 14964 14056
rect 13780 14016 13786 14028
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13957 1731 13991
rect 2498 13988 2504 14000
rect 2459 13960 2504 13988
rect 1673 13951 1731 13957
rect 2498 13948 2504 13960
rect 2556 13948 2562 14000
rect 8110 13988 8116 14000
rect 7576 13960 8116 13988
rect 1394 13920 1400 13932
rect 1355 13892 1400 13920
rect 1394 13880 1400 13892
rect 1452 13880 1458 13932
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 7576 13929 7604 13960
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 12621 13991 12679 13997
rect 12492 13960 12537 13988
rect 12492 13948 12498 13960
rect 12621 13957 12633 13991
rect 12667 13988 12679 13991
rect 13262 13988 13268 14000
rect 12667 13960 13268 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 13262 13948 13268 13960
rect 13320 13988 13326 14000
rect 13630 13988 13636 14000
rect 13320 13960 13636 13988
rect 13320 13948 13326 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 14458 13948 14464 14000
rect 14516 13988 14522 14000
rect 14826 13988 14832 14000
rect 14516 13960 14832 13988
rect 14516 13948 14522 13960
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 7561 13923 7619 13929
rect 2832 13892 2877 13920
rect 2832 13880 2838 13892
rect 7561 13889 7573 13923
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 7828 13923 7886 13929
rect 7828 13889 7840 13923
rect 7874 13920 7886 13923
rect 9582 13920 9588 13932
rect 7874 13892 8616 13920
rect 9543 13892 9588 13920
rect 7874 13889 7886 13892
rect 7828 13883 7886 13889
rect 2590 13852 2596 13864
rect 2551 13824 2596 13852
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 8588 13784 8616 13892
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 9766 13920 9772 13932
rect 9727 13892 9772 13920
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 11790 13920 11796 13932
rect 9916 13892 11796 13920
rect 9916 13880 9922 13892
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 13354 13920 13360 13932
rect 12584 13892 13360 13920
rect 12584 13880 12590 13892
rect 13354 13880 13360 13892
rect 13412 13920 13418 13932
rect 13538 13920 13544 13932
rect 13412 13892 13544 13920
rect 13412 13880 13418 13892
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14182 13880 14188 13932
rect 14240 13920 14246 13932
rect 14642 13920 14648 13932
rect 14240 13892 14648 13920
rect 14240 13880 14246 13892
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 14936 13929 14964 14028
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 17678 14056 17684 14068
rect 15611 14028 17684 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 29086 14056 29092 14068
rect 17828 14028 29092 14056
rect 17828 14016 17834 14028
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 29362 14056 29368 14068
rect 29323 14028 29368 14056
rect 29362 14016 29368 14028
rect 29420 14016 29426 14068
rect 29825 14059 29883 14065
rect 29825 14025 29837 14059
rect 29871 14056 29883 14059
rect 29914 14056 29920 14068
rect 29871 14028 29920 14056
rect 29871 14025 29883 14028
rect 29825 14019 29883 14025
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 30190 14056 30196 14068
rect 30151 14028 30196 14056
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 31754 14056 31760 14068
rect 30300 14028 31760 14056
rect 15764 13960 17080 13988
rect 15764 13932 15792 13960
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 15746 13920 15752 13932
rect 15659 13892 15752 13920
rect 14921 13883 14979 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 16022 13920 16028 13932
rect 15983 13892 16028 13920
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 17052 13929 17080 13960
rect 17218 13948 17224 14000
rect 17276 13988 17282 14000
rect 19334 13988 19340 14000
rect 17276 13960 19340 13988
rect 17276 13948 17282 13960
rect 19334 13948 19340 13960
rect 19392 13988 19398 14000
rect 22002 13988 22008 14000
rect 19392 13960 22008 13988
rect 19392 13948 19398 13960
rect 22002 13948 22008 13960
rect 22060 13948 22066 14000
rect 30300 13997 30328 14028
rect 31754 14016 31760 14028
rect 31812 14016 31818 14068
rect 33965 14059 34023 14065
rect 33965 14025 33977 14059
rect 34011 14056 34023 14059
rect 34422 14056 34428 14068
rect 34011 14028 34284 14056
rect 34383 14028 34428 14056
rect 34011 14025 34023 14028
rect 33965 14019 34023 14025
rect 25869 13991 25927 13997
rect 25869 13957 25881 13991
rect 25915 13988 25927 13991
rect 30285 13991 30343 13997
rect 30285 13988 30297 13991
rect 25915 13960 30297 13988
rect 25915 13957 25927 13960
rect 25869 13951 25927 13957
rect 30285 13957 30297 13960
rect 30331 13957 30343 13991
rect 33137 13991 33195 13997
rect 33137 13988 33149 13991
rect 30285 13951 30343 13957
rect 30392 13960 33149 13988
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 16172 13892 16773 13920
rect 16172 13880 16178 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17126 13920 17132 13932
rect 17083 13892 17132 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 17954 13920 17960 13932
rect 17736 13892 17960 13920
rect 17736 13880 17742 13892
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 25958 13920 25964 13932
rect 19484 13892 25964 13920
rect 19484 13880 19490 13892
rect 25958 13880 25964 13892
rect 26016 13880 26022 13932
rect 26050 13880 26056 13932
rect 26108 13920 26114 13932
rect 29178 13920 29184 13932
rect 26108 13892 26153 13920
rect 29139 13892 29184 13920
rect 26108 13880 26114 13892
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 30190 13880 30196 13932
rect 30248 13920 30254 13932
rect 30392 13920 30420 13960
rect 33137 13957 33149 13960
rect 33183 13988 33195 13991
rect 34057 13991 34115 13997
rect 34057 13988 34069 13991
rect 33183 13960 34069 13988
rect 33183 13957 33195 13960
rect 33137 13951 33195 13957
rect 34057 13957 34069 13960
rect 34103 13957 34115 13991
rect 34256 13988 34284 14028
rect 34422 14016 34428 14028
rect 34480 14016 34486 14068
rect 36078 14056 36084 14068
rect 34716 14028 36084 14056
rect 34716 13988 34744 14028
rect 36078 14016 36084 14028
rect 36136 14056 36142 14068
rect 36265 14059 36323 14065
rect 36265 14056 36277 14059
rect 36136 14028 36277 14056
rect 36136 14016 36142 14028
rect 36265 14025 36277 14028
rect 36311 14056 36323 14059
rect 37090 14056 37096 14068
rect 36311 14028 37096 14056
rect 36311 14025 36323 14028
rect 36265 14019 36323 14025
rect 37090 14016 37096 14028
rect 37148 14016 37154 14068
rect 34256 13960 34744 13988
rect 34057 13951 34115 13957
rect 34790 13948 34796 14000
rect 34848 13988 34854 14000
rect 35130 13991 35188 13997
rect 35130 13988 35142 13991
rect 34848 13960 35142 13988
rect 34848 13948 34854 13960
rect 35130 13957 35142 13960
rect 35176 13957 35188 13991
rect 35130 13951 35188 13957
rect 30248 13892 30420 13920
rect 30248 13880 30254 13892
rect 30558 13880 30564 13932
rect 30616 13920 30622 13932
rect 31205 13923 31263 13929
rect 31205 13920 31217 13923
rect 30616 13892 31217 13920
rect 30616 13880 30622 13892
rect 31205 13889 31217 13892
rect 31251 13889 31263 13923
rect 31205 13883 31263 13889
rect 34146 13880 34152 13932
rect 34204 13920 34210 13932
rect 34885 13923 34943 13929
rect 34885 13920 34897 13923
rect 34204 13892 34897 13920
rect 34204 13880 34210 13892
rect 34885 13889 34897 13892
rect 34931 13889 34943 13923
rect 34885 13883 34943 13889
rect 35894 13880 35900 13932
rect 35952 13920 35958 13932
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 35952 13892 37841 13920
rect 35952 13880 35958 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13262 13852 13268 13864
rect 13219 13824 13268 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15378 13852 15384 13864
rect 14875 13824 15384 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 16850 13852 16856 13864
rect 16040 13824 16856 13852
rect 16040 13796 16068 13824
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17862 13852 17868 13864
rect 17823 13824 17868 13852
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 20772 13824 25697 13852
rect 20772 13812 20778 13824
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 30469 13855 30527 13861
rect 30469 13821 30481 13855
rect 30515 13821 30527 13855
rect 30469 13815 30527 13821
rect 33873 13855 33931 13861
rect 33873 13821 33885 13855
rect 33919 13821 33931 13855
rect 33873 13815 33931 13821
rect 9401 13787 9459 13793
rect 9401 13784 9413 13787
rect 8588 13756 9413 13784
rect 9401 13753 9413 13756
rect 9447 13753 9459 13787
rect 15562 13784 15568 13796
rect 9401 13747 9459 13753
rect 14936 13756 15568 13784
rect 2498 13716 2504 13728
rect 2459 13688 2504 13716
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 2961 13719 3019 13725
rect 2961 13685 2973 13719
rect 3007 13716 3019 13719
rect 4062 13716 4068 13728
rect 3007 13688 4068 13716
rect 3007 13685 3019 13688
rect 2961 13679 3019 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 10413 13719 10471 13725
rect 10413 13685 10425 13719
rect 10459 13716 10471 13719
rect 10686 13716 10692 13728
rect 10459 13688 10692 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 14936 13725 14964 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 15838 13784 15844 13796
rect 15751 13756 15844 13784
rect 14921 13719 14979 13725
rect 14921 13685 14933 13719
rect 14967 13685 14979 13719
rect 14921 13679 14979 13685
rect 15105 13719 15163 13725
rect 15105 13685 15117 13719
rect 15151 13716 15163 13719
rect 15378 13716 15384 13728
rect 15151 13688 15384 13716
rect 15151 13685 15163 13688
rect 15105 13679 15163 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 15764 13716 15792 13756
rect 15838 13744 15844 13756
rect 15896 13744 15902 13796
rect 15933 13787 15991 13793
rect 15933 13753 15945 13787
rect 15979 13784 15991 13787
rect 16022 13784 16028 13796
rect 15979 13756 16028 13784
rect 15979 13753 15991 13756
rect 15933 13747 15991 13753
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 16945 13787 17003 13793
rect 16945 13753 16957 13787
rect 16991 13753 17003 13787
rect 16945 13747 17003 13753
rect 16960 13716 16988 13747
rect 17494 13744 17500 13796
rect 17552 13784 17558 13796
rect 20254 13784 20260 13796
rect 17552 13756 20260 13784
rect 17552 13744 17558 13756
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 21358 13744 21364 13796
rect 21416 13784 21422 13796
rect 21821 13787 21879 13793
rect 21821 13784 21833 13787
rect 21416 13756 21833 13784
rect 21416 13744 21422 13756
rect 21821 13753 21833 13756
rect 21867 13753 21879 13787
rect 21821 13747 21879 13753
rect 30374 13744 30380 13796
rect 30432 13784 30438 13796
rect 30484 13784 30512 13815
rect 30432 13756 30512 13784
rect 33888 13784 33916 13815
rect 34330 13784 34336 13796
rect 33888 13756 34336 13784
rect 30432 13744 30438 13756
rect 34330 13744 34336 13756
rect 34388 13744 34394 13796
rect 17218 13716 17224 13728
rect 15764 13688 16988 13716
rect 17179 13688 17224 13716
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 30926 13676 30932 13728
rect 30984 13716 30990 13728
rect 31021 13719 31079 13725
rect 31021 13716 31033 13719
rect 30984 13688 31033 13716
rect 30984 13676 30990 13688
rect 31021 13685 31033 13688
rect 31067 13685 31079 13719
rect 38010 13716 38016 13728
rect 37971 13688 38016 13716
rect 31021 13679 31079 13685
rect 38010 13676 38016 13688
rect 38068 13676 38074 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2774 13512 2780 13524
rect 2363 13484 2780 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 9582 13512 9588 13524
rect 9543 13484 9588 13512
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 10796 13484 12081 13512
rect 8389 13447 8447 13453
rect 8389 13413 8401 13447
rect 8435 13444 8447 13447
rect 10686 13444 10692 13456
rect 8435 13416 10692 13444
rect 8435 13413 8447 13416
rect 8389 13407 8447 13413
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 3694 13336 3700 13388
rect 3752 13376 3758 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 3752 13348 4261 13376
rect 3752 13336 3758 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 9490 13376 9496 13388
rect 4249 13339 4307 13345
rect 9140 13348 9496 13376
rect 9140 13320 9168 13348
rect 9490 13336 9496 13348
rect 9548 13376 9554 13388
rect 9548 13348 10364 13376
rect 9548 13336 9554 13348
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2130 13308 2136 13320
rect 2091 13280 2136 13308
rect 2130 13268 2136 13280
rect 2188 13308 2194 13320
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2188 13280 2789 13308
rect 2188 13268 2194 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 3786 13308 3792 13320
rect 3747 13280 3792 13308
rect 2777 13271 2835 13277
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 4062 13308 4068 13320
rect 4023 13280 4068 13308
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 7006 13308 7012 13320
rect 6967 13280 7012 13308
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8938 13308 8944 13320
rect 8899 13280 8944 13308
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9398 13308 9404 13320
rect 9359 13280 9404 13308
rect 9398 13268 9404 13280
rect 9456 13308 9462 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9456 13280 10241 13308
rect 9456 13268 9462 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10336 13308 10364 13348
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 10336 13280 10517 13308
rect 10229 13271 10287 13277
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10686 13308 10692 13320
rect 10647 13280 10692 13308
rect 10505 13271 10563 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 7276 13243 7334 13249
rect 7276 13209 7288 13243
rect 7322 13240 7334 13243
rect 7926 13240 7932 13252
rect 7322 13212 7932 13240
rect 7322 13209 7334 13212
rect 7276 13203 7334 13209
rect 7926 13200 7932 13212
rect 7984 13200 7990 13252
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 10045 13243 10103 13249
rect 10045 13240 10057 13243
rect 8168 13212 10057 13240
rect 8168 13200 8174 13212
rect 10045 13209 10057 13212
rect 10091 13209 10103 13243
rect 10045 13203 10103 13209
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 4341 13175 4399 13181
rect 4341 13141 4353 13175
rect 4387 13172 4399 13175
rect 10796 13172 10824 13484
rect 12069 13481 12081 13484
rect 12115 13512 12127 13515
rect 12250 13512 12256 13524
rect 12115 13484 12256 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 13872 13484 18705 13512
rect 13872 13472 13878 13484
rect 18693 13481 18705 13484
rect 18739 13512 18751 13515
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 18739 13484 19257 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 24670 13512 24676 13524
rect 20036 13484 24676 13512
rect 20036 13472 20042 13484
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 28534 13512 28540 13524
rect 28495 13484 28540 13512
rect 28534 13472 28540 13484
rect 28592 13472 28598 13524
rect 30193 13515 30251 13521
rect 30193 13481 30205 13515
rect 30239 13512 30251 13515
rect 30558 13512 30564 13524
rect 30239 13484 30564 13512
rect 30239 13481 30251 13484
rect 30193 13475 30251 13481
rect 30558 13472 30564 13484
rect 30616 13472 30622 13524
rect 32030 13512 32036 13524
rect 31943 13484 32036 13512
rect 32030 13472 32036 13484
rect 32088 13512 32094 13524
rect 35894 13512 35900 13524
rect 32088 13484 35900 13512
rect 32088 13472 32094 13484
rect 35894 13472 35900 13484
rect 35952 13472 35958 13524
rect 17126 13404 17132 13456
rect 17184 13444 17190 13456
rect 26513 13447 26571 13453
rect 26513 13444 26525 13447
rect 17184 13416 26525 13444
rect 17184 13404 17190 13416
rect 26513 13413 26525 13416
rect 26559 13413 26571 13447
rect 30006 13444 30012 13456
rect 29967 13416 30012 13444
rect 26513 13407 26571 13413
rect 30006 13404 30012 13416
rect 30064 13404 30070 13456
rect 34057 13447 34115 13453
rect 34057 13413 34069 13447
rect 34103 13444 34115 13447
rect 34701 13447 34759 13453
rect 34701 13444 34713 13447
rect 34103 13416 34713 13444
rect 34103 13413 34115 13416
rect 34057 13407 34115 13413
rect 34701 13413 34713 13416
rect 34747 13413 34759 13447
rect 34701 13407 34759 13413
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 14792 13348 15577 13376
rect 14792 13336 14798 13348
rect 15565 13345 15577 13348
rect 15611 13345 15623 13379
rect 15565 13339 15623 13345
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 15841 13379 15899 13385
rect 15841 13376 15853 13379
rect 15804 13348 15853 13376
rect 15804 13336 15810 13348
rect 15841 13345 15853 13348
rect 15887 13376 15899 13379
rect 15930 13376 15936 13388
rect 15887 13348 15936 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 17218 13376 17224 13388
rect 16899 13348 17224 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 20714 13376 20720 13388
rect 17327 13348 20720 13376
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 12986 13308 12992 13320
rect 12943 13280 12992 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13265 13311 13323 13317
rect 13136 13280 13181 13308
rect 13136 13268 13142 13280
rect 13265 13277 13277 13311
rect 13311 13308 13323 13311
rect 13354 13308 13360 13320
rect 13311 13280 13360 13308
rect 13311 13277 13323 13280
rect 13265 13271 13323 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 17327 13317 17355 13348
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 21637 13379 21695 13385
rect 21637 13376 21649 13379
rect 21008 13348 21649 13376
rect 21008 13320 21036 13348
rect 21637 13345 21649 13348
rect 21683 13345 21695 13379
rect 21637 13339 21695 13345
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 24728 13348 25237 13376
rect 24728 13336 24734 13348
rect 25225 13345 25237 13348
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 29733 13379 29791 13385
rect 29733 13345 29745 13379
rect 29779 13376 29791 13379
rect 30098 13376 30104 13388
rect 29779 13348 30104 13376
rect 29779 13345 29791 13348
rect 29733 13339 29791 13345
rect 30098 13336 30104 13348
rect 30156 13336 30162 13388
rect 34146 13336 34152 13388
rect 34204 13376 34210 13388
rect 34330 13376 34336 13388
rect 34204 13348 34336 13376
rect 34204 13336 34210 13348
rect 34330 13336 34336 13348
rect 34388 13376 34394 13388
rect 35253 13379 35311 13385
rect 35253 13376 35265 13379
rect 34388 13348 35265 13376
rect 34388 13336 34394 13348
rect 35253 13345 35265 13348
rect 35299 13345 35311 13379
rect 35253 13339 35311 13345
rect 37274 13336 37280 13388
rect 37332 13376 37338 13388
rect 37332 13348 37504 13376
rect 37332 13336 37338 13348
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 18966 13308 18972 13320
rect 18472 13280 18972 13308
rect 18472 13268 18478 13280
rect 18966 13268 18972 13280
rect 19024 13308 19030 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 19024 13280 19257 13308
rect 19024 13268 19030 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 20806 13308 20812 13320
rect 19392 13280 19437 13308
rect 20767 13280 20812 13308
rect 19392 13268 19398 13280
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 20990 13308 20996 13320
rect 20951 13280 20996 13308
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 13449 13243 13507 13249
rect 13449 13209 13461 13243
rect 13495 13240 13507 13243
rect 15102 13240 15108 13252
rect 13495 13212 15108 13240
rect 13495 13209 13507 13212
rect 13449 13203 13507 13209
rect 15102 13200 15108 13212
rect 15160 13200 15166 13252
rect 16666 13200 16672 13252
rect 16724 13240 16730 13252
rect 16991 13243 17049 13249
rect 16991 13240 17003 13243
rect 16724 13212 17003 13240
rect 16724 13200 16730 13212
rect 16991 13209 17003 13212
rect 17037 13209 17049 13243
rect 16991 13203 17049 13209
rect 17129 13243 17187 13249
rect 17129 13209 17141 13243
rect 17175 13209 17187 13243
rect 17129 13203 17187 13209
rect 17221 13243 17279 13249
rect 17221 13209 17233 13243
rect 17267 13240 17279 13243
rect 18049 13243 18107 13249
rect 18049 13240 18061 13243
rect 17267 13212 18061 13240
rect 17267 13209 17279 13212
rect 17221 13203 17279 13209
rect 18049 13209 18061 13212
rect 18095 13240 18107 13243
rect 19426 13240 19432 13252
rect 18095 13212 19432 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 11146 13172 11152 13184
rect 4387 13144 10824 13172
rect 11107 13144 11152 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 11146 13132 11152 13144
rect 11204 13172 11210 13184
rect 12069 13175 12127 13181
rect 12069 13172 12081 13175
rect 11204 13144 12081 13172
rect 11204 13132 11210 13144
rect 12069 13141 12081 13144
rect 12115 13141 12127 13175
rect 12069 13135 12127 13141
rect 12253 13175 12311 13181
rect 12253 13141 12265 13175
rect 12299 13172 12311 13175
rect 12526 13172 12532 13184
rect 12299 13144 12532 13172
rect 12299 13141 12311 13144
rect 12253 13135 12311 13141
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 14185 13175 14243 13181
rect 14185 13141 14197 13175
rect 14231 13172 14243 13175
rect 14274 13172 14280 13184
rect 14231 13144 14280 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 17144 13172 17172 13203
rect 19426 13200 19432 13212
rect 19484 13200 19490 13252
rect 20073 13243 20131 13249
rect 20073 13240 20085 13243
rect 19536 13212 20085 13240
rect 17310 13172 17316 13184
rect 16908 13144 17316 13172
rect 16908 13132 16914 13144
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 17494 13172 17500 13184
rect 17455 13144 17500 13172
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19536 13172 19564 13212
rect 20073 13209 20085 13212
rect 20119 13240 20131 13243
rect 21100 13240 21128 13271
rect 21358 13268 21364 13320
rect 21416 13308 21422 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21416 13280 21557 13308
rect 21416 13268 21422 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21818 13308 21824 13320
rect 21779 13280 21824 13308
rect 21545 13271 21603 13277
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 25317 13311 25375 13317
rect 25317 13308 25329 13311
rect 24820 13280 25329 13308
rect 24820 13268 24826 13280
rect 25317 13277 25329 13280
rect 25363 13277 25375 13311
rect 25317 13271 25375 13277
rect 25501 13311 25559 13317
rect 25501 13277 25513 13311
rect 25547 13308 25559 13311
rect 25590 13308 25596 13320
rect 25547 13280 25596 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 25685 13311 25743 13317
rect 25685 13277 25697 13311
rect 25731 13308 25743 13311
rect 26510 13308 26516 13320
rect 25731 13280 26516 13308
rect 25731 13277 25743 13280
rect 25685 13271 25743 13277
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 29546 13268 29552 13320
rect 29604 13308 29610 13320
rect 30282 13308 30288 13320
rect 29604 13280 30288 13308
rect 29604 13268 29610 13280
rect 30282 13268 30288 13280
rect 30340 13308 30346 13320
rect 30926 13317 30932 13320
rect 30653 13311 30711 13317
rect 30653 13308 30665 13311
rect 30340 13280 30665 13308
rect 30340 13268 30346 13280
rect 30653 13277 30665 13280
rect 30699 13277 30711 13311
rect 30920 13308 30932 13317
rect 30887 13280 30932 13308
rect 30653 13271 30711 13277
rect 30920 13271 30932 13280
rect 30926 13268 30932 13271
rect 30984 13268 30990 13320
rect 31202 13268 31208 13320
rect 31260 13308 31266 13320
rect 36998 13317 37004 13320
rect 35069 13311 35127 13317
rect 35069 13308 35081 13311
rect 31260 13280 35081 13308
rect 31260 13268 31266 13280
rect 35069 13277 35081 13280
rect 35115 13308 35127 13311
rect 35897 13311 35955 13317
rect 35897 13308 35909 13311
rect 35115 13280 35909 13308
rect 35115 13277 35127 13280
rect 35069 13271 35127 13277
rect 35897 13277 35909 13280
rect 35943 13277 35955 13311
rect 36996 13308 37004 13317
rect 36959 13280 37004 13308
rect 35897 13271 35955 13277
rect 36996 13271 37004 13280
rect 36998 13268 37004 13271
rect 37056 13268 37062 13320
rect 37182 13308 37188 13320
rect 37143 13280 37188 13308
rect 37182 13268 37188 13280
rect 37240 13268 37246 13320
rect 37476 13317 37504 13348
rect 37368 13311 37426 13317
rect 37368 13277 37380 13311
rect 37414 13277 37426 13311
rect 37368 13271 37426 13277
rect 37461 13311 37519 13317
rect 37461 13277 37473 13311
rect 37507 13277 37519 13311
rect 38102 13308 38108 13320
rect 38063 13280 38108 13308
rect 37461 13271 37519 13277
rect 20119 13212 21128 13240
rect 20119 13209 20131 13212
rect 20073 13203 20131 13209
rect 26050 13200 26056 13252
rect 26108 13240 26114 13252
rect 26145 13243 26203 13249
rect 26145 13240 26157 13243
rect 26108 13212 26157 13240
rect 26108 13200 26114 13212
rect 26145 13209 26157 13212
rect 26191 13209 26203 13243
rect 26145 13203 26203 13209
rect 26329 13243 26387 13249
rect 26329 13209 26341 13243
rect 26375 13240 26387 13243
rect 29638 13240 29644 13252
rect 26375 13212 29644 13240
rect 26375 13209 26387 13212
rect 26329 13203 26387 13209
rect 29638 13200 29644 13212
rect 29696 13200 29702 13252
rect 33689 13243 33747 13249
rect 33689 13209 33701 13243
rect 33735 13240 33747 13243
rect 34238 13240 34244 13252
rect 33735 13212 34244 13240
rect 33735 13209 33747 13212
rect 33689 13203 33747 13209
rect 34238 13200 34244 13212
rect 34296 13200 34302 13252
rect 35161 13243 35219 13249
rect 35161 13209 35173 13243
rect 35207 13240 35219 13243
rect 35986 13240 35992 13252
rect 35207 13212 35992 13240
rect 35207 13209 35219 13212
rect 35161 13203 35219 13209
rect 35986 13200 35992 13212
rect 36044 13240 36050 13252
rect 37093 13243 37151 13249
rect 37093 13240 37105 13243
rect 36044 13212 37105 13240
rect 36044 13200 36050 13212
rect 36924 13184 36952 13212
rect 37093 13209 37105 13212
rect 37139 13209 37151 13243
rect 37384 13240 37412 13271
rect 38102 13268 38108 13280
rect 38160 13268 38166 13320
rect 37384 13212 37964 13240
rect 37093 13203 37151 13209
rect 18932 13144 19564 13172
rect 19613 13175 19671 13181
rect 18932 13132 18938 13144
rect 19613 13141 19625 13175
rect 19659 13172 19671 13175
rect 19978 13172 19984 13184
rect 19659 13144 19984 13172
rect 19659 13141 19671 13144
rect 19613 13135 19671 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20622 13172 20628 13184
rect 20583 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 22005 13175 22063 13181
rect 22005 13141 22017 13175
rect 22051 13172 22063 13175
rect 22094 13172 22100 13184
rect 22051 13144 22100 13172
rect 22051 13141 22063 13144
rect 22005 13135 22063 13141
rect 22094 13132 22100 13144
rect 22152 13132 22158 13184
rect 22554 13172 22560 13184
rect 22467 13144 22560 13172
rect 22554 13132 22560 13144
rect 22612 13172 22618 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 22612 13144 23857 13172
rect 22612 13132 22618 13144
rect 23845 13141 23857 13144
rect 23891 13172 23903 13175
rect 24026 13172 24032 13184
rect 23891 13144 24032 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 34149 13175 34207 13181
rect 34149 13141 34161 13175
rect 34195 13172 34207 13175
rect 34974 13172 34980 13184
rect 34195 13144 34980 13172
rect 34195 13141 34207 13144
rect 34149 13135 34207 13141
rect 34974 13132 34980 13144
rect 35032 13132 35038 13184
rect 36814 13172 36820 13184
rect 36775 13144 36820 13172
rect 36814 13132 36820 13144
rect 36872 13132 36878 13184
rect 36906 13132 36912 13184
rect 36964 13132 36970 13184
rect 37936 13181 37964 13212
rect 37921 13175 37979 13181
rect 37921 13141 37933 13175
rect 37967 13141 37979 13175
rect 37921 13135 37979 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 6546 12968 6552 12980
rect 4203 12940 6552 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 11146 12968 11152 12980
rect 8076 12940 11152 12968
rect 8076 12928 8082 12940
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 12069 12971 12127 12977
rect 12069 12968 12081 12971
rect 11756 12940 12081 12968
rect 11756 12928 11762 12940
rect 12069 12937 12081 12940
rect 12115 12968 12127 12971
rect 13633 12971 13691 12977
rect 12115 12940 13584 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 2225 12903 2283 12909
rect 2225 12869 2237 12903
rect 2271 12900 2283 12903
rect 6914 12900 6920 12912
rect 2271 12872 6920 12900
rect 2271 12869 2283 12872
rect 2225 12863 2283 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 13078 12900 13084 12912
rect 12406 12872 13084 12900
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12832 1918 12844
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 1912 12804 2697 12832
rect 1912 12792 1918 12804
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 3510 12832 3516 12844
rect 3471 12804 3516 12832
rect 2685 12795 2743 12801
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 3694 12841 3700 12844
rect 3660 12835 3700 12841
rect 3660 12801 3672 12835
rect 3660 12795 3700 12801
rect 3694 12792 3700 12795
rect 3752 12792 3758 12844
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7064 12804 7757 12832
rect 7064 12792 7070 12804
rect 7745 12801 7757 12804
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 8012 12835 8070 12841
rect 8012 12801 8024 12835
rect 8058 12832 8070 12835
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 8058 12804 9597 12832
rect 8058 12801 8070 12804
rect 8012 12795 8070 12801
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 9766 12832 9772 12844
rect 9727 12804 9772 12832
rect 9585 12795 9643 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9916 12804 9965 12832
rect 9916 12792 9922 12804
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 12406 12832 12434 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 13556 12900 13584 12940
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13814 12968 13820 12980
rect 13679 12940 13820 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13814 12928 13820 12940
rect 13872 12968 13878 12980
rect 13998 12968 14004 12980
rect 13872 12940 14004 12968
rect 13872 12928 13878 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 27065 12971 27123 12977
rect 27065 12937 27077 12971
rect 27111 12968 27123 12971
rect 27154 12968 27160 12980
rect 27111 12940 27160 12968
rect 27111 12937 27123 12940
rect 27065 12931 27123 12937
rect 14274 12900 14280 12912
rect 13556 12872 14280 12900
rect 14274 12860 14280 12872
rect 14332 12900 14338 12912
rect 20254 12900 20260 12912
rect 14332 12872 18644 12900
rect 14332 12860 14338 12872
rect 12710 12832 12716 12844
rect 12299 12804 12434 12832
rect 12671 12804 12716 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 12710 12792 12716 12804
rect 12768 12832 12774 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 12768 12804 13461 12832
rect 12768 12792 12774 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13688 12804 14381 12832
rect 13688 12792 13694 12804
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15436 12804 15669 12832
rect 15436 12792 15442 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15838 12832 15844 12844
rect 15799 12804 15844 12832
rect 15657 12795 15715 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 16807 12835 16865 12841
rect 15988 12804 16033 12832
rect 15988 12792 15994 12804
rect 16807 12801 16819 12835
rect 16853 12801 16865 12835
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16807 12795 16865 12801
rect 3418 12724 3424 12776
rect 3476 12764 3482 12776
rect 3786 12764 3792 12776
rect 3476 12736 3792 12764
rect 3476 12724 3482 12736
rect 3786 12724 3792 12736
rect 3844 12764 3850 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3844 12736 3893 12764
rect 3844 12724 3850 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9732 12736 10057 12764
rect 9732 12724 9738 12736
rect 10045 12733 10057 12736
rect 10091 12764 10103 12767
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10091 12736 10517 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 13648 12764 13676 12792
rect 12676 12736 13676 12764
rect 15749 12767 15807 12773
rect 12676 12724 12682 12736
rect 15749 12733 15761 12767
rect 15795 12764 15807 12767
rect 16022 12764 16028 12776
rect 15795 12736 16028 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 16022 12724 16028 12736
rect 16080 12724 16086 12776
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16669 12767 16727 12773
rect 16669 12764 16681 12767
rect 16163 12736 16681 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16669 12733 16681 12736
rect 16715 12733 16727 12767
rect 16669 12727 16727 12733
rect 4062 12696 4068 12708
rect 3804 12668 4068 12696
rect 3804 12637 3832 12668
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 12897 12699 12955 12705
rect 12897 12665 12909 12699
rect 12943 12696 12955 12699
rect 13354 12696 13360 12708
rect 12943 12668 13360 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 13354 12656 13360 12668
rect 13412 12696 13418 12708
rect 16822 12696 16850 12795
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17052 12764 17080 12795
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17184 12804 17229 12832
rect 17184 12792 17190 12804
rect 18616 12776 18644 12872
rect 19904 12872 20260 12900
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 19904 12841 19932 12872
rect 20254 12860 20260 12872
rect 20312 12900 20318 12912
rect 22554 12900 22560 12912
rect 20312 12872 22560 12900
rect 20312 12860 20318 12872
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19852 12804 19901 12832
rect 19852 12792 19858 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 20156 12835 20214 12841
rect 20156 12801 20168 12835
rect 20202 12832 20214 12835
rect 20622 12832 20628 12844
rect 20202 12804 20628 12832
rect 20202 12801 20214 12804
rect 20156 12795 20214 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21836 12841 21864 12872
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 24762 12860 24768 12912
rect 24820 12900 24826 12912
rect 24820 12872 26280 12900
rect 24820 12860 24826 12872
rect 22094 12841 22100 12844
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 22088 12795 22100 12841
rect 22152 12832 22158 12844
rect 24302 12841 24308 12844
rect 22152 12804 22188 12832
rect 22094 12792 22100 12795
rect 22152 12792 22158 12804
rect 24296 12795 24308 12841
rect 24360 12832 24366 12844
rect 26053 12835 26111 12841
rect 24360 12804 24396 12832
rect 24302 12792 24308 12795
rect 24360 12792 24366 12804
rect 26053 12801 26065 12835
rect 26099 12832 26111 12835
rect 26142 12832 26148 12844
rect 26099 12804 26148 12832
rect 26099 12801 26111 12804
rect 26053 12795 26111 12801
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 26252 12841 26280 12872
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12832 26387 12835
rect 27080 12832 27108 12931
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 30006 12968 30012 12980
rect 29967 12940 30012 12968
rect 30006 12928 30012 12940
rect 30064 12928 30070 12980
rect 30377 12971 30435 12977
rect 30377 12937 30389 12971
rect 30423 12968 30435 12971
rect 30466 12968 30472 12980
rect 30423 12940 30472 12968
rect 30423 12937 30435 12940
rect 30377 12931 30435 12937
rect 30466 12928 30472 12940
rect 30524 12968 30530 12980
rect 31202 12968 31208 12980
rect 30524 12940 31208 12968
rect 30524 12928 30530 12940
rect 31202 12928 31208 12940
rect 31260 12928 31266 12980
rect 32030 12968 32036 12980
rect 31726 12940 32036 12968
rect 29454 12860 29460 12912
rect 29512 12900 29518 12912
rect 31297 12903 31355 12909
rect 31297 12900 31309 12903
rect 29512 12872 31309 12900
rect 29512 12860 29518 12872
rect 31297 12869 31309 12872
rect 31343 12869 31355 12903
rect 31297 12863 31355 12869
rect 26375 12804 27108 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 28534 12792 28540 12844
rect 28592 12832 28598 12844
rect 28813 12835 28871 12841
rect 28813 12832 28825 12835
rect 28592 12804 28825 12832
rect 28592 12792 28598 12804
rect 28813 12801 28825 12804
rect 28859 12801 28871 12835
rect 28813 12795 28871 12801
rect 28997 12835 29055 12841
rect 28997 12801 29009 12835
rect 29043 12832 29055 12835
rect 29086 12832 29092 12844
rect 29043 12804 29092 12832
rect 29043 12801 29055 12804
rect 28997 12795 29055 12801
rect 29086 12792 29092 12804
rect 29144 12792 29150 12844
rect 29638 12792 29644 12844
rect 29696 12832 29702 12844
rect 30469 12835 30527 12841
rect 30469 12832 30481 12835
rect 29696 12804 30481 12832
rect 29696 12792 29702 12804
rect 30469 12801 30481 12804
rect 30515 12832 30527 12835
rect 31726 12832 31754 12940
rect 32030 12928 32036 12940
rect 32088 12928 32094 12980
rect 37369 12971 37427 12977
rect 37369 12937 37381 12971
rect 37415 12968 37427 12971
rect 38102 12968 38108 12980
rect 37415 12940 38108 12968
rect 37415 12937 37427 12940
rect 37369 12931 37427 12937
rect 38102 12928 38108 12940
rect 38160 12928 38166 12980
rect 30515 12804 31754 12832
rect 30515 12801 30527 12804
rect 30469 12795 30527 12801
rect 33502 12792 33508 12844
rect 33560 12832 33566 12844
rect 33597 12835 33655 12841
rect 33597 12832 33609 12835
rect 33560 12804 33609 12832
rect 33560 12792 33566 12804
rect 33597 12801 33609 12804
rect 33643 12832 33655 12835
rect 34425 12835 34483 12841
rect 34425 12832 34437 12835
rect 33643 12804 34437 12832
rect 33643 12801 33655 12804
rect 33597 12795 33655 12801
rect 34425 12801 34437 12804
rect 34471 12801 34483 12835
rect 34425 12795 34483 12801
rect 34974 12792 34980 12844
rect 35032 12832 35038 12844
rect 35529 12835 35587 12841
rect 35529 12832 35541 12835
rect 35032 12804 35541 12832
rect 35032 12792 35038 12804
rect 35529 12801 35541 12804
rect 35575 12801 35587 12835
rect 35529 12795 35587 12801
rect 37829 12835 37887 12841
rect 37829 12801 37841 12835
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 17862 12764 17868 12776
rect 17052 12736 17868 12764
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18656 12736 18705 12764
rect 18656 12724 18662 12736
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 24026 12764 24032 12776
rect 23987 12736 24032 12764
rect 18693 12727 18751 12733
rect 24026 12724 24032 12736
rect 24084 12724 24090 12776
rect 28166 12724 28172 12776
rect 28224 12764 28230 12776
rect 28261 12767 28319 12773
rect 28261 12764 28273 12767
rect 28224 12736 28273 12764
rect 28224 12724 28230 12736
rect 28261 12733 28273 12736
rect 28307 12764 28319 12767
rect 28721 12767 28779 12773
rect 28721 12764 28733 12767
rect 28307 12736 28733 12764
rect 28307 12733 28319 12736
rect 28261 12727 28319 12733
rect 28721 12733 28733 12736
rect 28767 12733 28779 12767
rect 28721 12727 28779 12733
rect 30374 12724 30380 12776
rect 30432 12764 30438 12776
rect 30561 12767 30619 12773
rect 30561 12764 30573 12767
rect 30432 12736 30573 12764
rect 30432 12724 30438 12736
rect 30561 12733 30573 12736
rect 30607 12733 30619 12767
rect 34146 12764 34152 12776
rect 34107 12736 34152 12764
rect 30561 12727 30619 12733
rect 34146 12724 34152 12736
rect 34204 12724 34210 12776
rect 34333 12767 34391 12773
rect 34333 12733 34345 12767
rect 34379 12764 34391 12767
rect 37182 12764 37188 12776
rect 34379 12736 37188 12764
rect 34379 12733 34391 12736
rect 34333 12727 34391 12733
rect 37182 12724 37188 12736
rect 37240 12764 37246 12776
rect 37844 12764 37872 12795
rect 37240 12736 37872 12764
rect 37240 12724 37246 12736
rect 17034 12696 17040 12708
rect 13412 12668 15976 12696
rect 16822 12668 17040 12696
rect 13412 12656 13418 12668
rect 3789 12631 3847 12637
rect 3789 12597 3801 12631
rect 3835 12597 3847 12631
rect 3789 12591 3847 12597
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 8996 12600 9137 12628
rect 8996 12588 9002 12600
rect 9125 12597 9137 12600
rect 9171 12597 9183 12631
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 9125 12591 9183 12597
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 15948 12628 15976 12668
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 18874 12696 18880 12708
rect 17236 12668 18880 12696
rect 17236 12628 17264 12668
rect 18874 12656 18880 12668
rect 18932 12656 18938 12708
rect 15948 12600 17264 12628
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12628 17371 12631
rect 17402 12628 17408 12640
rect 17359 12600 17408 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18969 12631 19027 12637
rect 18969 12597 18981 12631
rect 19015 12628 19027 12631
rect 19334 12628 19340 12640
rect 19015 12600 19340 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 20898 12588 20904 12640
rect 20956 12628 20962 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20956 12600 21281 12628
rect 20956 12588 20962 12600
rect 21269 12597 21281 12600
rect 21315 12597 21327 12631
rect 21269 12591 21327 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 23201 12631 23259 12637
rect 23201 12628 23213 12631
rect 22520 12600 23213 12628
rect 22520 12588 22526 12600
rect 23201 12597 23213 12600
rect 23247 12597 23259 12631
rect 23201 12591 23259 12597
rect 25038 12588 25044 12640
rect 25096 12628 25102 12640
rect 25409 12631 25467 12637
rect 25409 12628 25421 12631
rect 25096 12600 25421 12628
rect 25096 12588 25102 12600
rect 25409 12597 25421 12600
rect 25455 12597 25467 12631
rect 25409 12591 25467 12597
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 25869 12631 25927 12637
rect 25869 12628 25881 12631
rect 25740 12600 25881 12628
rect 25740 12588 25746 12600
rect 25869 12597 25881 12600
rect 25915 12597 25927 12631
rect 25869 12591 25927 12597
rect 29181 12631 29239 12637
rect 29181 12597 29193 12631
rect 29227 12628 29239 12631
rect 29638 12628 29644 12640
rect 29227 12600 29644 12628
rect 29227 12597 29239 12600
rect 29181 12591 29239 12597
rect 29638 12588 29644 12600
rect 29696 12588 29702 12640
rect 31386 12628 31392 12640
rect 31347 12600 31392 12628
rect 31386 12588 31392 12600
rect 31444 12588 31450 12640
rect 34790 12628 34796 12640
rect 34751 12600 34796 12628
rect 34790 12588 34796 12600
rect 34848 12588 34854 12640
rect 35710 12628 35716 12640
rect 35671 12600 35716 12628
rect 35710 12588 35716 12600
rect 35768 12588 35774 12640
rect 38010 12628 38016 12640
rect 37971 12600 38016 12628
rect 38010 12588 38016 12600
rect 38068 12588 38074 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 2498 12424 2504 12436
rect 1627 12396 2504 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 4062 12424 4068 12436
rect 4023 12396 4068 12424
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 7282 12424 7288 12436
rect 4479 12396 7288 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 9585 12427 9643 12433
rect 9585 12393 9597 12427
rect 9631 12424 9643 12427
rect 9766 12424 9772 12436
rect 9631 12396 9772 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 16482 12424 16488 12436
rect 16395 12396 16488 12424
rect 16482 12384 16488 12396
rect 16540 12424 16546 12436
rect 16758 12424 16764 12436
rect 16540 12396 16764 12424
rect 16540 12384 16546 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 19794 12424 19800 12436
rect 19755 12396 19800 12424
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 20254 12384 20260 12436
rect 20312 12424 20318 12436
rect 20714 12424 20720 12436
rect 20312 12396 20720 12424
rect 20312 12384 20318 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 20806 12384 20812 12436
rect 20864 12424 20870 12436
rect 21729 12427 21787 12433
rect 21729 12424 21741 12427
rect 20864 12396 21741 12424
rect 20864 12384 20870 12396
rect 21729 12393 21741 12396
rect 21775 12393 21787 12427
rect 21729 12387 21787 12393
rect 24302 12384 24308 12436
rect 24360 12424 24366 12436
rect 24397 12427 24455 12433
rect 24397 12424 24409 12427
rect 24360 12396 24409 12424
rect 24360 12384 24366 12396
rect 24397 12393 24409 12396
rect 24443 12393 24455 12427
rect 24397 12387 24455 12393
rect 24670 12384 24676 12436
rect 24728 12424 24734 12436
rect 28629 12427 28687 12433
rect 28629 12424 28641 12427
rect 24728 12396 28641 12424
rect 24728 12384 24734 12396
rect 28629 12393 28641 12396
rect 28675 12393 28687 12427
rect 28629 12387 28687 12393
rect 36906 12384 36912 12436
rect 36964 12424 36970 12436
rect 37553 12427 37611 12433
rect 37553 12424 37565 12427
rect 36964 12396 37565 12424
rect 36964 12384 36970 12396
rect 37553 12393 37565 12396
rect 37599 12393 37611 12427
rect 37553 12387 37611 12393
rect 3694 12316 3700 12368
rect 3752 12356 3758 12368
rect 3927 12359 3985 12365
rect 3927 12356 3939 12359
rect 3752 12328 3939 12356
rect 3752 12316 3758 12328
rect 3927 12325 3939 12328
rect 3973 12325 3985 12359
rect 3927 12319 3985 12325
rect 8297 12359 8355 12365
rect 8297 12325 8309 12359
rect 8343 12356 8355 12359
rect 9858 12356 9864 12368
rect 8343 12328 9864 12356
rect 8343 12325 8355 12328
rect 8297 12319 8355 12325
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 17494 12356 17500 12368
rect 9968 12328 17500 12356
rect 3145 12291 3203 12297
rect 3145 12257 3157 12291
rect 3191 12288 3203 12291
rect 4157 12291 4215 12297
rect 4157 12288 4169 12291
rect 3191 12260 4169 12288
rect 3191 12257 3203 12260
rect 3145 12251 3203 12257
rect 4157 12257 4169 12260
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 9968 12288 9996 12328
rect 17494 12316 17500 12328
rect 17552 12316 17558 12368
rect 24762 12356 24768 12368
rect 21008 12328 24768 12356
rect 21008 12300 21036 12328
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 34790 12356 34796 12368
rect 34751 12328 34796 12356
rect 34790 12316 34796 12328
rect 34848 12316 34854 12368
rect 13449 12291 13507 12297
rect 7524 12260 9996 12288
rect 12406 12260 13400 12288
rect 7524 12248 7530 12260
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12220 1458 12232
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1452 12192 2053 12220
rect 1452 12180 1458 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 2041 12183 2099 12189
rect 3050 12180 3056 12192
rect 3108 12220 3114 12232
rect 3418 12220 3424 12232
rect 3108 12192 3424 12220
rect 3108 12180 3114 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 8389 12183 8447 12189
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3568 12124 3801 12152
rect 3568 12112 3574 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 8404 12152 8432 12183
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9398 12220 9404 12232
rect 9272 12192 9404 12220
rect 9272 12180 9278 12192
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 12406 12152 12434 12260
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 13044 12192 13185 12220
rect 13044 12180 13050 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13372 12220 13400 12260
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 13538 12288 13544 12300
rect 13495 12260 13544 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 20990 12288 20996 12300
rect 20763 12260 20996 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 21192 12260 22416 12288
rect 16758 12220 16764 12232
rect 13372 12192 16764 12220
rect 13173 12183 13231 12189
rect 16758 12180 16764 12192
rect 16816 12220 16822 12232
rect 17770 12220 17776 12232
rect 16816 12192 17776 12220
rect 16816 12180 16822 12192
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 20036 12192 20453 12220
rect 20036 12180 20042 12192
rect 20441 12189 20453 12192
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 20898 12180 20904 12232
rect 20956 12220 20962 12232
rect 21192 12220 21220 12260
rect 20956 12192 21220 12220
rect 21913 12223 21971 12229
rect 20956 12180 20962 12192
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22002 12220 22008 12232
rect 21959 12192 22008 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12220 22247 12223
rect 22278 12220 22284 12232
rect 22235 12192 22284 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22388 12229 22416 12260
rect 24026 12248 24032 12300
rect 24084 12288 24090 12300
rect 25406 12288 25412 12300
rect 24084 12260 25412 12288
rect 24084 12248 24090 12260
rect 25406 12248 25412 12260
rect 25464 12248 25470 12300
rect 34701 12291 34759 12297
rect 34701 12288 34713 12291
rect 33980 12260 34713 12288
rect 22373 12223 22431 12229
rect 22373 12189 22385 12223
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 24394 12180 24400 12232
rect 24452 12220 24458 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24452 12192 24593 12220
rect 24452 12180 24458 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24857 12223 24915 12229
rect 24857 12189 24869 12223
rect 24903 12220 24915 12223
rect 25314 12220 25320 12232
rect 24903 12192 25320 12220
rect 24903 12189 24915 12192
rect 24857 12183 24915 12189
rect 3789 12115 3847 12121
rect 7392 12124 12434 12152
rect 7392 12096 7420 12124
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 16393 12155 16451 12161
rect 16393 12152 16405 12155
rect 15160 12124 16405 12152
rect 15160 12112 15166 12124
rect 16393 12121 16405 12124
rect 16439 12121 16451 12155
rect 16393 12115 16451 12121
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24872 12152 24900 12183
rect 25314 12180 25320 12192
rect 25372 12180 25378 12232
rect 25682 12229 25688 12232
rect 25676 12183 25688 12229
rect 25740 12220 25746 12232
rect 27249 12223 27307 12229
rect 25740 12192 25776 12220
rect 25682 12180 25688 12183
rect 25740 12180 25746 12192
rect 27249 12189 27261 12223
rect 27295 12220 27307 12223
rect 29546 12220 29552 12232
rect 27295 12192 29552 12220
rect 27295 12189 27307 12192
rect 27249 12183 27307 12189
rect 29546 12180 29552 12192
rect 29604 12180 29610 12232
rect 29638 12180 29644 12232
rect 29696 12220 29702 12232
rect 33980 12229 34008 12260
rect 34701 12257 34713 12260
rect 34747 12257 34759 12291
rect 34701 12251 34759 12257
rect 29805 12223 29863 12229
rect 29805 12220 29817 12223
rect 29696 12192 29817 12220
rect 29696 12180 29702 12192
rect 29805 12189 29817 12192
rect 29851 12189 29863 12223
rect 29805 12183 29863 12189
rect 33965 12223 34023 12229
rect 33965 12189 33977 12223
rect 34011 12189 34023 12223
rect 33965 12183 34023 12189
rect 34054 12180 34060 12232
rect 34112 12220 34118 12232
rect 34422 12220 34428 12232
rect 34112 12192 34428 12220
rect 34112 12180 34118 12192
rect 34422 12180 34428 12192
rect 34480 12220 34486 12232
rect 35713 12223 35771 12229
rect 35713 12220 35725 12223
rect 34480 12192 35725 12220
rect 34480 12180 34486 12192
rect 35713 12189 35725 12192
rect 35759 12220 35771 12223
rect 36173 12223 36231 12229
rect 36173 12220 36185 12223
rect 35759 12192 36185 12220
rect 35759 12189 35771 12192
rect 35713 12183 35771 12189
rect 36173 12189 36185 12192
rect 36219 12220 36231 12223
rect 36262 12220 36268 12232
rect 36219 12192 36268 12220
rect 36219 12189 36231 12192
rect 36173 12183 36231 12189
rect 36262 12180 36268 12192
rect 36320 12180 36326 12232
rect 23891 12124 24900 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 7374 12084 7380 12096
rect 7335 12056 7380 12084
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 12710 12084 12716 12096
rect 7616 12056 12716 12084
rect 7616 12044 7622 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 16408 12084 16436 12115
rect 26510 12112 26516 12164
rect 26568 12152 26574 12164
rect 27494 12155 27552 12161
rect 27494 12152 27506 12155
rect 26568 12124 27506 12152
rect 26568 12112 26574 12124
rect 27494 12121 27506 12124
rect 27540 12121 27552 12155
rect 27494 12115 27552 12121
rect 34238 12112 34244 12164
rect 34296 12152 34302 12164
rect 35161 12155 35219 12161
rect 35161 12152 35173 12155
rect 34296 12124 35173 12152
rect 34296 12112 34302 12124
rect 35161 12121 35173 12124
rect 35207 12121 35219 12155
rect 35161 12115 35219 12121
rect 35802 12112 35808 12164
rect 35860 12152 35866 12164
rect 36418 12155 36476 12161
rect 36418 12152 36430 12155
rect 35860 12124 36430 12152
rect 35860 12112 35866 12124
rect 36418 12121 36430 12124
rect 36464 12121 36476 12155
rect 36418 12115 36476 12121
rect 18414 12084 18420 12096
rect 16408 12056 18420 12084
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18598 12084 18604 12096
rect 18559 12056 18604 12084
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 25314 12044 25320 12096
rect 25372 12084 25378 12096
rect 26602 12084 26608 12096
rect 25372 12056 26608 12084
rect 25372 12044 25378 12056
rect 26602 12044 26608 12056
rect 26660 12084 26666 12096
rect 26789 12087 26847 12093
rect 26789 12084 26801 12087
rect 26660 12056 26801 12084
rect 26660 12044 26666 12056
rect 26789 12053 26801 12056
rect 26835 12053 26847 12087
rect 30926 12084 30932 12096
rect 30887 12056 30932 12084
rect 26789 12047 26847 12053
rect 30926 12044 30932 12056
rect 30984 12044 30990 12096
rect 34146 12084 34152 12096
rect 34107 12056 34152 12084
rect 34146 12044 34152 12056
rect 34204 12044 34210 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 11388 11852 13277 11880
rect 11388 11840 11394 11852
rect 13265 11849 13277 11852
rect 13311 11880 13323 11883
rect 13446 11880 13452 11892
rect 13311 11852 13452 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 19242 11880 19248 11892
rect 14047 11852 19248 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 2590 11772 2596 11824
rect 2648 11812 2654 11824
rect 2648 11784 7604 11812
rect 2648 11772 2654 11784
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 7466 11744 7472 11756
rect 1719 11716 7472 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7576 11676 7604 11784
rect 8938 11772 8944 11824
rect 8996 11812 9002 11824
rect 11606 11812 11612 11824
rect 8996 11784 11612 11812
rect 8996 11772 9002 11784
rect 11606 11772 11612 11784
rect 11664 11772 11670 11824
rect 13357 11815 13415 11821
rect 13357 11781 13369 11815
rect 13403 11812 13415 11815
rect 14016 11812 14044 11843
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 21818 11880 21824 11892
rect 21779 11852 21824 11880
rect 21818 11840 21824 11852
rect 21876 11840 21882 11892
rect 24394 11880 24400 11892
rect 24355 11852 24400 11880
rect 24394 11840 24400 11852
rect 24452 11840 24458 11892
rect 26142 11880 26148 11892
rect 26103 11852 26148 11880
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 26878 11840 26884 11892
rect 26936 11880 26942 11892
rect 28534 11880 28540 11892
rect 26936 11852 28540 11880
rect 26936 11840 26942 11852
rect 28534 11840 28540 11852
rect 28592 11840 28598 11892
rect 29086 11880 29092 11892
rect 29047 11852 29092 11880
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 31726 11852 35572 11880
rect 13403 11784 14044 11812
rect 13403 11781 13415 11784
rect 13357 11775 13415 11781
rect 16390 11772 16396 11824
rect 16448 11812 16454 11824
rect 31726 11812 31754 11852
rect 16448 11784 31754 11812
rect 16448 11772 16454 11784
rect 34146 11772 34152 11824
rect 34204 11812 34210 11824
rect 34762 11815 34820 11821
rect 34762 11812 34774 11815
rect 34204 11784 34774 11812
rect 34204 11772 34210 11784
rect 34762 11781 34774 11784
rect 34808 11781 34820 11815
rect 34762 11775 34820 11781
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11744 9367 11747
rect 9858 11744 9864 11756
rect 9355 11716 9864 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 12618 11744 12624 11756
rect 12483 11716 12624 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 22002 11744 22008 11756
rect 20588 11716 22008 11744
rect 20588 11704 20594 11716
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22278 11744 22284 11756
rect 22239 11716 22284 11744
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 22830 11744 22836 11756
rect 22520 11716 22836 11744
rect 22520 11704 22526 11716
rect 22830 11704 22836 11716
rect 22888 11704 22894 11756
rect 24578 11744 24584 11756
rect 24539 11716 24584 11744
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11713 24915 11747
rect 25038 11744 25044 11756
rect 24999 11716 25044 11744
rect 24857 11707 24915 11713
rect 17402 11676 17408 11688
rect 7576 11648 17408 11676
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 20441 11679 20499 11685
rect 20441 11676 20453 11679
rect 19392 11648 20453 11676
rect 19392 11636 19398 11648
rect 20441 11645 20453 11648
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 22296 11676 22324 11704
rect 24872 11676 24900 11707
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25314 11704 25320 11756
rect 25372 11744 25378 11756
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 25372 11716 25513 11744
rect 25372 11704 25378 11716
rect 25501 11713 25513 11716
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11713 25743 11747
rect 25958 11744 25964 11756
rect 25919 11716 25964 11744
rect 25685 11707 25743 11713
rect 25130 11676 25136 11688
rect 20763 11648 25136 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 25130 11636 25136 11648
rect 25188 11676 25194 11688
rect 25700 11676 25728 11707
rect 25958 11704 25964 11716
rect 26016 11704 26022 11756
rect 29270 11744 29276 11756
rect 29231 11716 29276 11744
rect 29270 11704 29276 11716
rect 29328 11704 29334 11756
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11713 29607 11747
rect 29549 11707 29607 11713
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11744 29791 11747
rect 30745 11747 30803 11753
rect 30745 11744 30757 11747
rect 29779 11716 30757 11744
rect 29779 11713 29791 11716
rect 29733 11707 29791 11713
rect 30745 11713 30757 11716
rect 30791 11744 30803 11747
rect 30926 11744 30932 11756
rect 30791 11716 30932 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 25188 11648 25728 11676
rect 25188 11636 25194 11648
rect 28534 11636 28540 11688
rect 28592 11676 28598 11688
rect 29564 11676 29592 11707
rect 28592 11648 29592 11676
rect 28592 11636 28598 11648
rect 1486 11608 1492 11620
rect 1447 11580 1492 11608
rect 1486 11568 1492 11580
rect 1544 11568 1550 11620
rect 2593 11611 2651 11617
rect 2593 11577 2605 11611
rect 2639 11608 2651 11611
rect 2866 11608 2872 11620
rect 2639 11580 2872 11608
rect 2639 11577 2651 11580
rect 2593 11571 2651 11577
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 9858 11608 9864 11620
rect 9771 11580 9864 11608
rect 9858 11568 9864 11580
rect 9916 11608 9922 11620
rect 10134 11608 10140 11620
rect 9916 11580 10140 11608
rect 9916 11568 9922 11580
rect 10134 11568 10140 11580
rect 10192 11608 10198 11620
rect 18138 11608 18144 11620
rect 10192 11580 18144 11608
rect 10192 11568 10198 11580
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 24762 11568 24768 11620
rect 24820 11608 24826 11620
rect 25038 11608 25044 11620
rect 24820 11580 25044 11608
rect 24820 11568 24826 11580
rect 25038 11568 25044 11580
rect 25096 11568 25102 11620
rect 25314 11568 25320 11620
rect 25372 11608 25378 11620
rect 25372 11580 27660 11608
rect 25372 11568 25378 11580
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 2832 11512 3065 11540
rect 2832 11500 2838 11512
rect 3053 11509 3065 11512
rect 3099 11509 3111 11543
rect 3053 11503 3111 11509
rect 9125 11543 9183 11549
rect 9125 11509 9137 11543
rect 9171 11540 9183 11543
rect 9214 11540 9220 11552
rect 9171 11512 9220 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 12250 11540 12256 11552
rect 12211 11512 12256 11540
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 27632 11540 27660 11580
rect 28902 11568 28908 11620
rect 28960 11608 28966 11620
rect 29748 11608 29776 11707
rect 30926 11704 30932 11716
rect 30984 11704 30990 11756
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 31386 11744 31392 11756
rect 31076 11716 31392 11744
rect 31076 11704 31082 11716
rect 31386 11704 31392 11716
rect 31444 11744 31450 11756
rect 32585 11747 32643 11753
rect 32585 11744 32597 11747
rect 31444 11716 32597 11744
rect 31444 11704 31450 11716
rect 32585 11713 32597 11716
rect 32631 11713 32643 11747
rect 32585 11707 32643 11713
rect 32769 11747 32827 11753
rect 32769 11713 32781 11747
rect 32815 11744 32827 11747
rect 34057 11747 34115 11753
rect 34057 11744 34069 11747
rect 32815 11716 34069 11744
rect 32815 11713 32827 11716
rect 32769 11707 32827 11713
rect 34057 11713 34069 11716
rect 34103 11744 34115 11747
rect 34422 11744 34428 11756
rect 34103 11716 34428 11744
rect 34103 11713 34115 11716
rect 34057 11707 34115 11713
rect 34422 11704 34428 11716
rect 34480 11744 34486 11756
rect 34517 11747 34575 11753
rect 34517 11744 34529 11747
rect 34480 11716 34529 11744
rect 34480 11704 34486 11716
rect 34517 11713 34529 11716
rect 34563 11713 34575 11747
rect 34517 11707 34575 11713
rect 28960 11580 29776 11608
rect 30944 11608 30972 11704
rect 32490 11608 32496 11620
rect 30944 11580 32496 11608
rect 28960 11568 28966 11580
rect 32490 11568 32496 11580
rect 32548 11568 32554 11620
rect 30193 11543 30251 11549
rect 30193 11540 30205 11543
rect 27632 11512 30205 11540
rect 30193 11509 30205 11512
rect 30239 11540 30251 11543
rect 30466 11540 30472 11552
rect 30239 11512 30472 11540
rect 30239 11509 30251 11512
rect 30193 11503 30251 11509
rect 30466 11500 30472 11512
rect 30524 11500 30530 11552
rect 35544 11540 35572 11852
rect 36998 11840 37004 11892
rect 37056 11880 37062 11892
rect 37056 11852 37780 11880
rect 37056 11840 37062 11852
rect 37090 11772 37096 11824
rect 37148 11812 37154 11824
rect 37553 11815 37611 11821
rect 37553 11812 37565 11815
rect 37148 11784 37565 11812
rect 37148 11772 37154 11784
rect 37553 11781 37565 11784
rect 37599 11781 37611 11815
rect 37553 11775 37611 11781
rect 37274 11744 37280 11756
rect 37235 11716 37280 11744
rect 37274 11704 37280 11716
rect 37332 11704 37338 11756
rect 37366 11704 37372 11756
rect 37424 11744 37430 11756
rect 37752 11753 37780 11852
rect 37645 11747 37703 11753
rect 37424 11716 37469 11744
rect 37424 11704 37430 11716
rect 37645 11713 37657 11747
rect 37691 11713 37703 11747
rect 37645 11707 37703 11713
rect 37742 11747 37800 11753
rect 37742 11713 37754 11747
rect 37788 11713 37800 11747
rect 37742 11707 37800 11713
rect 37182 11676 37188 11688
rect 35912 11648 37188 11676
rect 35912 11617 35940 11648
rect 37182 11636 37188 11648
rect 37240 11676 37246 11688
rect 37660 11676 37688 11707
rect 37240 11648 37688 11676
rect 37240 11636 37246 11648
rect 35897 11611 35955 11617
rect 35897 11577 35909 11611
rect 35943 11577 35955 11611
rect 35897 11571 35955 11577
rect 37921 11543 37979 11549
rect 37921 11540 37933 11543
rect 35544 11512 37933 11540
rect 37921 11509 37933 11512
rect 37967 11509 37979 11543
rect 37921 11503 37979 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 7374 11336 7380 11348
rect 2179 11308 7380 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 10137 11339 10195 11345
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 10962 11336 10968 11348
rect 10183 11308 10968 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 1854 11132 1860 11144
rect 1767 11104 1860 11132
rect 1854 11092 1860 11104
rect 1912 11132 1918 11144
rect 2774 11132 2780 11144
rect 1912 11104 2780 11132
rect 1912 11092 1918 11104
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 9493 11135 9551 11141
rect 2924 11104 2969 11132
rect 2924 11092 2930 11104
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 10152 11132 10180 11299
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 12710 11336 12716 11348
rect 11072 11308 12572 11336
rect 12671 11308 12716 11336
rect 9539 11104 10180 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 11072 11064 11100 11308
rect 12437 11271 12495 11277
rect 12437 11237 12449 11271
rect 12483 11237 12495 11271
rect 12544 11268 12572 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 15378 11336 15384 11348
rect 12820 11308 15384 11336
rect 12820 11268 12848 11308
rect 15378 11296 15384 11308
rect 15436 11336 15442 11348
rect 15436 11308 15792 11336
rect 15436 11296 15442 11308
rect 12544 11240 12848 11268
rect 12437 11231 12495 11237
rect 12452 11200 12480 11231
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 14829 11271 14887 11277
rect 14829 11268 14841 11271
rect 13228 11240 14841 11268
rect 13228 11228 13234 11240
rect 14829 11237 14841 11240
rect 14875 11268 14887 11271
rect 15654 11268 15660 11280
rect 14875 11240 15660 11268
rect 14875 11237 14887 11240
rect 14829 11231 14887 11237
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 15764 11268 15792 11308
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15896 11308 16313 11336
rect 15896 11296 15902 11308
rect 16301 11305 16313 11308
rect 16347 11336 16359 11339
rect 16390 11336 16396 11348
rect 16347 11308 16396 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 16758 11336 16764 11348
rect 16719 11308 16764 11336
rect 16758 11296 16764 11308
rect 16816 11336 16822 11348
rect 17126 11336 17132 11348
rect 16816 11308 17132 11336
rect 16816 11296 16822 11308
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 25406 11296 25412 11348
rect 25464 11336 25470 11348
rect 26053 11339 26111 11345
rect 26053 11336 26065 11339
rect 25464 11308 26065 11336
rect 25464 11296 25470 11308
rect 26053 11305 26065 11308
rect 26099 11305 26111 11339
rect 26053 11299 26111 11305
rect 29270 11296 29276 11348
rect 29328 11336 29334 11348
rect 31754 11336 31760 11348
rect 29328 11308 31760 11336
rect 29328 11296 29334 11308
rect 31754 11296 31760 11308
rect 31812 11336 31818 11348
rect 33042 11336 33048 11348
rect 31812 11308 33048 11336
rect 31812 11296 31818 11308
rect 33042 11296 33048 11308
rect 33100 11296 33106 11348
rect 36633 11339 36691 11345
rect 36633 11305 36645 11339
rect 36679 11336 36691 11339
rect 37366 11336 37372 11348
rect 36679 11308 37372 11336
rect 36679 11305 36691 11308
rect 36633 11299 36691 11305
rect 37366 11296 37372 11308
rect 37424 11296 37430 11348
rect 38010 11336 38016 11348
rect 37971 11308 38016 11336
rect 38010 11296 38016 11308
rect 38068 11296 38074 11348
rect 25590 11268 25596 11280
rect 15764 11240 25452 11268
rect 25551 11240 25596 11268
rect 14737 11203 14795 11209
rect 12452 11172 14688 11200
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 11664 11104 12633 11132
rect 11664 11092 11670 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 14182 11132 14188 11144
rect 12943 11104 14188 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 9732 11036 11100 11064
rect 9732 11024 9738 11036
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 12728 11064 12756 11095
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 14660 11141 14688 11172
rect 14737 11169 14749 11203
rect 14783 11200 14795 11203
rect 15194 11200 15200 11212
rect 14783 11172 15200 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 17402 11160 17408 11212
rect 17460 11200 17466 11212
rect 25314 11200 25320 11212
rect 17460 11172 25320 11200
rect 17460 11160 17466 11172
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 25424 11200 25452 11240
rect 25590 11228 25596 11240
rect 25648 11228 25654 11280
rect 32490 11228 32496 11280
rect 32548 11268 32554 11280
rect 36078 11268 36084 11280
rect 32548 11240 36084 11268
rect 32548 11228 32554 11240
rect 36078 11228 36084 11240
rect 36136 11228 36142 11280
rect 37182 11228 37188 11280
rect 37240 11268 37246 11280
rect 37277 11271 37335 11277
rect 37277 11268 37289 11271
rect 37240 11240 37289 11268
rect 37240 11228 37246 11240
rect 37277 11237 37289 11240
rect 37323 11237 37335 11271
rect 37277 11231 37335 11237
rect 29549 11203 29607 11209
rect 29549 11200 29561 11203
rect 25424 11172 29561 11200
rect 29549 11169 29561 11172
rect 29595 11169 29607 11203
rect 29549 11163 29607 11169
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11132 14979 11135
rect 15930 11132 15936 11144
rect 14967 11104 15936 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 24670 11092 24676 11144
rect 24728 11132 24734 11144
rect 24949 11135 25007 11141
rect 24949 11132 24961 11135
rect 24728 11104 24961 11132
rect 24728 11092 24734 11104
rect 24949 11101 24961 11104
rect 24995 11101 25007 11135
rect 25130 11132 25136 11144
rect 25091 11104 25136 11132
rect 24949 11095 25007 11101
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25409 11135 25467 11141
rect 25409 11101 25421 11135
rect 25455 11132 25467 11135
rect 25958 11132 25964 11144
rect 25455 11104 25964 11132
rect 25455 11101 25467 11104
rect 25409 11095 25467 11101
rect 12492 11036 12756 11064
rect 16684 11036 16896 11064
rect 12492 11024 12498 11036
rect 2682 10996 2688 11008
rect 2643 10968 2688 10996
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 9398 10996 9404 11008
rect 9359 10968 9404 10996
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 15102 10996 15108 11008
rect 15063 10968 15108 10996
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 16684 10996 16712 11036
rect 15344 10968 16712 10996
rect 16868 10996 16896 11036
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19426 11064 19432 11076
rect 19116 11036 19432 11064
rect 19116 11024 19122 11036
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 24578 11024 24584 11076
rect 24636 11064 24642 11076
rect 25424 11064 25452 11095
rect 25958 11092 25964 11104
rect 26016 11092 26022 11144
rect 29564 11132 29592 11163
rect 30374 11160 30380 11212
rect 30432 11200 30438 11212
rect 30653 11203 30711 11209
rect 30653 11200 30665 11203
rect 30432 11172 30665 11200
rect 30432 11160 30438 11172
rect 30653 11169 30665 11172
rect 30699 11169 30711 11203
rect 30653 11163 30711 11169
rect 30469 11135 30527 11141
rect 30469 11132 30481 11135
rect 29564 11104 30481 11132
rect 30469 11101 30481 11104
rect 30515 11132 30527 11135
rect 33502 11132 33508 11144
rect 30515 11104 33508 11132
rect 30515 11101 30527 11104
rect 30469 11095 30527 11101
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 35989 11135 36047 11141
rect 35989 11101 36001 11135
rect 36035 11132 36047 11135
rect 36446 11132 36452 11144
rect 36035 11104 36452 11132
rect 36035 11101 36047 11104
rect 35989 11095 36047 11101
rect 36446 11092 36452 11104
rect 36504 11092 36510 11144
rect 37093 11135 37151 11141
rect 37093 11101 37105 11135
rect 37139 11132 37151 11135
rect 37642 11132 37648 11144
rect 37139 11104 37648 11132
rect 37139 11101 37151 11104
rect 37093 11095 37151 11101
rect 37642 11092 37648 11104
rect 37700 11092 37706 11144
rect 37829 11135 37887 11141
rect 37829 11101 37841 11135
rect 37875 11101 37887 11135
rect 37829 11095 37887 11101
rect 30558 11064 30564 11076
rect 24636 11036 25452 11064
rect 30519 11036 30564 11064
rect 24636 11024 24642 11036
rect 30558 11024 30564 11036
rect 30616 11064 30622 11076
rect 32674 11064 32680 11076
rect 30616 11036 32680 11064
rect 30616 11024 30622 11036
rect 32674 11024 32680 11036
rect 32732 11064 32738 11076
rect 37844 11064 37872 11095
rect 32732 11036 37872 11064
rect 32732 11024 32738 11036
rect 19150 10996 19156 11008
rect 16868 10968 19156 10996
rect 15344 10956 15350 10968
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 30101 10999 30159 11005
rect 30101 10965 30113 10999
rect 30147 10996 30159 10999
rect 30282 10996 30288 11008
rect 30147 10968 30288 10996
rect 30147 10965 30159 10968
rect 30101 10959 30159 10965
rect 30282 10956 30288 10968
rect 30340 10956 30346 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 8864 10764 9505 10792
rect 8864 10733 8892 10764
rect 9493 10761 9505 10764
rect 9539 10792 9551 10795
rect 9582 10792 9588 10804
rect 9539 10764 9588 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 16942 10792 16948 10804
rect 15764 10764 16948 10792
rect 8849 10727 8907 10733
rect 8849 10693 8861 10727
rect 8895 10693 8907 10727
rect 8849 10687 8907 10693
rect 11514 10684 11520 10736
rect 11572 10724 11578 10736
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 11572 10696 11989 10724
rect 11572 10684 11578 10696
rect 11977 10693 11989 10696
rect 12023 10724 12035 10727
rect 12250 10724 12256 10736
rect 12023 10696 12256 10724
rect 12023 10693 12035 10696
rect 11977 10687 12035 10693
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 12526 10684 12532 10736
rect 12584 10724 12590 10736
rect 13541 10727 13599 10733
rect 12584 10696 12940 10724
rect 12584 10684 12590 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2590 10656 2596 10668
rect 1719 10628 2596 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 8260 10628 11713 10656
rect 8260 10616 8266 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 11701 10619 11759 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12912 10665 12940 10696
rect 13541 10693 13553 10727
rect 13587 10724 13599 10727
rect 15286 10724 15292 10736
rect 13587 10696 15292 10724
rect 13587 10693 13599 10696
rect 13541 10687 13599 10693
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 15764 10733 15792 10764
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 21174 10752 21180 10804
rect 21232 10792 21238 10804
rect 22370 10792 22376 10804
rect 21232 10764 22376 10792
rect 21232 10752 21238 10764
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 25498 10752 25504 10804
rect 25556 10792 25562 10804
rect 25685 10795 25743 10801
rect 25685 10792 25697 10795
rect 25556 10764 25697 10792
rect 25556 10752 25562 10764
rect 25685 10761 25697 10764
rect 25731 10761 25743 10795
rect 25685 10755 25743 10761
rect 37274 10752 37280 10804
rect 37332 10792 37338 10804
rect 37369 10795 37427 10801
rect 37369 10792 37381 10795
rect 37332 10764 37381 10792
rect 37332 10752 37338 10764
rect 37369 10761 37381 10764
rect 37415 10792 37427 10795
rect 38286 10792 38292 10804
rect 37415 10764 38292 10792
rect 37415 10761 37427 10764
rect 37369 10755 37427 10761
rect 38286 10752 38292 10764
rect 38344 10752 38350 10804
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10693 15807 10727
rect 15749 10687 15807 10693
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 27614 10724 27620 10736
rect 15896 10696 15941 10724
rect 16776 10696 27620 10724
rect 15896 10684 15902 10696
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 12986 10656 12992 10668
rect 12943 10628 12992 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13136 10628 13229 10656
rect 13136 10616 13142 10628
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15160 10628 15485 10656
rect 15160 10616 15166 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15562 10616 15568 10668
rect 15620 10665 15626 10668
rect 15620 10659 15669 10665
rect 15620 10625 15623 10659
rect 15657 10625 15669 10659
rect 15620 10619 15669 10625
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16776 10656 16804 10696
rect 27614 10684 27620 10696
rect 27672 10684 27678 10736
rect 29825 10727 29883 10733
rect 29825 10693 29837 10727
rect 29871 10724 29883 10727
rect 31018 10724 31024 10736
rect 29871 10696 31024 10724
rect 29871 10693 29883 10696
rect 29825 10687 29883 10693
rect 31018 10684 31024 10696
rect 31076 10684 31082 10736
rect 15979 10628 16804 10656
rect 16853 10659 16911 10665
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 17494 10656 17500 10668
rect 16899 10628 17500 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 15620 10616 15626 10619
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 18012 10628 19073 10656
rect 18012 10616 18018 10628
rect 19061 10625 19073 10628
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19334 10656 19340 10668
rect 19291 10628 19340 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19978 10656 19984 10668
rect 19484 10628 19984 10656
rect 19484 10616 19490 10628
rect 19978 10616 19984 10628
rect 20036 10656 20042 10668
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 20036 10628 20085 10656
rect 20036 10616 20042 10628
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10656 25283 10659
rect 25406 10656 25412 10668
rect 25271 10628 25412 10656
rect 25271 10625 25283 10628
rect 25225 10619 25283 10625
rect 25406 10616 25412 10628
rect 25464 10656 25470 10668
rect 25774 10656 25780 10668
rect 25464 10628 25780 10656
rect 25464 10616 25470 10628
rect 25774 10616 25780 10628
rect 25832 10616 25838 10668
rect 32306 10616 32312 10668
rect 32364 10656 32370 10668
rect 37829 10659 37887 10665
rect 37829 10656 37841 10659
rect 32364 10628 37841 10656
rect 32364 10616 32370 10628
rect 37829 10625 37841 10628
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 12434 10588 12440 10600
rect 11931 10560 12440 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13096 10588 13124 10616
rect 12676 10560 13124 10588
rect 12676 10548 12682 10560
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 16816 10560 17049 10588
rect 16816 10548 16822 10560
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 17184 10560 17229 10588
rect 17184 10548 17190 10560
rect 18138 10548 18144 10600
rect 18196 10588 18202 10600
rect 22554 10588 22560 10600
rect 18196 10560 22560 10588
rect 18196 10548 18202 10560
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 29730 10588 29736 10600
rect 25884 10560 29736 10588
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 17957 10523 18015 10529
rect 17957 10520 17969 10523
rect 6972 10492 12848 10520
rect 6972 10480 6978 10492
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 2096 10424 2145 10452
rect 2096 10412 2102 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10452 2835 10455
rect 2958 10452 2964 10464
rect 2823 10424 2964 10452
rect 2823 10421 2835 10424
rect 2777 10415 2835 10421
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 8444 10424 8769 10452
rect 8444 10412 8450 10424
rect 8757 10421 8769 10424
rect 8803 10421 8815 10455
rect 8757 10415 8815 10421
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11020 10424 11529 10452
rect 11020 10412 11026 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 11977 10455 12035 10461
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12710 10452 12716 10464
rect 12023 10424 12716 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12820 10452 12848 10492
rect 15948 10492 17969 10520
rect 15948 10452 15976 10492
rect 17957 10489 17969 10492
rect 18003 10520 18015 10523
rect 18506 10520 18512 10532
rect 18003 10492 18512 10520
rect 18003 10489 18015 10492
rect 17957 10483 18015 10489
rect 18506 10480 18512 10492
rect 18564 10520 18570 10532
rect 25884 10520 25912 10560
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 18564 10492 25912 10520
rect 18564 10480 18570 10492
rect 29546 10480 29552 10532
rect 29604 10520 29610 10532
rect 29641 10523 29699 10529
rect 29641 10520 29653 10523
rect 29604 10492 29653 10520
rect 29604 10480 29610 10492
rect 29641 10489 29653 10492
rect 29687 10489 29699 10523
rect 29641 10483 29699 10489
rect 16114 10452 16120 10464
rect 12820 10424 15976 10452
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16669 10455 16727 10461
rect 16669 10421 16681 10455
rect 16715 10452 16727 10455
rect 16850 10452 16856 10464
rect 16715 10424 16856 10452
rect 16715 10421 16727 10424
rect 16669 10415 16727 10421
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 19889 10455 19947 10461
rect 19889 10452 19901 10455
rect 19024 10424 19901 10452
rect 19024 10412 19030 10424
rect 19889 10421 19901 10424
rect 19935 10452 19947 10455
rect 22094 10452 22100 10464
rect 19935 10424 22100 10452
rect 19935 10421 19947 10424
rect 19889 10415 19947 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22370 10412 22376 10464
rect 22428 10452 22434 10464
rect 22649 10455 22707 10461
rect 22649 10452 22661 10455
rect 22428 10424 22661 10452
rect 22428 10412 22434 10424
rect 22649 10421 22661 10424
rect 22695 10452 22707 10455
rect 28166 10452 28172 10464
rect 22695 10424 28172 10452
rect 22695 10421 22707 10424
rect 22649 10415 22707 10421
rect 28166 10412 28172 10424
rect 28224 10412 28230 10464
rect 38010 10452 38016 10464
rect 37971 10424 38016 10452
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2314 10248 2320 10260
rect 2179 10220 2320 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 10778 10248 10784 10260
rect 10735 10220 10784 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 10778 10208 10784 10220
rect 10836 10248 10842 10260
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 10836 10220 11621 10248
rect 10836 10208 10842 10220
rect 11609 10217 11621 10220
rect 11655 10248 11667 10251
rect 12710 10248 12716 10260
rect 11655 10220 12716 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 13538 10248 13544 10260
rect 12952 10220 13544 10248
rect 12952 10208 12958 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13964 10220 14105 10248
rect 13964 10208 13970 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17589 10251 17647 10257
rect 17589 10248 17601 10251
rect 17552 10220 17601 10248
rect 17552 10208 17558 10220
rect 17589 10217 17601 10220
rect 17635 10217 17647 10251
rect 22554 10248 22560 10260
rect 22515 10220 22560 10248
rect 17589 10211 17647 10217
rect 22554 10208 22560 10220
rect 22612 10248 22618 10260
rect 23750 10248 23756 10260
rect 22612 10220 23756 10248
rect 22612 10208 22618 10220
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 27614 10248 27620 10260
rect 27575 10220 27620 10248
rect 27614 10208 27620 10220
rect 27672 10208 27678 10260
rect 32585 10251 32643 10257
rect 32585 10217 32597 10251
rect 32631 10248 32643 10251
rect 32674 10248 32680 10260
rect 32631 10220 32680 10248
rect 32631 10217 32643 10220
rect 32585 10211 32643 10217
rect 32674 10208 32680 10220
rect 32732 10208 32738 10260
rect 35802 10248 35808 10260
rect 35763 10220 35808 10248
rect 35802 10208 35808 10220
rect 35860 10208 35866 10260
rect 36262 10248 36268 10260
rect 36223 10220 36268 10248
rect 36262 10208 36268 10220
rect 36320 10208 36326 10260
rect 2590 10140 2596 10192
rect 2648 10180 2654 10192
rect 16114 10180 16120 10192
rect 2648 10152 16120 10180
rect 2648 10140 2654 10152
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 16758 10140 16764 10192
rect 16816 10180 16822 10192
rect 18417 10183 18475 10189
rect 18417 10180 18429 10183
rect 16816 10152 18429 10180
rect 16816 10140 16822 10152
rect 18417 10149 18429 10152
rect 18463 10180 18475 10183
rect 19150 10180 19156 10192
rect 18463 10152 19156 10180
rect 18463 10149 18475 10152
rect 18417 10143 18475 10149
rect 19150 10140 19156 10152
rect 19208 10180 19214 10192
rect 19245 10183 19303 10189
rect 19245 10180 19257 10183
rect 19208 10152 19257 10180
rect 19208 10140 19214 10152
rect 19245 10149 19257 10152
rect 19291 10149 19303 10183
rect 30282 10180 30288 10192
rect 30243 10152 30288 10180
rect 19245 10143 19303 10149
rect 30282 10140 30288 10152
rect 30340 10140 30346 10192
rect 8294 10112 8300 10124
rect 8036 10084 8300 10112
rect 1854 10044 1860 10056
rect 1767 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10044 1918 10056
rect 3234 10044 3240 10056
rect 1912 10016 3240 10044
rect 1912 10004 1918 10016
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 8036 10053 8064 10084
rect 8294 10072 8300 10084
rect 8352 10112 8358 10124
rect 9398 10112 9404 10124
rect 8352 10084 9404 10112
rect 8352 10072 8358 10084
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 10594 10112 10600 10124
rect 10507 10084 10600 10112
rect 10594 10072 10600 10084
rect 10652 10112 10658 10124
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 10652 10084 11529 10112
rect 10652 10072 10658 10084
rect 11517 10081 11529 10084
rect 11563 10112 11575 10115
rect 12434 10112 12440 10124
rect 11563 10084 12440 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 12434 10072 12440 10084
rect 12492 10112 12498 10124
rect 12492 10084 12756 10112
rect 12492 10072 12498 10084
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 8021 10007 8079 10013
rect 7760 9976 7788 10007
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 9824 10016 10701 10044
rect 9824 10004 9830 10016
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 11112 10016 11621 10044
rect 11112 10004 11118 10016
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 9214 9976 9220 9988
rect 7760 9948 9220 9976
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 10413 9979 10471 9985
rect 10413 9945 10425 9979
rect 10459 9976 10471 9979
rect 11333 9979 11391 9985
rect 11333 9976 11345 9979
rect 10459 9948 11345 9976
rect 10459 9945 10471 9948
rect 10413 9939 10471 9945
rect 11333 9945 11345 9948
rect 11379 9976 11391 9979
rect 11514 9976 11520 9988
rect 11379 9948 11520 9976
rect 11379 9945 11391 9948
rect 11333 9939 11391 9945
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2832 9880 2877 9908
rect 2832 9868 2838 9880
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7340 9880 7573 9908
rect 7340 9868 7346 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 7561 9871 7619 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 11793 9911 11851 9917
rect 11793 9908 11805 9911
rect 11756 9880 11805 9908
rect 11756 9868 11762 9880
rect 11793 9877 11805 9880
rect 11839 9877 11851 9911
rect 12728 9908 12756 10084
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 15841 10115 15899 10121
rect 15841 10112 15853 10115
rect 15252 10084 15853 10112
rect 15252 10072 15258 10084
rect 15841 10081 15853 10084
rect 15887 10081 15899 10115
rect 17954 10112 17960 10124
rect 15841 10075 15899 10081
rect 17144 10084 17960 10112
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 13538 10044 13544 10056
rect 13499 10016 13544 10044
rect 12897 10007 12955 10013
rect 12912 9976 12940 10007
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16482 10044 16488 10056
rect 16163 10016 16488 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17144 10053 17172 10084
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18506 10112 18512 10124
rect 18467 10084 18512 10112
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 19978 10112 19984 10124
rect 19891 10084 19984 10112
rect 19978 10072 19984 10084
rect 20036 10112 20042 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 20036 10084 21281 10112
rect 20036 10072 20042 10084
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 25498 10112 25504 10124
rect 25459 10084 25504 10112
rect 21269 10075 21327 10081
rect 25498 10072 25504 10084
rect 25556 10072 25562 10124
rect 30558 10112 30564 10124
rect 27816 10084 30564 10112
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10013 17463 10047
rect 18230 10044 18236 10056
rect 18191 10016 18236 10044
rect 17405 10007 17463 10013
rect 13906 9976 13912 9988
rect 12912 9948 13912 9976
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 16500 9976 16528 10004
rect 17310 9976 17316 9988
rect 16500 9948 17316 9976
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 17420 9976 17448 10007
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 20070 10004 20076 10056
rect 20128 10044 20134 10056
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 20128 10016 20269 10044
rect 20128 10004 20134 10016
rect 20257 10013 20269 10016
rect 20303 10044 20315 10047
rect 20530 10044 20536 10056
rect 20303 10016 20536 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 23750 10004 23756 10056
rect 23808 10044 23814 10056
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 23808 10016 24409 10044
rect 23808 10004 23814 10016
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 25593 10047 25651 10053
rect 25593 10013 25605 10047
rect 25639 10013 25651 10047
rect 25774 10044 25780 10056
rect 25735 10016 25780 10044
rect 25593 10007 25651 10013
rect 20088 9976 20116 10004
rect 17420 9948 20116 9976
rect 25498 9936 25504 9988
rect 25556 9976 25562 9988
rect 25608 9976 25636 10007
rect 25774 10004 25780 10016
rect 25832 10004 25838 10056
rect 27816 10053 27844 10084
rect 30558 10072 30564 10084
rect 30616 10072 30622 10124
rect 36630 10072 36636 10124
rect 36688 10112 36694 10124
rect 37001 10115 37059 10121
rect 37001 10112 37013 10115
rect 36688 10084 37013 10112
rect 36688 10072 36694 10084
rect 37001 10081 37013 10084
rect 37047 10081 37059 10115
rect 37001 10075 37059 10081
rect 27801 10047 27859 10053
rect 27801 10013 27813 10047
rect 27847 10013 27859 10047
rect 27801 10007 27859 10013
rect 29546 10004 29552 10056
rect 29604 10044 29610 10056
rect 31205 10047 31263 10053
rect 31205 10044 31217 10047
rect 29604 10016 31217 10044
rect 29604 10004 29610 10016
rect 31205 10013 31217 10016
rect 31251 10013 31263 10047
rect 31205 10007 31263 10013
rect 37277 10047 37335 10053
rect 37277 10013 37289 10047
rect 37323 10044 37335 10047
rect 37734 10044 37740 10056
rect 37323 10016 37740 10044
rect 37323 10013 37335 10016
rect 37277 10007 37335 10013
rect 37734 10004 37740 10016
rect 37792 10004 37798 10056
rect 26421 9979 26479 9985
rect 26421 9976 26433 9979
rect 25556 9948 26433 9976
rect 25556 9936 25562 9948
rect 26421 9945 26433 9948
rect 26467 9976 26479 9979
rect 26970 9976 26976 9988
rect 26467 9948 26976 9976
rect 26467 9945 26479 9948
rect 26421 9939 26479 9945
rect 26970 9936 26976 9948
rect 27028 9936 27034 9988
rect 27706 9936 27712 9988
rect 27764 9976 27770 9988
rect 27985 9979 28043 9985
rect 27985 9976 27997 9979
rect 27764 9948 27997 9976
rect 27764 9936 27770 9948
rect 27985 9945 27997 9948
rect 28031 9945 28043 9979
rect 30006 9976 30012 9988
rect 29967 9948 30012 9976
rect 27985 9939 28043 9945
rect 30006 9936 30012 9948
rect 30064 9936 30070 9988
rect 30834 9936 30840 9988
rect 30892 9976 30898 9988
rect 31450 9979 31508 9985
rect 31450 9976 31462 9979
rect 30892 9948 31462 9976
rect 30892 9936 30898 9948
rect 31450 9945 31462 9948
rect 31496 9945 31508 9979
rect 31450 9939 31508 9945
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12728 9880 13369 9908
rect 11793 9871 11851 9877
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13924 9908 13952 9936
rect 17862 9908 17868 9920
rect 13924 9880 17868 9908
rect 13357 9871 13415 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18046 9908 18052 9920
rect 18007 9880 18052 9908
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22152 9880 22197 9908
rect 22152 9868 22158 9880
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 22922 9908 22928 9920
rect 22428 9880 22928 9908
rect 22428 9868 22434 9880
rect 22922 9868 22928 9880
rect 22980 9908 22986 9920
rect 23109 9911 23167 9917
rect 23109 9908 23121 9911
rect 22980 9880 23121 9908
rect 22980 9868 22986 9880
rect 23109 9877 23121 9880
rect 23155 9877 23167 9911
rect 24578 9908 24584 9920
rect 24539 9880 24584 9908
rect 23109 9871 23167 9877
rect 24578 9868 24584 9880
rect 24636 9868 24642 9920
rect 25961 9911 26019 9917
rect 25961 9877 25973 9911
rect 26007 9908 26019 9911
rect 26142 9908 26148 9920
rect 26007 9880 26148 9908
rect 26007 9877 26019 9880
rect 25961 9871 26019 9877
rect 26142 9868 26148 9880
rect 26200 9868 26206 9920
rect 30469 9911 30527 9917
rect 30469 9877 30481 9911
rect 30515 9908 30527 9911
rect 30650 9908 30656 9920
rect 30515 9880 30656 9908
rect 30515 9877 30527 9880
rect 30469 9871 30527 9877
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 8018 9704 8024 9716
rect 3936 9676 8024 9704
rect 3936 9664 3942 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 11514 9704 11520 9716
rect 10520 9676 11520 9704
rect 2774 9636 2780 9648
rect 1412 9608 2780 9636
rect 1412 9580 1440 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 8294 9636 8300 9648
rect 5092 9608 8300 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3033 9571 3091 9577
rect 3033 9568 3045 9571
rect 2924 9540 3045 9568
rect 2924 9528 2930 9540
rect 3033 9537 3045 9540
rect 3079 9537 3091 9571
rect 3033 9531 3091 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 4816 9500 4844 9531
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5092 9577 5120 9608
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 10520 9645 10548 9676
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 17402 9704 17408 9716
rect 11848 9676 17408 9704
rect 11848 9664 11854 9676
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 18874 9704 18880 9716
rect 17920 9676 18880 9704
rect 17920 9664 17926 9676
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 22370 9704 22376 9716
rect 22331 9676 22376 9704
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 23750 9664 23756 9716
rect 23808 9704 23814 9716
rect 23937 9707 23995 9713
rect 23937 9704 23949 9707
rect 23808 9676 23949 9704
rect 23808 9664 23814 9676
rect 23937 9673 23949 9676
rect 23983 9673 23995 9707
rect 26970 9704 26976 9716
rect 26931 9676 26976 9704
rect 23937 9667 23995 9673
rect 26970 9664 26976 9676
rect 27028 9664 27034 9716
rect 30834 9704 30840 9716
rect 30795 9676 30840 9704
rect 30834 9664 30840 9676
rect 30892 9664 30898 9716
rect 10505 9639 10563 9645
rect 10505 9605 10517 9639
rect 10551 9605 10563 9639
rect 10505 9599 10563 9605
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 10928 9608 13400 9636
rect 10928 9596 10934 9608
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 5040 9540 5089 9568
rect 5040 9528 5046 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5258 9568 5264 9580
rect 5219 9540 5264 9568
rect 5077 9531 5135 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7064 9540 7205 9568
rect 7064 9528 7070 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7460 9571 7518 9577
rect 7460 9537 7472 9571
rect 7506 9568 7518 9571
rect 8018 9568 8024 9580
rect 7506 9540 8024 9568
rect 7506 9537 7518 9540
rect 7460 9531 7518 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 9214 9568 9220 9580
rect 9175 9540 9220 9568
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 9456 9540 9505 9568
rect 9456 9528 9462 9540
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9766 9568 9772 9580
rect 9723 9540 9772 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 4816 9472 5488 9500
rect 2777 9463 2835 9469
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2498 9364 2504 9376
rect 2271 9336 2504 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2792 9364 2820 9463
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 5258 9432 5264 9444
rect 4203 9404 5264 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 5460 9376 5488 9472
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9432 8631 9435
rect 9692 9432 9720 9531
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 9916 9540 10793 9568
rect 9916 9528 9922 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12069 9571 12127 9577
rect 12381 9574 12439 9577
rect 12069 9568 12081 9571
rect 12032 9540 12081 9568
rect 12032 9528 12038 9540
rect 12069 9537 12081 9540
rect 12115 9537 12127 9571
rect 12268 9571 12439 9574
rect 12268 9568 12393 9571
rect 12069 9531 12127 9537
rect 12176 9546 12393 9568
rect 12176 9540 12296 9546
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 12176 9500 12204 9540
rect 12381 9537 12393 9546
rect 12427 9537 12439 9571
rect 12381 9531 12439 9537
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 10980 9472 12204 9500
rect 10980 9441 11008 9472
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 13096 9500 13124 9531
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 13372 9577 13400 9608
rect 13538 9596 13544 9648
rect 13596 9636 13602 9648
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 13596 9608 14105 9636
rect 13596 9596 13602 9608
rect 14093 9605 14105 9608
rect 14139 9605 14151 9639
rect 14093 9599 14151 9605
rect 17672 9639 17730 9645
rect 17672 9605 17684 9639
rect 17718 9636 17730 9639
rect 18046 9636 18052 9648
rect 17718 9608 18052 9636
rect 17718 9605 17730 9608
rect 17672 9599 17730 9605
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 19392 9608 20484 9636
rect 19392 9596 19398 9608
rect 13357 9571 13415 9577
rect 13228 9540 13273 9568
rect 13228 9528 13234 9540
rect 13357 9537 13369 9571
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 19300 9540 19441 9568
rect 19300 9528 19306 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19518 9528 19524 9580
rect 19576 9568 19582 9580
rect 20070 9568 20076 9580
rect 19576 9540 20076 9568
rect 19576 9528 19582 9540
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 20456 9577 20484 9608
rect 20622 9596 20628 9648
rect 20680 9636 20686 9648
rect 22281 9639 22339 9645
rect 20680 9608 22094 9636
rect 20680 9596 20686 9608
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9537 20499 9571
rect 20441 9531 20499 9537
rect 12308 9472 12353 9500
rect 13096 9472 13400 9500
rect 12308 9460 12314 9472
rect 13372 9444 13400 9472
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13688 9472 13921 9500
rect 13688 9460 13694 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 17184 9472 17417 9500
rect 17184 9460 17190 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 19150 9460 19156 9512
rect 19208 9500 19214 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19208 9472 19625 9500
rect 19208 9460 19214 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 8619 9404 9720 9432
rect 10965 9435 11023 9441
rect 8619 9401 8631 9404
rect 8573 9395 8631 9401
rect 10965 9401 10977 9435
rect 11011 9401 11023 9435
rect 12158 9432 12164 9444
rect 12119 9404 12164 9432
rect 10965 9395 11023 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 13265 9435 13323 9441
rect 13265 9432 13277 9435
rect 12452 9404 13277 9432
rect 3786 9364 3792 9376
rect 2792 9336 3792 9364
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4614 9364 4620 9376
rect 4575 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5813 9367 5871 9373
rect 5813 9364 5825 9367
rect 5500 9336 5825 9364
rect 5500 9324 5506 9336
rect 5813 9333 5825 9336
rect 5859 9364 5871 9367
rect 7374 9364 7380 9376
rect 5859 9336 7380 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 9033 9367 9091 9373
rect 9033 9364 9045 9367
rect 8352 9336 9045 9364
rect 8352 9324 8358 9336
rect 9033 9333 9045 9336
rect 9079 9333 9091 9367
rect 10778 9364 10784 9376
rect 10739 9336 10784 9364
rect 9033 9327 9091 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 12250 9364 12256 9376
rect 12124 9336 12256 9364
rect 12124 9324 12130 9336
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 12452 9364 12480 9404
rect 13265 9401 13277 9404
rect 13311 9401 13323 9435
rect 13265 9395 13323 9401
rect 12894 9364 12900 9376
rect 12308 9336 12480 9364
rect 12855 9336 12900 9364
rect 12308 9324 12314 9336
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13280 9364 13308 9395
rect 13354 9392 13360 9444
rect 13412 9392 13418 9444
rect 19720 9432 19748 9463
rect 20438 9432 20444 9444
rect 19720 9404 20444 9432
rect 20438 9392 20444 9404
rect 20496 9392 20502 9444
rect 22066 9432 22094 9608
rect 22281 9605 22293 9639
rect 22327 9636 22339 9639
rect 22554 9636 22560 9648
rect 22327 9608 22560 9636
rect 22327 9605 22339 9608
rect 22281 9599 22339 9605
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 23014 9596 23020 9648
rect 23072 9636 23078 9648
rect 23290 9636 23296 9648
rect 23072 9608 23296 9636
rect 23072 9596 23078 9608
rect 23290 9596 23296 9608
rect 23348 9596 23354 9648
rect 24673 9639 24731 9645
rect 24673 9605 24685 9639
rect 24719 9636 24731 9639
rect 24719 9608 27108 9636
rect 24719 9605 24731 9608
rect 24673 9599 24731 9605
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23201 9571 23259 9577
rect 23201 9568 23213 9571
rect 22796 9540 23213 9568
rect 22796 9528 22802 9540
rect 23201 9537 23213 9540
rect 23247 9537 23259 9571
rect 23382 9568 23388 9580
rect 23343 9540 23388 9568
rect 23201 9531 23259 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 24121 9571 24179 9577
rect 24121 9537 24133 9571
rect 24167 9568 24179 9571
rect 24486 9568 24492 9580
rect 24167 9540 24492 9568
rect 24167 9537 24179 9540
rect 24121 9531 24179 9537
rect 24486 9528 24492 9540
rect 24544 9568 24550 9580
rect 24688 9568 24716 9599
rect 24544 9540 24716 9568
rect 24544 9528 24550 9540
rect 25406 9528 25412 9580
rect 25464 9568 25470 9580
rect 25501 9571 25559 9577
rect 25501 9568 25513 9571
rect 25464 9540 25513 9568
rect 25464 9528 25470 9540
rect 25501 9537 25513 9540
rect 25547 9537 25559 9571
rect 25501 9531 25559 9537
rect 25590 9528 25596 9580
rect 25648 9568 25654 9580
rect 25777 9571 25835 9577
rect 25777 9568 25789 9571
rect 25648 9540 25789 9568
rect 25648 9528 25654 9540
rect 25777 9537 25789 9540
rect 25823 9537 25835 9571
rect 27080 9568 27108 9608
rect 27246 9596 27252 9648
rect 27304 9636 27310 9648
rect 27709 9639 27767 9645
rect 27709 9636 27721 9639
rect 27304 9608 27721 9636
rect 27304 9596 27310 9608
rect 27709 9605 27721 9608
rect 27755 9636 27767 9639
rect 28353 9639 28411 9645
rect 28353 9636 28365 9639
rect 27755 9608 28365 9636
rect 27755 9605 27767 9608
rect 27709 9599 27767 9605
rect 28353 9605 28365 9608
rect 28399 9605 28411 9639
rect 28353 9599 28411 9605
rect 31294 9596 31300 9648
rect 31352 9636 31358 9648
rect 31573 9639 31631 9645
rect 31573 9636 31585 9639
rect 31352 9608 31585 9636
rect 31352 9596 31358 9608
rect 31573 9605 31585 9608
rect 31619 9605 31631 9639
rect 31573 9599 31631 9605
rect 32582 9596 32588 9648
rect 32640 9636 32646 9648
rect 33137 9639 33195 9645
rect 33137 9636 33149 9639
rect 32640 9608 33149 9636
rect 32640 9596 32646 9608
rect 33137 9605 33149 9608
rect 33183 9636 33195 9639
rect 33689 9639 33747 9645
rect 33689 9636 33701 9639
rect 33183 9608 33701 9636
rect 33183 9605 33195 9608
rect 33137 9599 33195 9605
rect 33689 9605 33701 9608
rect 33735 9605 33747 9639
rect 33689 9599 33747 9605
rect 28626 9568 28632 9580
rect 27080 9540 28632 9568
rect 25777 9531 25835 9537
rect 28626 9528 28632 9540
rect 28684 9528 28690 9580
rect 30650 9568 30656 9580
rect 30611 9540 30656 9568
rect 30650 9528 30656 9540
rect 30708 9528 30714 9580
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9568 31447 9571
rect 31754 9568 31760 9580
rect 31435 9540 31760 9568
rect 31435 9537 31447 9540
rect 31389 9531 31447 9537
rect 31754 9528 31760 9540
rect 31812 9528 31818 9580
rect 34606 9528 34612 9580
rect 34664 9568 34670 9580
rect 35161 9571 35219 9577
rect 35161 9568 35173 9571
rect 34664 9540 35173 9568
rect 34664 9528 34670 9540
rect 35161 9537 35173 9540
rect 35207 9537 35219 9571
rect 35161 9531 35219 9537
rect 35802 9528 35808 9580
rect 35860 9568 35866 9580
rect 36725 9571 36783 9577
rect 36725 9568 36737 9571
rect 35860 9540 36737 9568
rect 35860 9528 35866 9540
rect 36725 9537 36737 9540
rect 36771 9537 36783 9571
rect 37274 9568 37280 9580
rect 37235 9540 37280 9568
rect 36725 9531 36783 9537
rect 37274 9528 37280 9540
rect 37332 9528 37338 9580
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 22925 9503 22983 9509
rect 22925 9500 22937 9503
rect 22336 9472 22937 9500
rect 22336 9460 22342 9472
rect 22925 9469 22937 9472
rect 22971 9469 22983 9503
rect 37550 9500 37556 9512
rect 22925 9463 22983 9469
rect 23032 9472 31754 9500
rect 37511 9472 37556 9500
rect 23032 9432 23060 9472
rect 22066 9404 23060 9432
rect 31726 9432 31754 9472
rect 37550 9460 37556 9472
rect 37608 9460 37614 9512
rect 37366 9432 37372 9444
rect 31726 9404 37372 9432
rect 37366 9392 37372 9404
rect 37424 9392 37430 9444
rect 15194 9364 15200 9376
rect 13280 9336 15200 9364
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18785 9367 18843 9373
rect 18785 9364 18797 9367
rect 17828 9336 18797 9364
rect 17828 9324 17834 9336
rect 18785 9333 18797 9336
rect 18831 9333 18843 9367
rect 18785 9327 18843 9333
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 19116 9336 19257 9364
rect 19116 9324 19122 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 20257 9367 20315 9373
rect 20257 9364 20269 9367
rect 19392 9336 20269 9364
rect 19392 9324 19398 9336
rect 20257 9333 20269 9336
rect 20303 9364 20315 9367
rect 22002 9364 22008 9376
rect 20303 9336 22008 9364
rect 20303 9333 20315 9336
rect 20257 9327 20315 9333
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 22094 9324 22100 9376
rect 22152 9364 22158 9376
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22152 9336 23029 9364
rect 22152 9324 22158 9336
rect 23017 9333 23029 9336
rect 23063 9364 23075 9367
rect 25498 9364 25504 9376
rect 23063 9336 25504 9364
rect 23063 9333 23075 9336
rect 23017 9327 23075 9333
rect 25498 9324 25504 9336
rect 25556 9364 25562 9376
rect 25593 9367 25651 9373
rect 25593 9364 25605 9367
rect 25556 9336 25605 9364
rect 25556 9324 25562 9336
rect 25593 9333 25605 9336
rect 25639 9333 25651 9367
rect 25593 9327 25651 9333
rect 25961 9367 26019 9373
rect 25961 9333 25973 9367
rect 26007 9364 26019 9367
rect 26050 9364 26056 9376
rect 26007 9336 26056 9364
rect 26007 9333 26019 9336
rect 25961 9327 26019 9333
rect 26050 9324 26056 9336
rect 26108 9324 26114 9376
rect 28445 9367 28503 9373
rect 28445 9333 28457 9367
rect 28491 9364 28503 9367
rect 30282 9364 30288 9376
rect 28491 9336 30288 9364
rect 28491 9333 28503 9336
rect 28445 9327 28503 9333
rect 30282 9324 30288 9336
rect 30340 9324 30346 9376
rect 33781 9367 33839 9373
rect 33781 9333 33793 9367
rect 33827 9364 33839 9367
rect 34514 9364 34520 9376
rect 33827 9336 34520 9364
rect 33827 9333 33839 9336
rect 33781 9327 33839 9333
rect 34514 9324 34520 9336
rect 34572 9324 34578 9376
rect 35345 9367 35403 9373
rect 35345 9333 35357 9367
rect 35391 9364 35403 9367
rect 35434 9364 35440 9376
rect 35391 9336 35440 9364
rect 35391 9333 35403 9336
rect 35345 9327 35403 9333
rect 35434 9324 35440 9336
rect 35492 9324 35498 9376
rect 36495 9367 36553 9373
rect 36495 9333 36507 9367
rect 36541 9364 36553 9367
rect 38010 9364 38016 9376
rect 36541 9336 38016 9364
rect 36541 9333 36553 9336
rect 36495 9327 36553 9333
rect 38010 9324 38016 9336
rect 38068 9324 38074 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 2501 9163 2559 9169
rect 2501 9160 2513 9163
rect 2372 9132 2513 9160
rect 2372 9120 2378 9132
rect 2501 9129 2513 9132
rect 2547 9129 2559 9163
rect 2501 9123 2559 9129
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3694 9160 3700 9172
rect 3007 9132 3700 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 7006 9160 7012 9172
rect 6656 9132 7012 9160
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 1636 9064 2820 9092
rect 1636 9052 1642 9064
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2792 8965 2820 9064
rect 6656 9033 6684 9132
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 22370 9160 22376 9172
rect 7432 9132 22376 9160
rect 7432 9120 7438 9132
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 22738 9160 22744 9172
rect 22699 9132 22744 9160
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 25501 9163 25559 9169
rect 25501 9129 25513 9163
rect 25547 9160 25559 9163
rect 25590 9160 25596 9172
rect 25547 9132 25596 9160
rect 25547 9129 25559 9132
rect 25501 9123 25559 9129
rect 25590 9120 25596 9132
rect 25648 9120 25654 9172
rect 27341 9163 27399 9169
rect 27341 9160 27353 9163
rect 25700 9132 27353 9160
rect 11057 9095 11115 9101
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 12066 9092 12072 9104
rect 11103 9064 12072 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 12526 9092 12532 9104
rect 12216 9064 12532 9092
rect 12216 9052 12222 9064
rect 12526 9052 12532 9064
rect 12584 9092 12590 9104
rect 13262 9092 13268 9104
rect 12584 9064 13268 9092
rect 12584 9052 12590 9064
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 18230 9052 18236 9104
rect 18288 9092 18294 9104
rect 18417 9095 18475 9101
rect 18417 9092 18429 9095
rect 18288 9064 18429 9092
rect 18288 9052 18294 9064
rect 18417 9061 18429 9064
rect 18463 9061 18475 9095
rect 19242 9092 19248 9104
rect 19203 9064 19248 9092
rect 18417 9055 18475 9061
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 20438 9092 20444 9104
rect 20399 9064 20444 9092
rect 20438 9052 20444 9064
rect 20496 9052 20502 9104
rect 22002 9052 22008 9104
rect 22060 9092 22066 9104
rect 22060 9064 23244 9092
rect 22060 9052 22066 9064
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 9024 11207 9027
rect 12176 9024 12204 9052
rect 11195 8996 12204 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 3786 8956 3792 8968
rect 3699 8928 3792 8956
rect 2777 8919 2835 8925
rect 3786 8916 3792 8928
rect 3844 8956 3850 8968
rect 6656 8956 6684 8987
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 12308 8996 12353 9024
rect 12308 8984 12314 8996
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 14921 9027 14979 9033
rect 14921 9024 14933 9027
rect 14792 8996 14933 9024
rect 14792 8984 14798 8996
rect 14921 8993 14933 8996
rect 14967 8993 14979 9027
rect 21361 9027 21419 9033
rect 14921 8987 14979 8993
rect 17972 8996 19748 9024
rect 17972 8968 18000 8996
rect 9582 8956 9588 8968
rect 3844 8928 6684 8956
rect 6840 8928 9588 8956
rect 3844 8916 3850 8928
rect 4062 8897 4068 8900
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 2041 8891 2099 8897
rect 1719 8860 1808 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 1780 8820 1808 8860
rect 2041 8857 2053 8891
rect 2087 8888 2099 8891
rect 2087 8860 2912 8888
rect 2087 8857 2099 8860
rect 2041 8851 2099 8857
rect 2774 8820 2780 8832
rect 1780 8792 2780 8820
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 2884 8820 2912 8860
rect 4056 8851 4068 8897
rect 4120 8888 4126 8900
rect 6840 8888 6868 8928
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 10962 8956 10968 8968
rect 10923 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11974 8956 11980 8968
rect 11287 8928 11980 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11974 8916 11980 8928
rect 12032 8956 12038 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 12032 8928 12081 8956
rect 12032 8916 12038 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 12069 8919 12127 8925
rect 12176 8928 12357 8956
rect 4120 8860 4156 8888
rect 4724 8860 6868 8888
rect 6908 8891 6966 8897
rect 4062 8848 4068 8851
rect 4120 8848 4126 8860
rect 4724 8820 4752 8860
rect 6908 8857 6920 8891
rect 6954 8888 6966 8891
rect 7098 8888 7104 8900
rect 6954 8860 7104 8888
rect 6954 8857 6966 8860
rect 6908 8851 6966 8857
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 9858 8888 9864 8900
rect 7208 8860 9864 8888
rect 2884 8792 4752 8820
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 4856 8792 5181 8820
rect 4856 8780 4862 8792
rect 5169 8789 5181 8792
rect 5215 8820 5227 8823
rect 7208 8820 7236 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 11330 8888 11336 8900
rect 10367 8860 11336 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 12176 8888 12204 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 13412 8928 14657 8956
rect 13412 8916 13418 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 16850 8916 16856 8968
rect 16908 8965 16914 8968
rect 16908 8956 16920 8965
rect 17126 8956 17132 8968
rect 16908 8928 16953 8956
rect 17087 8928 17132 8956
rect 16908 8919 16920 8928
rect 16908 8916 16914 8919
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8956 17831 8959
rect 17862 8956 17868 8968
rect 17819 8928 17868 8956
rect 17819 8925 17831 8928
rect 17773 8919 17831 8925
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18233 8959 18291 8965
rect 18012 8928 18057 8956
rect 18012 8916 18018 8928
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18279 8928 19441 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 19429 8925 19441 8928
rect 19475 8956 19487 8959
rect 19518 8956 19524 8968
rect 19475 8928 19524 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 19720 8965 19748 8996
rect 21361 8993 21373 9027
rect 21407 9024 21419 9027
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 21407 8996 22293 9024
rect 21407 8993 21419 8996
rect 21361 8987 21419 8993
rect 22281 8993 22293 8996
rect 22327 9024 22339 9027
rect 22462 9024 22468 9036
rect 22327 8996 22468 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20070 8956 20076 8968
rect 19935 8928 20076 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 21910 8916 21916 8968
rect 21968 8956 21974 8968
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21968 8928 22017 8956
rect 21968 8916 21974 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 22094 8916 22100 8968
rect 22152 8956 22158 8968
rect 22189 8959 22247 8965
rect 22189 8956 22201 8959
rect 22152 8928 22201 8956
rect 22152 8916 22158 8928
rect 22189 8925 22201 8928
rect 22235 8925 22247 8959
rect 22922 8956 22928 8968
rect 22883 8928 22928 8956
rect 22189 8919 22247 8925
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 23216 8965 23244 9064
rect 25130 9052 25136 9104
rect 25188 9092 25194 9104
rect 25700 9092 25728 9132
rect 27341 9129 27353 9132
rect 27387 9129 27399 9163
rect 27341 9123 27399 9129
rect 32122 9120 32128 9172
rect 32180 9160 32186 9172
rect 32309 9163 32367 9169
rect 32309 9160 32321 9163
rect 32180 9132 32321 9160
rect 32180 9120 32186 9132
rect 32309 9129 32321 9132
rect 32355 9160 32367 9163
rect 37458 9160 37464 9172
rect 32355 9132 37464 9160
rect 32355 9129 32367 9132
rect 32309 9123 32367 9129
rect 37458 9120 37464 9132
rect 37516 9120 37522 9172
rect 25188 9064 25728 9092
rect 25188 9052 25194 9064
rect 34698 9052 34704 9104
rect 34756 9092 34762 9104
rect 34977 9095 35035 9101
rect 34977 9092 34989 9095
rect 34756 9064 34989 9092
rect 34756 9052 34762 9064
rect 34977 9061 34989 9064
rect 35023 9061 35035 9095
rect 34977 9055 35035 9061
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 24636 8996 25360 9024
rect 24636 8984 24642 8996
rect 23201 8959 23259 8965
rect 23201 8925 23213 8959
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 23385 8959 23443 8965
rect 23385 8925 23397 8959
rect 23431 8956 23443 8959
rect 23474 8956 23480 8968
rect 23431 8928 23480 8956
rect 23431 8925 23443 8928
rect 23385 8919 23443 8925
rect 11756 8860 12204 8888
rect 12989 8891 13047 8897
rect 11756 8848 11762 8860
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13035 8860 17080 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 5215 8792 7236 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 7800 8792 8033 8820
rect 7800 8780 7806 8792
rect 8021 8789 8033 8792
rect 8067 8820 8079 8823
rect 8202 8820 8208 8832
rect 8067 8792 8208 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 10226 8820 10232 8832
rect 10187 8792 10232 8820
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 11422 8820 11428 8832
rect 11383 8792 11428 8820
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11848 8792 11897 8820
rect 11848 8780 11854 8792
rect 11885 8789 11897 8792
rect 11931 8789 11943 8823
rect 11885 8783 11943 8789
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 13004 8820 13032 8851
rect 12032 8792 13032 8820
rect 15749 8823 15807 8829
rect 12032 8780 12038 8792
rect 15749 8789 15761 8823
rect 15795 8820 15807 8823
rect 16390 8820 16396 8832
rect 15795 8792 16396 8820
rect 15795 8789 15807 8792
rect 15749 8783 15807 8789
rect 16390 8780 16396 8792
rect 16448 8820 16454 8832
rect 16942 8820 16948 8832
rect 16448 8792 16948 8820
rect 16448 8780 16454 8792
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17052 8820 17080 8860
rect 17218 8848 17224 8900
rect 17276 8888 17282 8900
rect 23216 8888 23244 8919
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 24854 8956 24860 8968
rect 24815 8928 24860 8956
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 25332 8965 25360 8996
rect 31754 8984 31760 9036
rect 31812 9024 31818 9036
rect 33137 9027 33195 9033
rect 33137 9024 33149 9027
rect 31812 8996 33149 9024
rect 31812 8984 31818 8996
rect 33137 8993 33149 8996
rect 33183 8993 33195 9027
rect 33137 8987 33195 8993
rect 25041 8959 25099 8965
rect 25041 8925 25053 8959
rect 25087 8925 25099 8959
rect 25041 8919 25099 8925
rect 25317 8959 25375 8965
rect 25317 8925 25329 8959
rect 25363 8956 25375 8959
rect 25590 8956 25596 8968
rect 25363 8928 25596 8956
rect 25363 8925 25375 8928
rect 25317 8919 25375 8925
rect 25056 8888 25084 8919
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 25958 8956 25964 8968
rect 25919 8928 25964 8956
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 26228 8959 26286 8965
rect 26228 8925 26240 8959
rect 26274 8925 26286 8959
rect 30650 8956 30656 8968
rect 30611 8928 30656 8956
rect 26228 8919 26286 8925
rect 25222 8888 25228 8900
rect 17276 8860 22094 8888
rect 23216 8860 25228 8888
rect 17276 8848 17282 8860
rect 20622 8820 20628 8832
rect 17052 8792 20628 8820
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 21818 8820 21824 8832
rect 21779 8792 21824 8820
rect 21818 8780 21824 8792
rect 21876 8780 21882 8832
rect 22066 8820 22094 8860
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 26142 8848 26148 8900
rect 26200 8888 26206 8900
rect 26252 8888 26280 8919
rect 30650 8916 30656 8928
rect 30708 8916 30714 8968
rect 31665 8959 31723 8965
rect 31665 8925 31677 8959
rect 31711 8956 31723 8959
rect 32122 8956 32128 8968
rect 31711 8928 32128 8956
rect 31711 8925 31723 8928
rect 31665 8919 31723 8925
rect 26200 8860 26280 8888
rect 26200 8848 26206 8860
rect 28626 8848 28632 8900
rect 28684 8888 28690 8900
rect 31680 8888 31708 8919
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 33413 8959 33471 8965
rect 33413 8925 33425 8959
rect 33459 8956 33471 8959
rect 34330 8956 34336 8968
rect 33459 8928 34336 8956
rect 33459 8925 33471 8928
rect 33413 8919 33471 8925
rect 34330 8916 34336 8928
rect 34388 8956 34394 8968
rect 34701 8959 34759 8965
rect 34701 8956 34713 8959
rect 34388 8928 34713 8956
rect 34388 8916 34394 8928
rect 34701 8925 34713 8928
rect 34747 8925 34759 8959
rect 34701 8919 34759 8925
rect 36081 8959 36139 8965
rect 36081 8925 36093 8959
rect 36127 8956 36139 8959
rect 36170 8956 36176 8968
rect 36127 8928 36176 8956
rect 36127 8925 36139 8928
rect 36081 8919 36139 8925
rect 36170 8916 36176 8928
rect 36228 8916 36234 8968
rect 38102 8956 38108 8968
rect 38063 8928 38108 8956
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 36354 8897 36360 8900
rect 28684 8860 31708 8888
rect 28684 8848 28690 8860
rect 36348 8851 36360 8897
rect 36412 8888 36418 8900
rect 36412 8860 36448 8888
rect 36354 8848 36360 8851
rect 36412 8848 36418 8860
rect 27246 8820 27252 8832
rect 22066 8792 27252 8820
rect 27246 8780 27252 8792
rect 27304 8780 27310 8832
rect 27982 8820 27988 8832
rect 27943 8792 27988 8820
rect 27982 8780 27988 8792
rect 28040 8780 28046 8832
rect 29730 8820 29736 8832
rect 29691 8792 29736 8820
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 30837 8823 30895 8829
rect 30837 8789 30849 8823
rect 30883 8820 30895 8823
rect 31018 8820 31024 8832
rect 30883 8792 31024 8820
rect 30883 8789 30895 8792
rect 30837 8783 30895 8789
rect 31018 8780 31024 8792
rect 31076 8780 31082 8832
rect 31573 8823 31631 8829
rect 31573 8789 31585 8823
rect 31619 8820 31631 8823
rect 31754 8820 31760 8832
rect 31619 8792 31760 8820
rect 31619 8789 31631 8792
rect 31573 8783 31631 8789
rect 31754 8780 31760 8792
rect 31812 8780 31818 8832
rect 35161 8823 35219 8829
rect 35161 8789 35173 8823
rect 35207 8820 35219 8823
rect 35802 8820 35808 8832
rect 35207 8792 35808 8820
rect 35207 8789 35219 8792
rect 35161 8783 35219 8789
rect 35802 8780 35808 8792
rect 35860 8780 35866 8832
rect 37461 8823 37519 8829
rect 37461 8789 37473 8823
rect 37507 8820 37519 8823
rect 37642 8820 37648 8832
rect 37507 8792 37648 8820
rect 37507 8789 37519 8792
rect 37461 8783 37519 8789
rect 37642 8780 37648 8792
rect 37700 8780 37706 8832
rect 37918 8820 37924 8832
rect 37879 8792 37924 8820
rect 37918 8780 37924 8792
rect 37976 8780 37982 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1486 8616 1492 8628
rect 1447 8588 1492 8616
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 4065 8619 4123 8625
rect 4065 8585 4077 8619
rect 4111 8616 4123 8619
rect 5350 8616 5356 8628
rect 4111 8588 5356 8616
rect 4111 8585 4123 8588
rect 4065 8579 4123 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5500 8588 5641 8616
rect 5500 8576 5506 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 5629 8579 5687 8585
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 25774 8616 25780 8628
rect 8536 8588 25636 8616
rect 25735 8588 25780 8616
rect 8536 8576 8542 8588
rect 3786 8548 3792 8560
rect 2700 8520 3792 8548
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2590 8480 2596 8492
rect 1719 8452 2596 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2700 8489 2728 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 5460 8548 5488 8576
rect 9125 8551 9183 8557
rect 4724 8520 5488 8548
rect 5552 8520 9076 8548
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2952 8483 3010 8489
rect 2952 8449 2964 8483
rect 2998 8480 3010 8483
rect 3326 8480 3332 8492
rect 2998 8452 3332 8480
rect 2998 8449 3010 8452
rect 2952 8443 3010 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 4724 8489 4752 8520
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4982 8480 4988 8492
rect 4943 8452 4988 8480
rect 4709 8443 4767 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5350 8480 5356 8492
rect 5215 8452 5356 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5552 8412 5580 8520
rect 7282 8480 7288 8492
rect 7243 8452 7288 8480
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 8205 8483 8263 8489
rect 7524 8452 7696 8480
rect 7524 8440 7530 8452
rect 5316 8384 5580 8412
rect 6641 8415 6699 8421
rect 5316 8372 5322 8384
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7558 8412 7564 8424
rect 6687 8384 7564 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7668 8412 7696 8452
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 8294 8480 8300 8492
rect 8251 8452 8300 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 9048 8480 9076 8520
rect 9125 8517 9137 8551
rect 9171 8548 9183 8551
rect 10226 8548 10232 8560
rect 9171 8520 10232 8548
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 11974 8508 11980 8560
rect 12032 8548 12038 8560
rect 12162 8551 12220 8557
rect 12162 8548 12174 8551
rect 12032 8520 12174 8548
rect 12032 8508 12038 8520
rect 12162 8517 12174 8520
rect 12208 8517 12220 8551
rect 12162 8511 12220 8517
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 12434 8557 12440 8560
rect 12391 8551 12440 8557
rect 12308 8520 12353 8548
rect 12308 8508 12314 8520
rect 12391 8517 12403 8551
rect 12437 8517 12440 8551
rect 12391 8511 12440 8517
rect 12434 8508 12440 8511
rect 12492 8508 12498 8560
rect 14277 8551 14335 8557
rect 14277 8517 14289 8551
rect 14323 8548 14335 8551
rect 17126 8548 17132 8560
rect 14323 8520 17132 8548
rect 14323 8517 14335 8520
rect 14277 8511 14335 8517
rect 17126 8508 17132 8520
rect 17184 8548 17190 8560
rect 21542 8548 21548 8560
rect 17184 8520 21548 8548
rect 17184 8508 17190 8520
rect 11054 8480 11060 8492
rect 8444 8452 8489 8480
rect 9048 8452 11060 8480
rect 8444 8440 8450 8452
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12894 8480 12900 8492
rect 12575 8452 12900 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13078 8480 13084 8492
rect 13039 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13354 8480 13360 8492
rect 13315 8452 13360 8480
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 18800 8489 18828 8520
rect 21542 8508 21548 8520
rect 21600 8508 21606 8560
rect 21910 8548 21916 8560
rect 21871 8520 21916 8548
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 22002 8508 22008 8560
rect 22060 8548 22066 8560
rect 23284 8551 23342 8557
rect 22060 8520 22416 8548
rect 22060 8508 22066 8520
rect 19058 8489 19064 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 19052 8480 19064 8489
rect 19019 8452 19064 8480
rect 18785 8443 18843 8449
rect 19052 8443 19064 8452
rect 8404 8412 8432 8440
rect 7668 8384 8432 8412
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 13262 8412 13268 8424
rect 8536 8384 8581 8412
rect 13223 8384 13268 8412
rect 8536 8372 8542 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 2133 8347 2191 8353
rect 2133 8344 2145 8347
rect 1636 8316 2145 8344
rect 1636 8304 1642 8316
rect 2133 8313 2145 8316
rect 2179 8313 2191 8347
rect 4525 8347 4583 8353
rect 4525 8344 4537 8347
rect 2133 8307 2191 8313
rect 3620 8316 4537 8344
rect 3620 8288 3648 8316
rect 4525 8313 4537 8316
rect 4571 8313 4583 8347
rect 4525 8307 4583 8313
rect 7006 8304 7012 8356
rect 7064 8344 7070 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 7064 8316 8953 8344
rect 7064 8304 7070 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 8941 8307 8999 8313
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10284 8316 12020 8344
rect 10284 8304 10290 8316
rect 3602 8236 3608 8288
rect 3660 8236 3666 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11885 8279 11943 8285
rect 11885 8276 11897 8279
rect 11112 8248 11897 8276
rect 11112 8236 11118 8248
rect 11885 8245 11897 8248
rect 11931 8245 11943 8279
rect 11992 8276 12020 8316
rect 12802 8304 12808 8356
rect 12860 8344 12866 8356
rect 12986 8344 12992 8356
rect 12860 8316 12992 8344
rect 12860 8304 12866 8316
rect 12986 8304 12992 8316
rect 13044 8344 13050 8356
rect 13173 8347 13231 8353
rect 13173 8344 13185 8347
rect 13044 8316 13185 8344
rect 13044 8304 13050 8316
rect 13173 8313 13185 8316
rect 13219 8313 13231 8347
rect 13538 8344 13544 8356
rect 13499 8316 13544 8344
rect 13173 8307 13231 8313
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 14108 8276 14136 8443
rect 19058 8440 19064 8443
rect 19116 8440 19122 8492
rect 22388 8489 22416 8520
rect 23284 8517 23296 8551
rect 23330 8548 23342 8551
rect 23382 8548 23388 8560
rect 23330 8520 23388 8548
rect 23330 8517 23342 8520
rect 23284 8511 23342 8517
rect 23382 8508 23388 8520
rect 23440 8508 23446 8560
rect 25608 8548 25636 8588
rect 25774 8576 25780 8588
rect 25832 8576 25838 8628
rect 27246 8576 27252 8628
rect 27304 8616 27310 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 27304 8588 27353 8616
rect 27304 8576 27310 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 29730 8616 29736 8628
rect 27341 8579 27399 8585
rect 27448 8588 29736 8616
rect 27448 8548 27476 8588
rect 29730 8576 29736 8588
rect 29788 8616 29794 8628
rect 30285 8619 30343 8625
rect 30285 8616 30297 8619
rect 29788 8588 30297 8616
rect 29788 8576 29794 8588
rect 30285 8585 30297 8588
rect 30331 8616 30343 8619
rect 34054 8616 34060 8628
rect 30331 8588 34060 8616
rect 30331 8585 30343 8588
rect 30285 8579 30343 8585
rect 34054 8576 34060 8588
rect 34112 8576 34118 8628
rect 34425 8619 34483 8625
rect 34425 8585 34437 8619
rect 34471 8616 34483 8619
rect 36722 8616 36728 8628
rect 34471 8588 36728 8616
rect 34471 8585 34483 8588
rect 34425 8579 34483 8585
rect 36722 8576 36728 8588
rect 36780 8576 36786 8628
rect 37366 8616 37372 8628
rect 37327 8588 37372 8616
rect 37366 8576 37372 8588
rect 37424 8576 37430 8628
rect 25608 8520 27476 8548
rect 27525 8551 27583 8557
rect 27525 8517 27537 8551
rect 27571 8548 27583 8551
rect 30377 8551 30435 8557
rect 30377 8548 30389 8551
rect 27571 8520 30389 8548
rect 27571 8517 27583 8520
rect 27525 8511 27583 8517
rect 30377 8517 30389 8520
rect 30423 8548 30435 8551
rect 32306 8548 32312 8560
rect 30423 8520 32312 8548
rect 30423 8517 30435 8520
rect 30377 8511 30435 8517
rect 32306 8508 32312 8520
rect 32364 8508 32370 8560
rect 36170 8548 36176 8560
rect 35360 8520 36176 8548
rect 35360 8492 35388 8520
rect 36170 8508 36176 8520
rect 36228 8508 36234 8560
rect 37734 8548 37740 8560
rect 37695 8520 37740 8548
rect 37734 8508 37740 8520
rect 37792 8508 37798 8560
rect 22122 8483 22180 8489
rect 22122 8449 22134 8483
rect 22168 8480 22180 8483
rect 22373 8483 22431 8489
rect 22168 8452 22324 8480
rect 22168 8449 22180 8452
rect 22122 8443 22180 8449
rect 20070 8304 20076 8356
rect 20128 8344 20134 8356
rect 20165 8347 20223 8353
rect 20165 8344 20177 8347
rect 20128 8316 20177 8344
rect 20128 8304 20134 8316
rect 20165 8313 20177 8316
rect 20211 8313 20223 8347
rect 20165 8307 20223 8313
rect 21269 8347 21327 8353
rect 21269 8313 21281 8347
rect 21315 8344 21327 8347
rect 22094 8344 22100 8356
rect 21315 8316 22100 8344
rect 21315 8313 21327 8316
rect 21269 8307 21327 8313
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 22296 8344 22324 8452
rect 22373 8449 22385 8483
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 22474 8483 22532 8489
rect 22474 8449 22486 8483
rect 22520 8449 22532 8483
rect 25130 8480 25136 8492
rect 25091 8452 25136 8480
rect 22474 8443 22532 8449
rect 22480 8412 22508 8443
rect 25130 8440 25136 8452
rect 25188 8440 25194 8492
rect 25222 8440 25228 8492
rect 25280 8480 25286 8492
rect 25317 8483 25375 8489
rect 25317 8480 25329 8483
rect 25280 8452 25329 8480
rect 25280 8440 25286 8452
rect 25317 8449 25329 8452
rect 25363 8449 25375 8483
rect 25590 8480 25596 8492
rect 25551 8452 25596 8480
rect 25317 8443 25375 8449
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 27706 8480 27712 8492
rect 27667 8452 27712 8480
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 34517 8483 34575 8489
rect 34517 8449 34529 8483
rect 34563 8449 34575 8483
rect 35342 8480 35348 8492
rect 35255 8452 35348 8480
rect 34517 8443 34575 8449
rect 22554 8412 22560 8424
rect 22480 8384 22560 8412
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 23017 8415 23075 8421
rect 23017 8381 23029 8415
rect 23063 8381 23075 8415
rect 23017 8375 23075 8381
rect 22922 8344 22928 8356
rect 22296 8316 22928 8344
rect 22922 8304 22928 8316
rect 22980 8304 22986 8356
rect 11992 8248 14136 8276
rect 11885 8239 11943 8245
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 23032 8276 23060 8375
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 27430 8412 27436 8424
rect 24912 8384 27436 8412
rect 24912 8372 24918 8384
rect 27430 8372 27436 8384
rect 27488 8372 27494 8424
rect 27982 8372 27988 8424
rect 28040 8412 28046 8424
rect 28169 8415 28227 8421
rect 28169 8412 28181 8415
rect 28040 8384 28181 8412
rect 28040 8372 28046 8384
rect 28169 8381 28181 8384
rect 28215 8381 28227 8415
rect 28169 8375 28227 8381
rect 28445 8415 28503 8421
rect 28445 8381 28457 8415
rect 28491 8412 28503 8415
rect 30006 8412 30012 8424
rect 28491 8384 30012 8412
rect 28491 8381 28503 8384
rect 28445 8375 28503 8381
rect 30006 8372 30012 8384
rect 30064 8372 30070 8424
rect 30282 8372 30288 8424
rect 30340 8412 30346 8424
rect 30469 8415 30527 8421
rect 30469 8412 30481 8415
rect 30340 8384 30481 8412
rect 30340 8372 30346 8384
rect 30469 8381 30481 8384
rect 30515 8381 30527 8415
rect 30469 8375 30527 8381
rect 34333 8415 34391 8421
rect 34333 8381 34345 8415
rect 34379 8412 34391 8415
rect 34422 8412 34428 8424
rect 34379 8384 34428 8412
rect 34379 8381 34391 8384
rect 34333 8375 34391 8381
rect 34422 8372 34428 8384
rect 34480 8372 34486 8424
rect 24397 8347 24455 8353
rect 24397 8344 24409 8347
rect 23952 8316 24409 8344
rect 21600 8248 23060 8276
rect 21600 8236 21606 8248
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 23952 8276 23980 8316
rect 24397 8313 24409 8316
rect 24443 8313 24455 8347
rect 24397 8307 24455 8313
rect 25958 8304 25964 8356
rect 26016 8344 26022 8356
rect 29546 8344 29552 8356
rect 26016 8316 29552 8344
rect 26016 8304 26022 8316
rect 29546 8304 29552 8316
rect 29604 8304 29610 8356
rect 33594 8344 33600 8356
rect 33555 8316 33600 8344
rect 33594 8304 33600 8316
rect 33652 8344 33658 8356
rect 34532 8344 34560 8443
rect 35342 8440 35348 8452
rect 35400 8440 35406 8492
rect 35434 8440 35440 8492
rect 35492 8480 35498 8492
rect 37550 8489 37556 8492
rect 35601 8483 35659 8489
rect 35601 8480 35613 8483
rect 35492 8452 35613 8480
rect 35492 8440 35498 8452
rect 35601 8449 35613 8452
rect 35647 8449 35659 8483
rect 37548 8480 37556 8489
rect 37511 8452 37556 8480
rect 35601 8443 35659 8449
rect 37548 8443 37556 8452
rect 37550 8440 37556 8443
rect 37608 8440 37614 8492
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 37918 8480 37924 8492
rect 37700 8452 37745 8480
rect 37879 8452 37924 8480
rect 37700 8440 37706 8452
rect 37918 8440 37924 8452
rect 37976 8440 37982 8492
rect 38010 8440 38016 8492
rect 38068 8480 38074 8492
rect 38068 8452 38113 8480
rect 38068 8440 38074 8452
rect 33652 8316 34560 8344
rect 33652 8304 33658 8316
rect 23440 8248 23980 8276
rect 29917 8279 29975 8285
rect 23440 8236 23446 8248
rect 29917 8245 29929 8279
rect 29963 8276 29975 8279
rect 30098 8276 30104 8288
rect 29963 8248 30104 8276
rect 29963 8245 29975 8248
rect 29917 8239 29975 8245
rect 30098 8236 30104 8248
rect 30156 8236 30162 8288
rect 34790 8236 34796 8288
rect 34848 8276 34854 8288
rect 34885 8279 34943 8285
rect 34885 8276 34897 8279
rect 34848 8248 34897 8276
rect 34848 8236 34854 8248
rect 34885 8245 34897 8248
rect 34931 8245 34943 8279
rect 34885 8239 34943 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2866 8072 2872 8084
rect 2823 8044 2872 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 11054 8072 11060 8084
rect 2976 8044 11060 8072
rect 2976 8004 3004 8044
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12618 8072 12624 8084
rect 12579 8044 12624 8072
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13078 8072 13084 8084
rect 13039 8044 13084 8072
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 17402 8072 17408 8084
rect 16623 8044 17408 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 25792 8044 32720 8072
rect 2746 7976 3004 8004
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1688 7800 1716 7831
rect 2746 7800 2774 7976
rect 4614 7964 4620 8016
rect 4672 7964 4678 8016
rect 5353 8007 5411 8013
rect 5353 7973 5365 8007
rect 5399 8004 5411 8007
rect 5442 8004 5448 8016
rect 5399 7976 5448 8004
rect 5399 7973 5411 7976
rect 5353 7967 5411 7973
rect 4632 7936 4660 7964
rect 4982 7936 4988 7948
rect 2976 7908 4660 7936
rect 4724 7908 4988 7936
rect 2976 7877 3004 7908
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 3142 7868 3148 7880
rect 3103 7840 3148 7868
rect 2961 7831 3019 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4724 7868 4752 7908
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 4663 7840 4752 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 1688 7772 2774 7800
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 2225 7735 2283 7741
rect 2225 7732 2237 7735
rect 1820 7704 2237 7732
rect 1820 7692 1826 7704
rect 2225 7701 2237 7704
rect 2271 7732 2283 7735
rect 3252 7732 3280 7831
rect 4356 7800 4384 7831
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 5258 7868 5264 7880
rect 4856 7840 5264 7868
rect 4856 7828 4862 7840
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5368 7800 5396 7967
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 12406 7976 12940 8004
rect 12406 7936 12434 7976
rect 5460 7908 12434 7936
rect 5460 7880 5488 7908
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 11572 7840 12633 7868
rect 11572 7828 11578 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12621 7831 12679 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 12912 7877 12940 7976
rect 21450 7896 21456 7948
rect 21508 7936 21514 7948
rect 25792 7936 25820 8044
rect 27982 8004 27988 8016
rect 26988 7976 27988 8004
rect 21508 7908 21680 7936
rect 21508 7896 21514 7908
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 21542 7868 21548 7880
rect 21503 7840 21548 7868
rect 12897 7831 12955 7837
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 21652 7868 21680 7908
rect 25608 7908 25820 7936
rect 25608 7868 25636 7908
rect 25958 7896 25964 7948
rect 26016 7936 26022 7948
rect 26016 7908 26061 7936
rect 26016 7896 26022 7908
rect 21652 7840 25636 7868
rect 26050 7828 26056 7880
rect 26108 7868 26114 7880
rect 26217 7871 26275 7877
rect 26217 7868 26229 7871
rect 26108 7840 26229 7868
rect 26108 7828 26114 7840
rect 26217 7837 26229 7840
rect 26263 7837 26275 7871
rect 26988 7868 27016 7976
rect 27982 7964 27988 7976
rect 28040 7964 28046 8016
rect 28626 8004 28632 8016
rect 28587 7976 28632 8004
rect 28626 7964 28632 7976
rect 28684 7964 28690 8016
rect 30098 8004 30104 8016
rect 30059 7976 30104 8004
rect 30098 7964 30104 7976
rect 30156 7964 30162 8016
rect 30285 8007 30343 8013
rect 30285 7973 30297 8007
rect 30331 8004 30343 8007
rect 30650 8004 30656 8016
rect 30331 7976 30656 8004
rect 30331 7973 30343 7976
rect 30285 7967 30343 7973
rect 30650 7964 30656 7976
rect 30708 7964 30714 8016
rect 32306 8004 32312 8016
rect 32267 7976 32312 8004
rect 32306 7964 32312 7976
rect 32364 7964 32370 8016
rect 32692 8004 32720 8044
rect 32766 8032 32772 8084
rect 32824 8072 32830 8084
rect 32861 8075 32919 8081
rect 32861 8072 32873 8075
rect 32824 8044 32873 8072
rect 32824 8032 32830 8044
rect 32861 8041 32873 8044
rect 32907 8072 32919 8075
rect 35342 8072 35348 8084
rect 32907 8044 35348 8072
rect 32907 8041 32919 8044
rect 32861 8035 32919 8041
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 36081 8075 36139 8081
rect 36081 8041 36093 8075
rect 36127 8072 36139 8075
rect 36354 8072 36360 8084
rect 36127 8044 36360 8072
rect 36127 8041 36139 8044
rect 36081 8035 36139 8041
rect 36354 8032 36360 8044
rect 36412 8032 36418 8084
rect 38010 8072 38016 8084
rect 37971 8044 38016 8072
rect 38010 8032 38016 8044
rect 38068 8032 38074 8084
rect 38930 8004 38936 8016
rect 32692 7976 38936 8004
rect 38930 7964 38936 7976
rect 38988 7964 38994 8016
rect 26217 7831 26275 7837
rect 26344 7840 27016 7868
rect 27801 7871 27859 7877
rect 4356 7772 5396 7800
rect 7834 7760 7840 7812
rect 7892 7800 7898 7812
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 7892 7772 9321 7800
rect 7892 7760 7898 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 9493 7803 9551 7809
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 10137 7803 10195 7809
rect 10137 7800 10149 7803
rect 9539 7772 10149 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 10137 7769 10149 7772
rect 10183 7800 10195 7803
rect 18966 7800 18972 7812
rect 10183 7772 18972 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 21818 7809 21824 7812
rect 21812 7800 21824 7809
rect 21779 7772 21824 7800
rect 21812 7763 21824 7772
rect 21818 7760 21824 7763
rect 21876 7760 21882 7812
rect 26344 7800 26372 7840
rect 27801 7837 27813 7871
rect 27847 7868 27859 7871
rect 28644 7868 28672 7964
rect 29825 7939 29883 7945
rect 29825 7905 29837 7939
rect 29871 7936 29883 7939
rect 30006 7936 30012 7948
rect 29871 7908 30012 7936
rect 29871 7905 29883 7908
rect 29825 7899 29883 7905
rect 30006 7896 30012 7908
rect 30064 7896 30070 7948
rect 34054 7936 34060 7948
rect 34015 7908 34060 7936
rect 34054 7896 34060 7908
rect 34112 7936 34118 7948
rect 35253 7939 35311 7945
rect 34112 7908 35112 7936
rect 34112 7896 34118 7908
rect 27847 7840 28672 7868
rect 27847 7837 27859 7840
rect 27801 7831 27859 7837
rect 30834 7828 30840 7880
rect 30892 7868 30898 7880
rect 30929 7871 30987 7877
rect 30929 7868 30941 7871
rect 30892 7840 30941 7868
rect 30892 7828 30898 7840
rect 30929 7837 30941 7840
rect 30975 7837 30987 7871
rect 30929 7831 30987 7837
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 35084 7877 35112 7908
rect 35253 7905 35265 7939
rect 35299 7905 35311 7939
rect 35253 7899 35311 7905
rect 37369 7939 37427 7945
rect 37369 7905 37381 7939
rect 37415 7936 37427 7939
rect 38102 7936 38108 7948
rect 37415 7908 38108 7936
rect 37415 7905 37427 7908
rect 37369 7899 37427 7905
rect 31185 7871 31243 7877
rect 31185 7868 31197 7871
rect 31076 7840 31197 7868
rect 31076 7828 31082 7840
rect 31185 7837 31197 7840
rect 31231 7837 31243 7871
rect 31185 7831 31243 7837
rect 35069 7871 35127 7877
rect 35069 7837 35081 7871
rect 35115 7837 35127 7871
rect 35069 7831 35127 7837
rect 22480 7772 26372 7800
rect 2271 7704 3280 7732
rect 4157 7735 4215 7741
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 4157 7701 4169 7735
rect 4203 7732 4215 7735
rect 4430 7732 4436 7744
rect 4203 7704 4436 7732
rect 4203 7701 4215 7704
rect 4157 7695 4215 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 7926 7732 7932 7744
rect 7887 7704 7932 7732
rect 7926 7692 7932 7704
rect 7984 7732 7990 7744
rect 8478 7732 8484 7744
rect 7984 7704 8484 7732
rect 7984 7692 7990 7704
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 22480 7732 22508 7772
rect 34514 7760 34520 7812
rect 34572 7800 34578 7812
rect 35268 7800 35296 7899
rect 38102 7896 38108 7908
rect 38160 7896 38166 7948
rect 35802 7828 35808 7880
rect 35860 7868 35866 7880
rect 35897 7871 35955 7877
rect 35897 7868 35909 7871
rect 35860 7840 35909 7868
rect 35860 7828 35866 7840
rect 35897 7837 35909 7840
rect 35943 7837 35955 7871
rect 35897 7831 35955 7837
rect 36722 7828 36728 7880
rect 36780 7868 36786 7880
rect 37182 7868 37188 7880
rect 36780 7840 37188 7868
rect 36780 7828 36786 7840
rect 37182 7828 37188 7840
rect 37240 7868 37246 7880
rect 37829 7871 37887 7877
rect 37829 7868 37841 7871
rect 37240 7840 37841 7868
rect 37240 7828 37246 7840
rect 37829 7837 37841 7840
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 34572 7772 35296 7800
rect 34572 7760 34578 7772
rect 20036 7704 22508 7732
rect 20036 7692 20042 7704
rect 22554 7692 22560 7744
rect 22612 7732 22618 7744
rect 22925 7735 22983 7741
rect 22925 7732 22937 7735
rect 22612 7704 22937 7732
rect 22612 7692 22618 7704
rect 22925 7701 22937 7704
rect 22971 7732 22983 7735
rect 23385 7735 23443 7741
rect 23385 7732 23397 7735
rect 22971 7704 23397 7732
rect 22971 7701 22983 7704
rect 22925 7695 22983 7701
rect 23385 7701 23397 7704
rect 23431 7701 23443 7735
rect 23385 7695 23443 7701
rect 27341 7735 27399 7741
rect 27341 7701 27353 7735
rect 27387 7732 27399 7735
rect 27430 7732 27436 7744
rect 27387 7704 27436 7732
rect 27387 7701 27399 7704
rect 27341 7695 27399 7701
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 34698 7732 34704 7744
rect 34659 7704 34704 7732
rect 34698 7692 34704 7704
rect 34756 7692 34762 7744
rect 35161 7735 35219 7741
rect 35161 7701 35173 7735
rect 35207 7732 35219 7735
rect 37642 7732 37648 7744
rect 35207 7704 37648 7732
rect 35207 7701 35219 7704
rect 35161 7695 35219 7701
rect 37642 7692 37648 7704
rect 37700 7692 37706 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 3326 7528 3332 7540
rect 3287 7500 3332 7528
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4249 7531 4307 7537
rect 4249 7528 4261 7531
rect 4120 7500 4261 7528
rect 4120 7488 4126 7500
rect 4249 7497 4261 7500
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 6917 7531 6975 7537
rect 6917 7528 6929 7531
rect 4580 7500 6929 7528
rect 4580 7488 4586 7500
rect 6917 7497 6929 7500
rect 6963 7528 6975 7531
rect 7926 7528 7932 7540
rect 6963 7500 7932 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 19334 7528 19340 7540
rect 9784 7500 19340 7528
rect 6365 7463 6423 7469
rect 6365 7460 6377 7463
rect 1412 7432 6377 7460
rect 1412 7404 1440 7432
rect 6365 7429 6377 7432
rect 6411 7429 6423 7463
rect 6365 7423 6423 7429
rect 1394 7392 1400 7404
rect 1307 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3602 7392 3608 7404
rect 3559 7364 3608 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3712 7364 3801 7392
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 3712 7324 3740 7364
rect 3789 7361 3801 7364
rect 3835 7392 3847 7395
rect 4062 7392 4068 7404
rect 3835 7364 4068 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 7466 7392 7472 7404
rect 4672 7364 7472 7392
rect 4672 7352 4678 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 7834 7392 7840 7404
rect 7795 7364 7840 7392
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 9784 7401 9812 7500
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 22649 7531 22707 7537
rect 22649 7497 22661 7531
rect 22695 7528 22707 7531
rect 22922 7528 22928 7540
rect 22695 7500 22928 7528
rect 22695 7497 22707 7500
rect 22649 7491 22707 7497
rect 22922 7488 22928 7500
rect 22980 7488 22986 7540
rect 33594 7528 33600 7540
rect 30208 7500 33600 7528
rect 30208 7469 30236 7500
rect 33594 7488 33600 7500
rect 33652 7488 33658 7540
rect 34606 7488 34612 7540
rect 34664 7528 34670 7540
rect 34885 7531 34943 7537
rect 34885 7528 34897 7531
rect 34664 7500 34897 7528
rect 34664 7488 34670 7500
rect 34885 7497 34897 7500
rect 34931 7497 34943 7531
rect 35342 7528 35348 7540
rect 35303 7500 35348 7528
rect 34885 7491 34943 7497
rect 35342 7488 35348 7500
rect 35400 7528 35406 7540
rect 35802 7528 35808 7540
rect 35400 7500 35808 7528
rect 35400 7488 35406 7500
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 36078 7488 36084 7540
rect 36136 7528 36142 7540
rect 36265 7531 36323 7537
rect 36265 7528 36277 7531
rect 36136 7500 36277 7528
rect 36136 7488 36142 7500
rect 36265 7497 36277 7500
rect 36311 7497 36323 7531
rect 36265 7491 36323 7497
rect 29273 7463 29331 7469
rect 29273 7460 29285 7463
rect 12406 7432 29285 7460
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 2915 7296 3740 7324
rect 4709 7327 4767 7333
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 4798 7324 4804 7336
rect 4755 7296 4804 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 7926 7324 7932 7336
rect 7887 7296 7932 7324
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 8444 7296 9505 7324
rect 8444 7284 8450 7296
rect 9493 7293 9505 7296
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 4522 7256 4528 7268
rect 1627 7228 4528 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 4522 7216 4528 7228
rect 4580 7216 4586 7268
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 12406 7256 12434 7432
rect 29273 7429 29285 7432
rect 29319 7460 29331 7463
rect 30193 7463 30251 7469
rect 30193 7460 30205 7463
rect 29319 7432 30205 7460
rect 29319 7429 29331 7432
rect 29273 7423 29331 7429
rect 30193 7429 30205 7432
rect 30239 7429 30251 7463
rect 30193 7423 30251 7429
rect 30282 7420 30288 7472
rect 30340 7420 30346 7472
rect 34330 7420 34336 7472
rect 34388 7460 34394 7472
rect 34425 7463 34483 7469
rect 34425 7460 34437 7463
rect 34388 7432 34437 7460
rect 34388 7420 34394 7432
rect 34425 7429 34437 7432
rect 34471 7429 34483 7463
rect 34425 7423 34483 7429
rect 37182 7420 37188 7472
rect 37240 7460 37246 7472
rect 37645 7463 37703 7469
rect 37645 7460 37657 7463
rect 37240 7432 37657 7460
rect 37240 7420 37246 7432
rect 37645 7429 37657 7432
rect 37691 7429 37703 7463
rect 37645 7423 37703 7429
rect 37734 7420 37740 7472
rect 37792 7460 37798 7472
rect 37792 7432 37837 7460
rect 37792 7420 37798 7432
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15378 7392 15384 7404
rect 15243 7364 15384 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15838 7392 15844 7404
rect 15799 7364 15844 7392
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17402 7392 17408 7404
rect 17175 7364 17408 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7392 19579 7395
rect 19978 7392 19984 7404
rect 19567 7364 19984 7392
rect 19567 7361 19579 7364
rect 19521 7355 19579 7361
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 15396 7324 15424 7352
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15396 7296 16129 7324
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 19242 7324 19248 7336
rect 19203 7296 19248 7324
rect 16117 7287 16175 7293
rect 19242 7284 19248 7296
rect 19300 7284 19306 7336
rect 27724 7324 27752 7355
rect 27798 7352 27804 7404
rect 27856 7392 27862 7404
rect 27893 7395 27951 7401
rect 27893 7392 27905 7395
rect 27856 7364 27905 7392
rect 27856 7352 27862 7364
rect 27893 7361 27905 7364
rect 27939 7361 27951 7395
rect 30300 7392 30328 7420
rect 30300 7364 30420 7392
rect 27893 7355 27951 7361
rect 30282 7324 30288 7336
rect 27724 7296 30288 7324
rect 30282 7284 30288 7296
rect 30340 7284 30346 7336
rect 30392 7333 30420 7364
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 37550 7401 37556 7404
rect 31021 7395 31079 7401
rect 31021 7392 31033 7395
rect 30524 7364 31033 7392
rect 30524 7352 30530 7364
rect 31021 7361 31033 7364
rect 31067 7361 31079 7395
rect 37548 7392 37556 7401
rect 37511 7364 37556 7392
rect 31021 7355 31079 7361
rect 37548 7355 37556 7364
rect 37550 7352 37556 7355
rect 37608 7352 37614 7404
rect 37865 7395 37923 7401
rect 37865 7392 37877 7395
rect 37844 7361 37877 7392
rect 37911 7361 37923 7395
rect 37844 7355 37923 7361
rect 30377 7327 30435 7333
rect 30377 7293 30389 7327
rect 30423 7293 30435 7327
rect 30377 7287 30435 7293
rect 36630 7284 36636 7336
rect 36688 7324 36694 7336
rect 37844 7324 37872 7355
rect 38010 7352 38016 7404
rect 38068 7392 38074 7404
rect 38068 7364 38113 7392
rect 38068 7352 38074 7364
rect 36688 7296 37872 7324
rect 36688 7284 36694 7296
rect 7616 7228 12434 7256
rect 16025 7259 16083 7265
rect 7616 7216 7622 7228
rect 16025 7225 16037 7259
rect 16071 7256 16083 7259
rect 16758 7256 16764 7268
rect 16071 7228 16764 7256
rect 16071 7225 16083 7228
rect 16025 7219 16083 7225
rect 16758 7216 16764 7228
rect 16816 7256 16822 7268
rect 17037 7259 17095 7265
rect 17037 7256 17049 7259
rect 16816 7228 17049 7256
rect 16816 7216 16822 7228
rect 17037 7225 17049 7228
rect 17083 7225 17095 7259
rect 34790 7256 34796 7268
rect 34751 7228 34796 7256
rect 17037 7219 17095 7225
rect 34790 7216 34796 7228
rect 34848 7216 34854 7268
rect 37366 7256 37372 7268
rect 37327 7228 37372 7256
rect 37366 7216 37372 7228
rect 37424 7216 37430 7268
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3200 7160 3709 7188
rect 3200 7148 3206 7160
rect 3697 7157 3709 7160
rect 3743 7188 3755 7191
rect 4614 7188 4620 7200
rect 3743 7160 4620 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4948 7160 5273 7188
rect 4948 7148 4954 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5718 7188 5724 7200
rect 5679 7160 5724 7188
rect 5261 7151 5319 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 7340 7160 7481 7188
rect 7340 7148 7346 7160
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 7469 7151 7527 7157
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12952 7160 13277 7188
rect 12952 7148 12958 7160
rect 13265 7157 13277 7160
rect 13311 7188 13323 7191
rect 13630 7188 13636 7200
rect 13311 7160 13636 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 16540 7160 16681 7188
rect 16540 7148 16546 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 27522 7188 27528 7200
rect 27483 7160 27528 7188
rect 16669 7151 16727 7157
rect 27522 7148 27528 7160
rect 27580 7148 27586 7200
rect 29825 7191 29883 7197
rect 29825 7157 29837 7191
rect 29871 7188 29883 7191
rect 30098 7188 30104 7200
rect 29871 7160 30104 7188
rect 29871 7157 29883 7160
rect 29825 7151 29883 7157
rect 30098 7148 30104 7160
rect 30156 7148 30162 7200
rect 31110 7148 31116 7200
rect 31168 7188 31174 7200
rect 31205 7191 31263 7197
rect 31205 7188 31217 7191
rect 31168 7160 31217 7188
rect 31168 7148 31174 7160
rect 31205 7157 31217 7160
rect 31251 7157 31263 7191
rect 31205 7151 31263 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 4890 6984 4896 6996
rect 3936 6956 4896 6984
rect 3936 6944 3942 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 11756 6956 12265 6984
rect 11756 6944 11762 6956
rect 12253 6953 12265 6956
rect 12299 6953 12311 6987
rect 12253 6947 12311 6953
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 15933 6987 15991 6993
rect 15933 6984 15945 6987
rect 15896 6956 15945 6984
rect 15896 6944 15902 6956
rect 15933 6953 15945 6956
rect 15979 6953 15991 6987
rect 15933 6947 15991 6953
rect 16850 6944 16856 6996
rect 16908 6984 16914 6996
rect 17037 6987 17095 6993
rect 17037 6984 17049 6987
rect 16908 6956 17049 6984
rect 16908 6944 16914 6956
rect 17037 6953 17049 6956
rect 17083 6953 17095 6987
rect 17037 6947 17095 6953
rect 30834 6944 30840 6996
rect 30892 6984 30898 6996
rect 32766 6984 32772 6996
rect 30892 6956 32772 6984
rect 30892 6944 30898 6956
rect 32766 6944 32772 6956
rect 32824 6944 32830 6996
rect 36630 6984 36636 6996
rect 36591 6956 36636 6984
rect 36630 6944 36636 6956
rect 36688 6944 36694 6996
rect 38010 6984 38016 6996
rect 37971 6956 38016 6984
rect 38010 6944 38016 6956
rect 38068 6944 38074 6996
rect 27522 6916 27528 6928
rect 12084 6888 27528 6916
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 4028 6820 6285 6848
rect 4028 6808 4034 6820
rect 6273 6817 6285 6820
rect 6319 6817 6331 6851
rect 7006 6848 7012 6860
rect 6967 6820 7012 6848
rect 6273 6811 6331 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 11422 6808 11428 6860
rect 11480 6848 11486 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11480 6820 11621 6848
rect 11480 6808 11486 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11974 6848 11980 6860
rect 11609 6811 11667 6817
rect 11900 6820 11980 6848
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 7282 6789 7288 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 2096 6752 2145 6780
rect 2096 6740 2102 6752
rect 2133 6749 2145 6752
rect 2179 6780 2191 6783
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 2179 6752 5181 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 7276 6780 7288 6789
rect 7243 6752 7288 6780
rect 5169 6743 5227 6749
rect 7276 6743 7288 6752
rect 7282 6740 7288 6743
rect 7340 6740 7346 6792
rect 11900 6789 11928 6820
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12084 6789 12112 6888
rect 27522 6876 27528 6888
rect 27580 6876 27586 6928
rect 30098 6916 30104 6928
rect 30059 6888 30104 6916
rect 30098 6876 30104 6888
rect 30156 6876 30162 6928
rect 12802 6848 12808 6860
rect 12176 6820 12808 6848
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 4617 6715 4675 6721
rect 4617 6712 4629 6715
rect 2924 6684 4629 6712
rect 2924 6672 2930 6684
rect 4617 6681 4629 6684
rect 4663 6681 4675 6715
rect 4617 6675 4675 6681
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 5592 6684 8708 6712
rect 5592 6672 5598 6684
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2464 6616 2789 6644
rect 2464 6604 2470 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 2777 6607 2835 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5721 6647 5779 6653
rect 5721 6644 5733 6647
rect 4764 6616 5733 6644
rect 4764 6604 4770 6616
rect 5721 6613 5733 6616
rect 5767 6613 5779 6647
rect 5721 6607 5779 6613
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8570 6644 8576 6656
rect 8435 6616 8576 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8680 6644 8708 6684
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 11747 6715 11805 6721
rect 11747 6712 11759 6715
rect 11296 6684 11759 6712
rect 11296 6672 11302 6684
rect 11747 6681 11759 6684
rect 11793 6681 11805 6715
rect 11747 6675 11805 6681
rect 11977 6715 12035 6721
rect 11977 6681 11989 6715
rect 12023 6712 12035 6715
rect 12176 6712 12204 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 19242 6848 19248 6860
rect 16132 6820 19248 6848
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 16132 6789 16160 6820
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 12584 6752 16129 6780
rect 12584 6740 12590 6752
rect 16117 6749 16129 6752
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16356 6752 16405 6780
rect 16356 6740 16362 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16494 6783 16552 6789
rect 16494 6749 16506 6783
rect 16540 6749 16552 6783
rect 16494 6743 16552 6749
rect 17144 6774 17172 6820
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 23290 6848 23296 6860
rect 22066 6820 23296 6848
rect 17214 6777 17272 6783
rect 17494 6780 17500 6792
rect 17214 6774 17226 6777
rect 17144 6746 17226 6774
rect 17214 6743 17226 6746
rect 17260 6743 17272 6777
rect 17455 6752 17500 6780
rect 12023 6684 12204 6712
rect 12023 6681 12035 6684
rect 11977 6675 12035 6681
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 16500 6712 16528 6743
rect 17214 6737 17272 6743
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17598 6783 17656 6789
rect 17598 6749 17610 6783
rect 17644 6749 17656 6783
rect 17598 6743 17656 6749
rect 15804 6684 16528 6712
rect 15804 6672 15810 6684
rect 14458 6644 14464 6656
rect 8680 6616 14464 6644
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 17604 6644 17632 6743
rect 18414 6740 18420 6792
rect 18472 6780 18478 6792
rect 20441 6783 20499 6789
rect 20441 6780 20453 6783
rect 18472 6752 20453 6780
rect 18472 6740 18478 6752
rect 20441 6749 20453 6752
rect 20487 6780 20499 6783
rect 21818 6780 21824 6792
rect 20487 6752 21824 6780
rect 20487 6749 20499 6752
rect 20441 6743 20499 6749
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 17770 6672 17776 6724
rect 17828 6712 17834 6724
rect 22066 6712 22094 6820
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 24486 6848 24492 6860
rect 23584 6820 24492 6848
rect 23584 6789 23612 6820
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 25314 6808 25320 6860
rect 25372 6848 25378 6860
rect 26050 6848 26056 6860
rect 25372 6820 26056 6848
rect 25372 6808 25378 6820
rect 26050 6808 26056 6820
rect 26108 6808 26114 6860
rect 29086 6808 29092 6860
rect 29144 6848 29150 6860
rect 29825 6851 29883 6857
rect 29825 6848 29837 6851
rect 29144 6820 29837 6848
rect 29144 6808 29150 6820
rect 29825 6817 29837 6820
rect 29871 6848 29883 6851
rect 30006 6848 30012 6860
rect 29871 6820 30012 6848
rect 29871 6817 29883 6820
rect 29825 6811 29883 6817
rect 30006 6808 30012 6820
rect 30064 6808 30070 6860
rect 30285 6851 30343 6857
rect 30285 6817 30297 6851
rect 30331 6848 30343 6851
rect 30466 6848 30472 6860
rect 30331 6820 30472 6848
rect 30331 6817 30343 6820
rect 30285 6811 30343 6817
rect 30466 6808 30472 6820
rect 30524 6808 30530 6860
rect 30834 6848 30840 6860
rect 30795 6820 30840 6848
rect 30834 6808 30840 6820
rect 30892 6808 30898 6860
rect 31110 6789 31116 6792
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6749 23627 6783
rect 31104 6780 31116 6789
rect 31071 6752 31116 6780
rect 23569 6743 23627 6749
rect 31104 6743 31116 6752
rect 31110 6740 31116 6743
rect 31168 6740 31174 6792
rect 35989 6783 36047 6789
rect 35989 6749 36001 6783
rect 36035 6780 36047 6783
rect 36446 6780 36452 6792
rect 36035 6752 36452 6780
rect 36035 6749 36047 6752
rect 35989 6743 36047 6749
rect 36446 6740 36452 6752
rect 36504 6740 36510 6792
rect 37090 6780 37096 6792
rect 37051 6752 37096 6780
rect 37090 6740 37096 6752
rect 37148 6740 37154 6792
rect 37829 6783 37887 6789
rect 37829 6749 37841 6783
rect 37875 6749 37887 6783
rect 37829 6743 37887 6749
rect 17828 6684 22094 6712
rect 17828 6672 17834 6684
rect 30282 6672 30288 6724
rect 30340 6712 30346 6724
rect 37844 6712 37872 6743
rect 30340 6684 37872 6712
rect 30340 6672 30346 6684
rect 20622 6644 20628 6656
rect 16908 6616 17632 6644
rect 20583 6616 20628 6644
rect 16908 6604 16914 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 32232 6653 32260 6684
rect 32217 6647 32275 6653
rect 32217 6613 32229 6647
rect 32263 6613 32275 6647
rect 37274 6644 37280 6656
rect 37235 6616 37280 6644
rect 32217 6607 32275 6613
rect 37274 6604 37280 6616
rect 37332 6604 37338 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2133 6443 2191 6449
rect 2133 6409 2145 6443
rect 2179 6440 2191 6443
rect 6917 6443 6975 6449
rect 6917 6440 6929 6443
rect 2179 6412 6929 6440
rect 2179 6409 2191 6412
rect 2133 6403 2191 6409
rect 6917 6409 6929 6412
rect 6963 6440 6975 6443
rect 7558 6440 7564 6452
rect 6963 6412 7564 6440
rect 6963 6409 6975 6412
rect 6917 6403 6975 6409
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7708 6412 7941 6440
rect 7708 6400 7714 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 12216 6412 13185 6440
rect 12216 6400 12222 6412
rect 13173 6409 13185 6412
rect 13219 6440 13231 6443
rect 36814 6440 36820 6452
rect 13219 6412 36820 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 36814 6400 36820 6412
rect 36872 6400 36878 6452
rect 1854 6372 1860 6384
rect 1767 6344 1860 6372
rect 1854 6332 1860 6344
rect 1912 6372 1918 6384
rect 5718 6372 5724 6384
rect 1912 6344 5724 6372
rect 1912 6332 1918 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 7156 6344 15608 6372
rect 7156 6332 7162 6344
rect 2866 6304 2872 6316
rect 2827 6276 2872 6304
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4798 6304 4804 6316
rect 4212 6276 4804 6304
rect 4212 6264 4218 6276
rect 4798 6264 4804 6276
rect 4856 6304 4862 6316
rect 7116 6304 7144 6332
rect 8110 6304 8116 6316
rect 4856 6276 7144 6304
rect 8071 6276 8116 6304
rect 4856 6264 4862 6276
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8386 6304 8392 6316
rect 8347 6276 8392 6304
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9582 6304 9588 6316
rect 8628 6276 9588 6304
rect 8628 6264 8634 6276
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 12710 6304 12716 6316
rect 10836 6276 12716 6304
rect 10836 6264 10842 6276
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 15580 6304 15608 6344
rect 15654 6332 15660 6384
rect 15712 6372 15718 6384
rect 15850 6375 15908 6381
rect 15850 6372 15862 6375
rect 15712 6344 15862 6372
rect 15712 6332 15718 6344
rect 15850 6341 15862 6344
rect 15896 6341 15908 6375
rect 15850 6335 15908 6341
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 19613 6375 19671 6381
rect 19613 6372 19625 6375
rect 19392 6344 19625 6372
rect 19392 6332 19398 6344
rect 19613 6341 19625 6344
rect 19659 6372 19671 6375
rect 20257 6375 20315 6381
rect 20257 6372 20269 6375
rect 19659 6344 20269 6372
rect 19659 6341 19671 6344
rect 19613 6335 19671 6341
rect 20257 6341 20269 6344
rect 20303 6372 20315 6375
rect 20530 6372 20536 6384
rect 20303 6344 20536 6372
rect 20303 6341 20315 6344
rect 20257 6335 20315 6341
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 23106 6372 23112 6384
rect 23067 6344 23112 6372
rect 23106 6332 23112 6344
rect 23164 6332 23170 6384
rect 24578 6372 24584 6384
rect 23584 6344 24584 6372
rect 16117 6307 16175 6313
rect 15580 6276 16068 6304
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 11698 6236 11704 6248
rect 1728 6208 11704 6236
rect 1728 6196 1734 6208
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 16040 6236 16068 6276
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16574 6304 16580 6316
rect 16163 6276 16580 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16574 6264 16580 6276
rect 16632 6304 16638 6316
rect 17126 6304 17132 6316
rect 16632 6276 17132 6304
rect 16632 6264 16638 6276
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 21818 6304 21824 6316
rect 21779 6276 21824 6304
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 22097 6239 22155 6245
rect 16040 6208 16160 6236
rect 3694 6128 3700 6180
rect 3752 6168 3758 6180
rect 4709 6171 4767 6177
rect 4709 6168 4721 6171
rect 3752 6140 4721 6168
rect 3752 6128 3758 6140
rect 4709 6137 4721 6140
rect 4755 6137 4767 6171
rect 4709 6131 4767 6137
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 15102 6168 15108 6180
rect 11204 6140 15108 6168
rect 11204 6128 11210 6140
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 16132 6168 16160 6208
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 22462 6236 22468 6248
rect 22143 6208 22468 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 22462 6196 22468 6208
rect 22520 6236 22526 6248
rect 23308 6236 23336 6267
rect 23382 6264 23388 6316
rect 23440 6304 23446 6316
rect 23584 6313 23612 6344
rect 24578 6332 24584 6344
rect 24636 6332 24642 6384
rect 23569 6307 23627 6313
rect 23440 6276 23533 6304
rect 23440 6264 23446 6276
rect 23569 6273 23581 6307
rect 23615 6273 23627 6307
rect 23569 6267 23627 6273
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 23716 6276 23761 6304
rect 23716 6264 23722 6276
rect 34790 6264 34796 6316
rect 34848 6304 34854 6316
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 34848 6276 37841 6304
rect 34848 6264 34854 6276
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 22520 6208 23336 6236
rect 23400 6236 23428 6264
rect 34698 6236 34704 6248
rect 23400 6208 34704 6236
rect 22520 6196 22526 6208
rect 34698 6196 34704 6208
rect 34756 6196 34762 6248
rect 28994 6168 29000 6180
rect 16132 6140 29000 6168
rect 28994 6128 29000 6140
rect 29052 6168 29058 6180
rect 34514 6168 34520 6180
rect 29052 6140 34520 6168
rect 29052 6128 29058 6140
rect 34514 6128 34520 6140
rect 34572 6128 34578 6180
rect 35897 6171 35955 6177
rect 35897 6137 35909 6171
rect 35943 6168 35955 6171
rect 37182 6168 37188 6180
rect 35943 6140 37188 6168
rect 35943 6137 35955 6140
rect 35897 6131 35955 6137
rect 37182 6128 37188 6140
rect 37240 6128 37246 6180
rect 37369 6171 37427 6177
rect 37369 6137 37381 6171
rect 37415 6168 37427 6171
rect 38102 6168 38108 6180
rect 37415 6140 38108 6168
rect 37415 6137 37427 6140
rect 37369 6131 37427 6137
rect 38102 6128 38108 6140
rect 38160 6128 38166 6180
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3292 6072 3617 6100
rect 3292 6060 3298 6072
rect 3605 6069 3617 6072
rect 3651 6100 3663 6103
rect 4062 6100 4068 6112
rect 3651 6072 4068 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4614 6100 4620 6112
rect 4295 6072 4620 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 4856 6072 5273 6100
rect 4856 6060 4862 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8110 6100 8116 6112
rect 7616 6072 8116 6100
rect 7616 6060 7622 6072
rect 8110 6060 8116 6072
rect 8168 6100 8174 6112
rect 12526 6100 12532 6112
rect 8168 6072 12532 6100
rect 8168 6060 8174 6072
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 12621 6103 12679 6109
rect 12621 6069 12633 6103
rect 12667 6100 12679 6103
rect 12710 6100 12716 6112
rect 12667 6072 12716 6100
rect 12667 6069 12679 6072
rect 12621 6063 12679 6069
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 13412 6072 13645 6100
rect 13412 6060 13418 6072
rect 13633 6069 13645 6072
rect 13679 6069 13691 6103
rect 13633 6063 13691 6069
rect 14737 6103 14795 6109
rect 14737 6069 14749 6103
rect 14783 6100 14795 6103
rect 15746 6100 15752 6112
rect 14783 6072 15752 6100
rect 14783 6069 14795 6072
rect 14737 6063 14795 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 20346 6100 20352 6112
rect 20307 6072 20352 6100
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 24213 6103 24271 6109
rect 24213 6100 24225 6103
rect 22612 6072 24225 6100
rect 22612 6060 22618 6072
rect 24213 6069 24225 6072
rect 24259 6100 24271 6103
rect 25958 6100 25964 6112
rect 24259 6072 25964 6100
rect 24259 6069 24271 6072
rect 24213 6063 24271 6069
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 26050 6060 26056 6112
rect 26108 6100 26114 6112
rect 35345 6103 35403 6109
rect 35345 6100 35357 6103
rect 26108 6072 35357 6100
rect 26108 6060 26114 6072
rect 35345 6069 35357 6072
rect 35391 6100 35403 6103
rect 35618 6100 35624 6112
rect 35391 6072 35624 6100
rect 35391 6069 35403 6072
rect 35345 6063 35403 6069
rect 35618 6060 35624 6072
rect 35676 6060 35682 6112
rect 35710 6060 35716 6112
rect 35768 6100 35774 6112
rect 36357 6103 36415 6109
rect 36357 6100 36369 6103
rect 35768 6072 36369 6100
rect 35768 6060 35774 6072
rect 36357 6069 36369 6072
rect 36403 6069 36415 6103
rect 38010 6100 38016 6112
rect 37971 6072 38016 6100
rect 36357 6063 36415 6069
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 7098 5896 7104 5908
rect 6319 5868 7104 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7374 5896 7380 5908
rect 7287 5868 7380 5896
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 7834 5896 7840 5908
rect 7432 5868 7840 5896
rect 7432 5856 7438 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 11333 5899 11391 5905
rect 11333 5865 11345 5899
rect 11379 5896 11391 5899
rect 12434 5896 12440 5908
rect 11379 5868 12440 5896
rect 11379 5865 11391 5868
rect 11333 5859 11391 5865
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14231 5868 16620 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 2556 5800 3801 5828
rect 2556 5788 2562 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 6362 5828 6368 5840
rect 4571 5800 6368 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 4540 5760 4568 5791
rect 6362 5788 6368 5800
rect 6420 5788 6426 5840
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 13173 5831 13231 5837
rect 13173 5828 13185 5831
rect 13044 5800 13185 5828
rect 13044 5788 13050 5800
rect 13173 5797 13185 5800
rect 13219 5797 13231 5831
rect 13173 5791 13231 5797
rect 7466 5760 7472 5772
rect 3476 5732 4568 5760
rect 7427 5732 7472 5760
rect 3476 5720 3482 5732
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 11793 5763 11851 5769
rect 9640 5732 11100 5760
rect 9640 5720 9646 5732
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3160 5624 3188 5655
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3970 5692 3976 5704
rect 3384 5664 3976 5692
rect 3384 5652 3390 5664
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10778 5692 10784 5704
rect 10376 5664 10784 5692
rect 10376 5652 10382 5664
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11072 5701 11100 5732
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 11882 5760 11888 5772
rect 11839 5732 11888 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 14200 5704 14228 5859
rect 16592 5828 16620 5868
rect 18322 5856 18328 5908
rect 18380 5896 18386 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 18380 5868 19809 5896
rect 18380 5856 18386 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 19797 5859 19855 5865
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 21637 5899 21695 5905
rect 21637 5896 21649 5899
rect 20588 5868 21649 5896
rect 20588 5856 20594 5868
rect 21637 5865 21649 5868
rect 21683 5865 21695 5899
rect 21637 5859 21695 5865
rect 22186 5856 22192 5908
rect 22244 5896 22250 5908
rect 22281 5899 22339 5905
rect 22281 5896 22293 5899
rect 22244 5868 22293 5896
rect 22244 5856 22250 5868
rect 22281 5865 22293 5868
rect 22327 5865 22339 5899
rect 22281 5859 22339 5865
rect 23198 5856 23204 5908
rect 23256 5896 23262 5908
rect 23293 5899 23351 5905
rect 23293 5896 23305 5899
rect 23256 5868 23305 5896
rect 23256 5856 23262 5868
rect 23293 5865 23305 5868
rect 23339 5865 23351 5899
rect 23658 5896 23664 5908
rect 23293 5859 23351 5865
rect 23492 5868 23664 5896
rect 20622 5828 20628 5840
rect 16592 5800 20628 5828
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 16574 5760 16580 5772
rect 16535 5732 16580 5760
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 23492 5760 23520 5868
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 24118 5856 24124 5908
rect 24176 5896 24182 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 24176 5868 24409 5896
rect 24176 5856 24182 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 24397 5859 24455 5865
rect 25777 5899 25835 5905
rect 25777 5865 25789 5899
rect 25823 5896 25835 5899
rect 25866 5896 25872 5908
rect 25823 5868 25872 5896
rect 25823 5865 25835 5868
rect 25777 5859 25835 5865
rect 25866 5856 25872 5868
rect 25924 5856 25930 5908
rect 28905 5899 28963 5905
rect 28905 5865 28917 5899
rect 28951 5896 28963 5899
rect 28994 5896 29000 5908
rect 28951 5868 29000 5896
rect 28951 5865 28963 5868
rect 28905 5859 28963 5865
rect 28994 5856 29000 5868
rect 29052 5856 29058 5908
rect 33410 5896 33416 5908
rect 33371 5868 33416 5896
rect 33410 5856 33416 5868
rect 33468 5856 33474 5908
rect 36814 5896 36820 5908
rect 36775 5868 36820 5896
rect 36814 5856 36820 5868
rect 36872 5856 36878 5908
rect 23566 5788 23572 5840
rect 23624 5828 23630 5840
rect 25130 5828 25136 5840
rect 23624 5800 25136 5828
rect 23624 5788 23630 5800
rect 25130 5788 25136 5800
rect 25188 5788 25194 5840
rect 22066 5732 24992 5760
rect 11057 5695 11115 5701
rect 10928 5664 10973 5692
rect 10928 5652 10934 5664
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 12066 5692 12072 5704
rect 11204 5664 11249 5692
rect 12027 5664 12072 5692
rect 11204 5652 11210 5664
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12250 5692 12256 5704
rect 12211 5664 12256 5692
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5692 13415 5695
rect 14182 5692 14188 5704
rect 13403 5664 14188 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 16321 5695 16379 5701
rect 16321 5661 16333 5695
rect 16367 5692 16379 5695
rect 16482 5692 16488 5704
rect 16367 5664 16488 5692
rect 16367 5661 16379 5664
rect 16321 5655 16379 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18288 5664 19257 5692
rect 18288 5652 18294 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19521 5695 19579 5701
rect 19392 5664 19437 5692
rect 19392 5652 19398 5664
rect 19521 5661 19533 5695
rect 19567 5661 19579 5695
rect 19521 5655 19579 5661
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19978 5692 19984 5704
rect 19659 5664 19984 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 3160 5596 11468 5624
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 2774 5556 2780 5568
rect 2271 5528 2780 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 7098 5556 7104 5568
rect 7055 5528 7104 5556
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 11440 5556 11468 5596
rect 11514 5584 11520 5636
rect 11572 5624 11578 5636
rect 11931 5627 11989 5633
rect 11931 5624 11943 5627
rect 11572 5596 11943 5624
rect 11572 5584 11578 5596
rect 11931 5593 11943 5596
rect 11977 5593 11989 5627
rect 11931 5587 11989 5593
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 19536 5624 19564 5655
rect 19978 5652 19984 5664
rect 20036 5652 20042 5704
rect 20070 5624 20076 5636
rect 12216 5596 12261 5624
rect 19536 5596 20076 5624
rect 12216 5584 12222 5596
rect 20070 5584 20076 5596
rect 20128 5584 20134 5636
rect 12437 5559 12495 5565
rect 12437 5556 12449 5559
rect 11440 5528 12449 5556
rect 12437 5525 12449 5528
rect 12483 5525 12495 5559
rect 15194 5556 15200 5568
rect 15155 5528 15200 5556
rect 12437 5519 12495 5525
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 20622 5556 20628 5568
rect 20404 5528 20628 5556
rect 20404 5516 20410 5528
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 21726 5516 21732 5568
rect 21784 5556 21790 5568
rect 22066 5556 22094 5732
rect 22462 5692 22468 5704
rect 22423 5664 22468 5692
rect 22462 5652 22468 5664
rect 22520 5652 22526 5704
rect 22554 5652 22560 5704
rect 22612 5692 22618 5704
rect 22738 5692 22744 5704
rect 22612 5664 22657 5692
rect 22699 5664 22744 5692
rect 22612 5652 22618 5664
rect 22738 5652 22744 5664
rect 22796 5652 22802 5704
rect 22848 5701 22876 5732
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 23477 5695 23535 5701
rect 23477 5661 23489 5695
rect 23523 5661 23535 5695
rect 23477 5655 23535 5661
rect 22480 5624 22508 5652
rect 23492 5624 23520 5655
rect 23566 5652 23572 5704
rect 23624 5692 23630 5704
rect 23750 5692 23756 5704
rect 23624 5664 23669 5692
rect 23711 5664 23756 5692
rect 23624 5652 23630 5664
rect 23750 5652 23756 5664
rect 23808 5652 23814 5704
rect 23860 5701 23888 5732
rect 23845 5695 23903 5701
rect 23845 5661 23857 5695
rect 23891 5661 23903 5695
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23845 5655 23903 5661
rect 24136 5664 24593 5692
rect 24136 5636 24164 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5661 24731 5695
rect 24854 5692 24860 5704
rect 24815 5664 24860 5692
rect 24673 5655 24731 5661
rect 24118 5624 24124 5636
rect 22480 5596 24124 5624
rect 24118 5584 24124 5596
rect 24176 5584 24182 5636
rect 24688 5624 24716 5655
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 24964 5701 24992 5732
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 25148 5692 25176 5788
rect 25884 5760 25912 5856
rect 25958 5788 25964 5840
rect 26016 5828 26022 5840
rect 32858 5828 32864 5840
rect 26016 5800 32864 5828
rect 26016 5788 26022 5800
rect 32858 5788 32864 5800
rect 32916 5788 32922 5840
rect 36265 5831 36323 5837
rect 36265 5797 36277 5831
rect 36311 5828 36323 5831
rect 36311 5800 37320 5828
rect 36311 5797 36323 5800
rect 36265 5791 36323 5797
rect 26237 5763 26295 5769
rect 26237 5760 26249 5763
rect 25884 5732 26249 5760
rect 26237 5729 26249 5732
rect 26283 5760 26295 5763
rect 26418 5760 26424 5772
rect 26283 5732 26424 5760
rect 26283 5729 26295 5732
rect 26237 5723 26295 5729
rect 26418 5720 26424 5732
rect 26476 5720 26482 5772
rect 26513 5763 26571 5769
rect 26513 5729 26525 5763
rect 26559 5760 26571 5763
rect 27706 5760 27712 5772
rect 26559 5732 27712 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 27706 5720 27712 5732
rect 27764 5720 27770 5772
rect 34606 5720 34612 5772
rect 34664 5760 34670 5772
rect 34793 5763 34851 5769
rect 34793 5760 34805 5763
rect 34664 5732 34805 5760
rect 34664 5720 34670 5732
rect 34793 5729 34805 5732
rect 34839 5729 34851 5763
rect 34793 5723 34851 5729
rect 26050 5692 26056 5704
rect 25148 5664 26056 5692
rect 24949 5655 25007 5661
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 34514 5652 34520 5704
rect 34572 5692 34578 5704
rect 35069 5695 35127 5701
rect 35069 5692 35081 5695
rect 34572 5664 35081 5692
rect 34572 5652 34578 5664
rect 35069 5661 35081 5664
rect 35115 5661 35127 5695
rect 35069 5655 35127 5661
rect 35710 5652 35716 5704
rect 35768 5692 35774 5704
rect 37090 5701 37096 5704
rect 36081 5695 36139 5701
rect 36081 5692 36093 5695
rect 35768 5664 36093 5692
rect 35768 5652 35774 5664
rect 36081 5661 36093 5664
rect 36127 5661 36139 5695
rect 36081 5655 36139 5661
rect 36996 5695 37054 5701
rect 36996 5661 37008 5695
rect 37042 5661 37054 5695
rect 36996 5655 37054 5661
rect 37084 5655 37096 5701
rect 37148 5692 37154 5704
rect 37292 5701 37320 5800
rect 37292 5695 37371 5701
rect 37148 5664 37184 5692
rect 37292 5664 37325 5695
rect 27522 5624 27528 5636
rect 24688 5596 27528 5624
rect 27522 5584 27528 5596
rect 27580 5584 27586 5636
rect 34977 5627 35035 5633
rect 34977 5593 34989 5627
rect 35023 5624 35035 5627
rect 36906 5624 36912 5636
rect 35023 5596 36912 5624
rect 35023 5593 35035 5596
rect 34977 5587 35035 5593
rect 36906 5584 36912 5596
rect 36964 5584 36970 5636
rect 21784 5528 22094 5556
rect 34149 5559 34207 5565
rect 21784 5516 21790 5528
rect 34149 5525 34161 5559
rect 34195 5556 34207 5559
rect 34422 5556 34428 5568
rect 34195 5528 34428 5556
rect 34195 5525 34207 5528
rect 34149 5519 34207 5525
rect 34422 5516 34428 5528
rect 34480 5516 34486 5568
rect 35434 5556 35440 5568
rect 35395 5528 35440 5556
rect 35434 5516 35440 5528
rect 35492 5516 35498 5568
rect 37016 5556 37044 5655
rect 37090 5652 37096 5655
rect 37148 5652 37154 5664
rect 37313 5661 37325 5664
rect 37359 5661 37371 5695
rect 37313 5655 37371 5661
rect 37461 5695 37519 5701
rect 37461 5661 37473 5695
rect 37507 5692 37519 5695
rect 37918 5692 37924 5704
rect 37507 5664 37924 5692
rect 37507 5661 37519 5664
rect 37461 5655 37519 5661
rect 37918 5652 37924 5664
rect 37976 5652 37982 5704
rect 38102 5692 38108 5704
rect 38063 5664 38108 5692
rect 38102 5652 38108 5664
rect 38160 5652 38166 5704
rect 37185 5627 37243 5633
rect 37185 5593 37197 5627
rect 37231 5624 37243 5627
rect 37734 5624 37740 5636
rect 37231 5596 37740 5624
rect 37231 5593 37243 5596
rect 37185 5587 37243 5593
rect 37734 5584 37740 5596
rect 37792 5584 37798 5636
rect 37550 5556 37556 5568
rect 37016 5528 37556 5556
rect 37550 5516 37556 5528
rect 37608 5516 37614 5568
rect 37918 5556 37924 5568
rect 37879 5528 37924 5556
rect 37918 5516 37924 5528
rect 37976 5516 37982 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3786 5352 3792 5364
rect 3747 5324 3792 5352
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7248 5324 7389 5352
rect 7248 5312 7254 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 11238 5352 11244 5364
rect 10919 5324 11244 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 12710 5352 12716 5364
rect 12406 5324 12716 5352
rect 2406 5244 2412 5296
rect 2464 5284 2470 5296
rect 6914 5284 6920 5296
rect 2464 5256 6592 5284
rect 2464 5244 2470 5256
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2682 5216 2688 5228
rect 2363 5188 2688 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 3418 5216 3424 5228
rect 3379 5188 3424 5216
rect 2869 5179 2927 5185
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 2884 5148 2912 5179
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 5166 5216 5172 5228
rect 5127 5188 5172 5216
rect 4893 5179 4951 5185
rect 2648 5120 2912 5148
rect 4908 5148 4936 5179
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 5534 5216 5540 5228
rect 5399 5188 5540 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 5626 5148 5632 5160
rect 4908 5120 5632 5148
rect 2648 5108 2654 5120
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 3050 5080 3056 5092
rect 1811 5052 3056 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 3050 5040 3056 5052
rect 3108 5040 3114 5092
rect 6564 5080 6592 5256
rect 6656 5256 6920 5284
rect 6656 5225 6684 5256
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 8110 5284 8116 5296
rect 8023 5256 8116 5284
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7190 5216 7196 5228
rect 6871 5188 7196 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7190 5176 7196 5188
rect 7248 5216 7254 5228
rect 7374 5216 7380 5228
rect 7248 5188 7380 5216
rect 7248 5176 7254 5188
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7558 5216 7564 5228
rect 7519 5188 7564 5216
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 8036 5225 8064 5256
rect 8110 5244 8116 5256
rect 8168 5284 8174 5296
rect 12066 5284 12072 5296
rect 8168 5256 10640 5284
rect 12027 5256 12072 5284
rect 8168 5244 8174 5256
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 10318 5216 10324 5228
rect 10279 5188 10324 5216
rect 8021 5179 8079 5185
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 7282 5148 7288 5160
rect 6963 5120 7288 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7852 5148 7880 5179
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 10410 5176 10416 5228
rect 10468 5216 10474 5228
rect 10612 5225 10640 5256
rect 12066 5244 12072 5256
rect 12124 5244 12130 5296
rect 12161 5287 12219 5293
rect 12161 5253 12173 5287
rect 12207 5284 12219 5287
rect 12406 5284 12434 5324
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 12894 5352 12900 5364
rect 12855 5324 12900 5352
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13998 5352 14004 5364
rect 13959 5324 14004 5352
rect 13998 5312 14004 5324
rect 14056 5352 14062 5364
rect 14458 5352 14464 5364
rect 14056 5324 14464 5352
rect 14056 5312 14062 5324
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 20533 5355 20591 5361
rect 20533 5352 20545 5355
rect 19484 5324 20545 5352
rect 19484 5312 19490 5324
rect 20533 5321 20545 5324
rect 20579 5321 20591 5355
rect 20533 5315 20591 5321
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 23382 5352 23388 5364
rect 20680 5324 23388 5352
rect 20680 5312 20686 5324
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 23934 5352 23940 5364
rect 23895 5324 23940 5352
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 26142 5312 26148 5364
rect 26200 5352 26206 5364
rect 27249 5355 27307 5361
rect 27249 5352 27261 5355
rect 26200 5324 27261 5352
rect 26200 5312 26206 5324
rect 27249 5321 27261 5324
rect 27295 5321 27307 5355
rect 27249 5315 27307 5321
rect 28537 5355 28595 5361
rect 28537 5321 28549 5355
rect 28583 5321 28595 5355
rect 28537 5315 28595 5321
rect 13262 5284 13268 5296
rect 12207 5256 12434 5284
rect 13223 5256 13268 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 13262 5244 13268 5256
rect 13320 5244 13326 5296
rect 13403 5287 13461 5293
rect 13403 5253 13415 5287
rect 13449 5284 13461 5287
rect 13538 5284 13544 5296
rect 13449 5256 13544 5284
rect 13449 5253 13461 5256
rect 13403 5247 13461 5253
rect 13538 5244 13544 5256
rect 13596 5244 13602 5296
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 14792 5256 15117 5284
rect 14792 5244 14798 5256
rect 15105 5253 15117 5256
rect 15151 5253 15163 5287
rect 15286 5284 15292 5296
rect 15199 5256 15292 5284
rect 15105 5247 15163 5253
rect 10597 5219 10655 5225
rect 10468 5188 10513 5216
rect 10468 5176 10474 5188
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 8386 5148 8392 5160
rect 7524 5120 8392 5148
rect 7524 5108 7530 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 10704 5080 10732 5179
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11931 5219 11989 5225
rect 11931 5216 11943 5219
rect 11112 5188 11943 5216
rect 11112 5176 11118 5188
rect 11931 5185 11943 5188
rect 11977 5185 11989 5219
rect 11931 5179 11989 5185
rect 11790 5148 11796 5160
rect 11751 5120 11796 5148
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 12084 5148 12112 5244
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 13081 5219 13139 5225
rect 12308 5188 12353 5216
rect 12308 5176 12314 5188
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 13096 5148 13124 5179
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 13228 5188 13273 5216
rect 13228 5176 13234 5188
rect 13538 5148 13544 5160
rect 12084 5120 13124 5148
rect 13499 5120 13544 5148
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 15120 5148 15148 5247
rect 15286 5244 15292 5256
rect 15344 5284 15350 5296
rect 21726 5284 21732 5296
rect 15344 5256 21732 5284
rect 15344 5244 15350 5256
rect 21726 5244 21732 5256
rect 21784 5244 21790 5296
rect 24302 5284 24308 5296
rect 22066 5256 24308 5284
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17310 5216 17316 5228
rect 17175 5188 17316 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17310 5176 17316 5188
rect 17368 5216 17374 5228
rect 18230 5216 18236 5228
rect 17368 5188 18092 5216
rect 18191 5188 18236 5216
rect 17368 5176 17374 5188
rect 17954 5148 17960 5160
rect 15120 5120 17960 5148
rect 17954 5108 17960 5120
rect 18012 5108 18018 5160
rect 18064 5148 18092 5188
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 19058 5216 19064 5228
rect 18656 5188 19064 5216
rect 18656 5176 18662 5188
rect 19058 5176 19064 5188
rect 19116 5176 19122 5228
rect 19521 5219 19579 5225
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 19978 5216 19984 5228
rect 19567 5188 19984 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 19978 5176 19984 5188
rect 20036 5216 20042 5228
rect 20622 5216 20628 5228
rect 20036 5188 20628 5216
rect 20036 5176 20042 5188
rect 20622 5176 20628 5188
rect 20680 5216 20686 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 20680 5188 20729 5216
rect 20680 5176 20686 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 20990 5216 20996 5228
rect 20864 5188 20909 5216
rect 20951 5188 20996 5216
rect 20864 5176 20870 5188
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 21082 5176 21088 5228
rect 21140 5216 21146 5228
rect 22066 5216 22094 5256
rect 24302 5244 24308 5256
rect 24360 5284 24366 5296
rect 27617 5287 27675 5293
rect 24360 5256 24532 5284
rect 24360 5244 24366 5256
rect 24118 5216 24124 5228
rect 21140 5188 22094 5216
rect 24079 5188 24124 5216
rect 21140 5176 21146 5188
rect 24118 5176 24124 5188
rect 24176 5176 24182 5228
rect 24213 5219 24271 5225
rect 24213 5185 24225 5219
rect 24259 5185 24271 5219
rect 24394 5216 24400 5228
rect 24355 5188 24400 5216
rect 24213 5179 24271 5185
rect 19245 5151 19303 5157
rect 19245 5148 19257 5151
rect 18064 5120 19257 5148
rect 19245 5117 19257 5120
rect 19291 5117 19303 5151
rect 19245 5111 19303 5117
rect 20530 5108 20536 5160
rect 20588 5148 20594 5160
rect 21821 5151 21879 5157
rect 21821 5148 21833 5151
rect 20588 5120 21833 5148
rect 20588 5108 20594 5120
rect 21821 5117 21833 5120
rect 21867 5117 21879 5151
rect 21821 5111 21879 5117
rect 22097 5151 22155 5157
rect 22097 5117 22109 5151
rect 22143 5148 22155 5151
rect 22370 5148 22376 5160
rect 22143 5120 22376 5148
rect 22143 5117 22155 5120
rect 22097 5111 22155 5117
rect 22370 5108 22376 5120
rect 22428 5108 22434 5160
rect 23934 5108 23940 5160
rect 23992 5148 23998 5160
rect 24228 5148 24256 5179
rect 24394 5176 24400 5188
rect 24452 5176 24458 5228
rect 24504 5225 24532 5256
rect 27617 5253 27629 5287
rect 27663 5284 27675 5287
rect 27706 5284 27712 5296
rect 27663 5256 27712 5284
rect 27663 5253 27675 5256
rect 27617 5247 27675 5253
rect 27706 5244 27712 5256
rect 27764 5244 27770 5296
rect 28552 5284 28580 5315
rect 28994 5312 29000 5364
rect 29052 5352 29058 5364
rect 29365 5355 29423 5361
rect 29365 5352 29377 5355
rect 29052 5324 29377 5352
rect 29052 5312 29058 5324
rect 29365 5321 29377 5324
rect 29411 5321 29423 5355
rect 32214 5352 32220 5364
rect 32175 5324 32220 5352
rect 29365 5315 29423 5321
rect 32214 5312 32220 5324
rect 32272 5312 32278 5364
rect 32858 5352 32864 5364
rect 32819 5324 32864 5352
rect 32858 5312 32864 5324
rect 32916 5312 32922 5364
rect 34330 5312 34336 5364
rect 34388 5352 34394 5364
rect 34388 5324 35204 5352
rect 34388 5312 34394 5324
rect 35176 5293 35204 5324
rect 37826 5312 37832 5364
rect 37884 5352 37890 5364
rect 37884 5324 38056 5352
rect 37884 5312 37890 5324
rect 35161 5287 35219 5293
rect 28552 5256 30420 5284
rect 30392 5225 30420 5256
rect 35161 5253 35173 5287
rect 35207 5253 35219 5287
rect 37645 5287 37703 5293
rect 37645 5284 37657 5287
rect 35161 5247 35219 5253
rect 35544 5256 37657 5284
rect 35544 5228 35572 5256
rect 37645 5253 37657 5256
rect 37691 5253 37703 5287
rect 37645 5247 37703 5253
rect 37734 5244 37740 5296
rect 37792 5284 37798 5296
rect 37792 5256 37837 5284
rect 37792 5244 37798 5256
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5185 24547 5219
rect 24489 5179 24547 5185
rect 27433 5219 27491 5225
rect 27433 5185 27445 5219
rect 27479 5216 27491 5219
rect 30377 5219 30435 5225
rect 27479 5188 29316 5216
rect 27479 5185 27491 5188
rect 27433 5179 27491 5185
rect 24670 5148 24676 5160
rect 23992 5120 24676 5148
rect 23992 5108 23998 5120
rect 24670 5108 24676 5120
rect 24728 5108 24734 5160
rect 28077 5151 28135 5157
rect 28077 5117 28089 5151
rect 28123 5148 28135 5151
rect 29086 5148 29092 5160
rect 28123 5120 29092 5148
rect 28123 5117 28135 5120
rect 28077 5111 28135 5117
rect 29086 5108 29092 5120
rect 29144 5108 29150 5160
rect 29288 5148 29316 5188
rect 30377 5185 30389 5219
rect 30423 5185 30435 5219
rect 34333 5219 34391 5225
rect 34333 5216 34345 5219
rect 30377 5179 30435 5185
rect 33428 5188 34345 5216
rect 29454 5148 29460 5160
rect 29288 5120 29460 5148
rect 29454 5108 29460 5120
rect 29512 5108 29518 5160
rect 29641 5151 29699 5157
rect 29641 5117 29653 5151
rect 29687 5148 29699 5151
rect 30190 5148 30196 5160
rect 29687 5120 30196 5148
rect 29687 5117 29699 5120
rect 29641 5111 29699 5117
rect 10962 5080 10968 5092
rect 6564 5052 6960 5080
rect 10704 5052 10968 5080
rect 4709 5015 4767 5021
rect 4709 4981 4721 5015
rect 4755 5012 4767 5015
rect 5074 5012 5080 5024
rect 4755 4984 5080 5012
rect 4755 4981 4767 4984
rect 4709 4975 4767 4981
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6328 4984 6469 5012
rect 6328 4972 6334 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6932 5012 6960 5052
rect 10962 5040 10968 5052
rect 11020 5080 11026 5092
rect 12986 5080 12992 5092
rect 11020 5052 12992 5080
rect 11020 5040 11026 5052
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 24210 5040 24216 5092
rect 24268 5080 24274 5092
rect 27798 5080 27804 5092
rect 24268 5052 27804 5080
rect 24268 5040 24274 5052
rect 27798 5040 27804 5052
rect 27856 5040 27862 5092
rect 28445 5083 28503 5089
rect 28445 5049 28457 5083
rect 28491 5080 28503 5083
rect 28997 5083 29055 5089
rect 28997 5080 29009 5083
rect 28491 5052 29009 5080
rect 28491 5049 28503 5052
rect 28445 5043 28503 5049
rect 28997 5049 29009 5052
rect 29043 5049 29055 5083
rect 28997 5043 29055 5049
rect 29178 5040 29184 5092
rect 29236 5080 29242 5092
rect 29656 5080 29684 5111
rect 30190 5108 30196 5120
rect 30248 5108 30254 5160
rect 33428 5089 33456 5188
rect 34333 5185 34345 5188
rect 34379 5185 34391 5219
rect 34333 5179 34391 5185
rect 34425 5219 34483 5225
rect 34425 5185 34437 5219
rect 34471 5216 34483 5219
rect 35526 5216 35532 5228
rect 34471 5188 35532 5216
rect 34471 5185 34483 5188
rect 34425 5179 34483 5185
rect 35526 5176 35532 5188
rect 35584 5176 35590 5228
rect 37550 5225 37556 5228
rect 36081 5219 36139 5225
rect 36081 5216 36093 5219
rect 35636 5188 36093 5216
rect 34606 5148 34612 5160
rect 34567 5120 34612 5148
rect 34606 5108 34612 5120
rect 34664 5108 34670 5160
rect 35636 5157 35664 5188
rect 36081 5185 36093 5188
rect 36127 5185 36139 5219
rect 37548 5216 37556 5225
rect 37511 5188 37556 5216
rect 36081 5179 36139 5185
rect 37548 5179 37556 5188
rect 37550 5176 37556 5179
rect 37608 5176 37614 5228
rect 37918 5216 37924 5228
rect 37879 5188 37924 5216
rect 37918 5176 37924 5188
rect 37976 5176 37982 5228
rect 38028 5225 38056 5324
rect 38013 5219 38071 5225
rect 38013 5185 38025 5219
rect 38059 5185 38071 5219
rect 38013 5179 38071 5185
rect 35621 5151 35679 5157
rect 35621 5117 35633 5151
rect 35667 5117 35679 5151
rect 35621 5111 35679 5117
rect 33413 5083 33471 5089
rect 33413 5080 33425 5083
rect 29236 5052 29684 5080
rect 29748 5052 33425 5080
rect 29236 5040 29242 5052
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 6932 4984 12449 5012
rect 6457 4975 6515 4981
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 17218 5012 17224 5024
rect 17179 4984 17224 5012
rect 12437 4975 12495 4981
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 23106 4972 23112 5024
rect 23164 5012 23170 5024
rect 23201 5015 23259 5021
rect 23201 5012 23213 5015
rect 23164 4984 23213 5012
rect 23164 4972 23170 4984
rect 23201 4981 23213 4984
rect 23247 5012 23259 5015
rect 25317 5015 25375 5021
rect 25317 5012 25329 5015
rect 23247 4984 25329 5012
rect 23247 4981 23259 4984
rect 23201 4975 23259 4981
rect 25317 4981 25329 4984
rect 25363 5012 25375 5015
rect 25682 5012 25688 5024
rect 25363 4984 25688 5012
rect 25363 4981 25375 4984
rect 25317 4975 25375 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 25774 4972 25780 5024
rect 25832 5012 25838 5024
rect 25832 4984 25877 5012
rect 25832 4972 25838 4984
rect 28626 4972 28632 5024
rect 28684 5012 28690 5024
rect 29748 5012 29776 5052
rect 33413 5049 33425 5052
rect 33459 5049 33471 5083
rect 35434 5080 35440 5092
rect 35395 5052 35440 5080
rect 33413 5043 33471 5049
rect 35434 5040 35440 5052
rect 35492 5040 35498 5092
rect 37366 5080 37372 5092
rect 37327 5052 37372 5080
rect 37366 5040 37372 5052
rect 37424 5040 37430 5092
rect 30190 5012 30196 5024
rect 28684 4984 29776 5012
rect 30151 4984 30196 5012
rect 28684 4972 28690 4984
rect 30190 4972 30196 4984
rect 30248 4972 30254 5024
rect 33594 4972 33600 5024
rect 33652 5012 33658 5024
rect 33965 5015 34023 5021
rect 33965 5012 33977 5015
rect 33652 4984 33977 5012
rect 33652 4972 33658 4984
rect 33965 4981 33977 4984
rect 34011 4981 34023 5015
rect 36262 5012 36268 5024
rect 36223 4984 36268 5012
rect 33965 4975 34023 4981
rect 36262 4972 36268 4984
rect 36320 4972 36326 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1946 4768 1952 4820
rect 2004 4808 2010 4820
rect 2590 4808 2596 4820
rect 2004 4780 2596 4808
rect 2004 4768 2010 4780
rect 2590 4768 2596 4780
rect 2648 4808 2654 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2648 4780 2789 4808
rect 2648 4768 2654 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3510 4808 3516 4820
rect 3099 4780 3516 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5684 4780 5825 4808
rect 5684 4768 5690 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 7006 4808 7012 4820
rect 5813 4771 5871 4777
rect 6748 4780 7012 4808
rect 2133 4743 2191 4749
rect 2133 4709 2145 4743
rect 2179 4740 2191 4743
rect 4890 4740 4896 4752
rect 2179 4712 4896 4740
rect 2179 4709 2191 4712
rect 2133 4703 2191 4709
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 4246 4672 4252 4684
rect 4207 4644 4252 4672
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 5644 4672 5672 4768
rect 4908 4644 5672 4672
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3234 4604 3240 4616
rect 2915 4576 3240 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3234 4564 3240 4576
rect 3292 4604 3298 4616
rect 3602 4604 3608 4616
rect 3292 4576 3608 4604
rect 3292 4564 3298 4576
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 4154 4604 4160 4616
rect 4115 4576 4160 4604
rect 3973 4567 4031 4573
rect 1854 4536 1860 4548
rect 1767 4508 1860 4536
rect 1854 4496 1860 4508
rect 1912 4536 1918 4548
rect 3878 4536 3884 4548
rect 1912 4508 3884 4536
rect 1912 4496 1918 4508
rect 3878 4496 3884 4508
rect 3936 4496 3942 4548
rect 3988 4536 4016 4567
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4908 4613 4936 4644
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6748 4681 6776 4780
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 8110 4808 8116 4820
rect 8071 4780 8116 4808
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 11054 4808 11060 4820
rect 11015 4780 11060 4808
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 13630 4768 13636 4820
rect 13688 4808 13694 4820
rect 15562 4808 15568 4820
rect 13688 4780 14412 4808
rect 15523 4780 15568 4808
rect 13688 4768 13694 4780
rect 13262 4700 13268 4752
rect 13320 4740 13326 4752
rect 14274 4740 14280 4752
rect 13320 4712 14280 4740
rect 13320 4700 13326 4712
rect 14274 4700 14280 4712
rect 14332 4700 14338 4752
rect 14384 4749 14412 4780
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 17034 4808 17040 4820
rect 16623 4780 17040 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 17586 4808 17592 4820
rect 17547 4780 17592 4808
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 18598 4808 18604 4820
rect 18559 4780 18604 4808
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 22557 4811 22615 4817
rect 22557 4777 22569 4811
rect 22603 4808 22615 4811
rect 22646 4808 22652 4820
rect 22603 4780 22652 4808
rect 22603 4777 22615 4780
rect 22557 4771 22615 4777
rect 22646 4768 22652 4780
rect 22704 4768 22710 4820
rect 23293 4811 23351 4817
rect 23293 4777 23305 4811
rect 23339 4808 23351 4811
rect 23750 4808 23756 4820
rect 23339 4780 23756 4808
rect 23339 4777 23351 4780
rect 23293 4771 23351 4777
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 24946 4808 24952 4820
rect 24907 4780 24952 4808
rect 24946 4768 24952 4780
rect 25004 4768 25010 4820
rect 26786 4808 26792 4820
rect 26747 4780 26792 4808
rect 26786 4768 26792 4780
rect 26844 4768 26850 4820
rect 27430 4808 27436 4820
rect 27391 4780 27436 4808
rect 27430 4768 27436 4780
rect 27488 4768 27494 4820
rect 29454 4768 29460 4820
rect 29512 4808 29518 4820
rect 30929 4811 30987 4817
rect 30929 4808 30941 4811
rect 29512 4780 30941 4808
rect 29512 4768 29518 4780
rect 30929 4777 30941 4780
rect 30975 4808 30987 4811
rect 34790 4808 34796 4820
rect 30975 4780 34796 4808
rect 30975 4777 30987 4780
rect 30929 4771 30987 4777
rect 34790 4768 34796 4780
rect 34848 4768 34854 4820
rect 37090 4768 37096 4820
rect 37148 4808 37154 4820
rect 37737 4811 37795 4817
rect 37737 4808 37749 4811
rect 37148 4780 37749 4808
rect 37148 4768 37154 4780
rect 37737 4777 37749 4780
rect 37783 4777 37795 4811
rect 37737 4771 37795 4777
rect 14369 4743 14427 4749
rect 14369 4709 14381 4743
rect 14415 4709 14427 4743
rect 20346 4740 20352 4752
rect 14369 4703 14427 4709
rect 14476 4712 20352 4740
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6052 4644 6745 4672
rect 6052 4632 6058 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 12618 4632 12624 4684
rect 12676 4672 12682 4684
rect 14476 4672 14504 4712
rect 20346 4700 20352 4712
rect 20404 4700 20410 4752
rect 20622 4700 20628 4752
rect 20680 4740 20686 4752
rect 20680 4712 22416 4740
rect 20680 4700 20686 4712
rect 17218 4672 17224 4684
rect 12676 4644 14504 4672
rect 15764 4644 17224 4672
rect 12676 4632 12682 4644
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 5166 4604 5172 4616
rect 5079 4576 5172 4604
rect 4893 4567 4951 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5442 4604 5448 4616
rect 5399 4576 5448 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 7006 4613 7012 4616
rect 7000 4604 7012 4613
rect 6967 4576 7012 4604
rect 7000 4567 7012 4576
rect 7006 4564 7012 4567
rect 7064 4564 7070 4616
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10505 4607 10563 4613
rect 10505 4604 10517 4607
rect 10376 4576 10517 4604
rect 10376 4564 10382 4576
rect 10505 4573 10517 4576
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10778 4604 10784 4616
rect 10739 4576 10784 4604
rect 10597 4567 10655 4573
rect 4709 4539 4767 4545
rect 4709 4536 4721 4539
rect 3988 4508 4721 4536
rect 4709 4505 4721 4508
rect 4755 4505 4767 4539
rect 5184 4536 5212 4564
rect 7466 4536 7472 4548
rect 5184 4508 7472 4536
rect 4709 4499 4767 4505
rect 7466 4496 7472 4508
rect 7524 4496 7530 4548
rect 10612 4536 10640 4567
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 10962 4604 10968 4616
rect 10919 4576 10968 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11698 4564 11704 4616
rect 11756 4604 11762 4616
rect 14292 4613 14320 4644
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 11756 4576 12541 4604
rect 11756 4564 11762 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 14277 4607 14335 4613
rect 12851 4576 14228 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 10686 4536 10692 4548
rect 10612 4508 10692 4536
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 3786 4468 3792 4480
rect 3747 4440 3792 4468
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 4028 4440 8953 4468
rect 4028 4428 4034 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 8941 4431 8999 4437
rect 13541 4471 13599 4477
rect 13541 4437 13553 4471
rect 13587 4468 13599 4471
rect 13630 4468 13636 4480
rect 13587 4440 13636 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13872 4440 14105 4468
rect 13872 4428 13878 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14200 4468 14228 4576
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14458 4604 14464 4616
rect 14419 4576 14464 4604
rect 14277 4567 14335 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4604 14611 4607
rect 14734 4604 14740 4616
rect 14599 4576 14740 4604
rect 14599 4573 14611 4576
rect 14553 4567 14611 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15102 4564 15108 4616
rect 15160 4604 15166 4616
rect 15764 4613 15792 4644
rect 16776 4616 16804 4644
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17954 4632 17960 4684
rect 18012 4672 18018 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 18012 4644 19257 4672
rect 18012 4632 18018 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4672 19579 4675
rect 21082 4672 21088 4684
rect 19567 4644 21088 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 21082 4632 21088 4644
rect 21140 4672 21146 4684
rect 22388 4672 22416 4712
rect 23106 4700 23112 4752
rect 23164 4740 23170 4752
rect 23569 4743 23627 4749
rect 23569 4740 23581 4743
rect 23164 4712 23581 4740
rect 23164 4700 23170 4712
rect 23569 4709 23581 4712
rect 23615 4709 23627 4743
rect 23569 4703 23627 4709
rect 24578 4700 24584 4752
rect 24636 4740 24642 4752
rect 25409 4743 25467 4749
rect 25409 4740 25421 4743
rect 24636 4712 25421 4740
rect 24636 4700 24642 4712
rect 25409 4709 25421 4712
rect 25455 4709 25467 4743
rect 25682 4740 25688 4752
rect 25643 4712 25688 4740
rect 25409 4703 25467 4709
rect 25682 4700 25688 4712
rect 25740 4700 25746 4752
rect 25774 4700 25780 4752
rect 25832 4740 25838 4752
rect 31662 4740 31668 4752
rect 25832 4712 25877 4740
rect 31623 4712 31668 4740
rect 25832 4700 25838 4712
rect 31662 4700 31668 4712
rect 31720 4700 31726 4752
rect 33965 4743 34023 4749
rect 33965 4709 33977 4743
rect 34011 4740 34023 4743
rect 34701 4743 34759 4749
rect 34701 4740 34713 4743
rect 34011 4712 34713 4740
rect 34011 4709 34023 4712
rect 33965 4703 34023 4709
rect 34701 4709 34713 4712
rect 34747 4709 34759 4743
rect 34701 4703 34759 4709
rect 24026 4672 24032 4684
rect 21140 4644 22048 4672
rect 21140 4632 21146 4644
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15160 4576 15761 4604
rect 15160 4564 15166 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 16025 4607 16083 4613
rect 15896 4576 15941 4604
rect 15896 4564 15902 4576
rect 16025 4573 16037 4607
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16758 4604 16764 4616
rect 16671 4576 16764 4604
rect 16117 4567 16175 4573
rect 14366 4496 14372 4548
rect 14424 4536 14430 4548
rect 16040 4536 16068 4567
rect 14424 4508 16068 4536
rect 16132 4536 16160 4567
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16850 4564 16856 4616
rect 16908 4604 16914 4616
rect 17034 4604 17040 4616
rect 16908 4576 16953 4604
rect 16995 4576 17040 4604
rect 16908 4564 16914 4576
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4573 17187 4607
rect 17236 4604 17264 4632
rect 17773 4607 17831 4613
rect 17773 4604 17785 4607
rect 17236 4576 17785 4604
rect 17129 4567 17187 4573
rect 17773 4573 17785 4576
rect 17819 4573 17831 4607
rect 17773 4567 17831 4573
rect 17144 4536 17172 4567
rect 17862 4564 17868 4616
rect 17920 4604 17926 4616
rect 18046 4604 18052 4616
rect 17920 4576 17965 4604
rect 18007 4576 18052 4604
rect 17920 4564 17926 4576
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4604 18199 4607
rect 18230 4604 18236 4616
rect 18187 4576 18236 4604
rect 18187 4573 18199 4576
rect 18141 4567 18199 4573
rect 17218 4536 17224 4548
rect 16132 4508 17224 4536
rect 14424 4496 14430 4508
rect 17218 4496 17224 4508
rect 17276 4536 17282 4548
rect 18156 4536 18184 4567
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 18782 4564 18788 4616
rect 18840 4604 18846 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 18840 4576 20729 4604
rect 18840 4564 18846 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20717 4567 20775 4573
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4604 21051 4607
rect 21542 4604 21548 4616
rect 21039 4576 21548 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 22020 4613 22048 4644
rect 22388 4644 24032 4672
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 22094 4564 22100 4616
rect 22152 4604 22158 4616
rect 22388 4613 22416 4644
rect 24026 4632 24032 4644
rect 24084 4672 24090 4684
rect 24084 4644 24808 4672
rect 24084 4632 24090 4644
rect 22281 4607 22339 4613
rect 22152 4576 22197 4604
rect 22152 4564 22158 4576
rect 22281 4573 22293 4607
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 17276 4508 18184 4536
rect 22296 4536 22324 4567
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 23477 4607 23535 4613
rect 23477 4604 23489 4607
rect 23440 4576 23489 4604
rect 23440 4564 23446 4576
rect 23477 4573 23489 4576
rect 23523 4573 23535 4607
rect 23658 4604 23664 4616
rect 23619 4576 23664 4604
rect 23477 4567 23535 4573
rect 22830 4536 22836 4548
rect 22296 4508 22836 4536
rect 17276 4496 17282 4508
rect 22830 4496 22836 4508
rect 22888 4496 22894 4548
rect 23492 4536 23520 4567
rect 23658 4564 23664 4576
rect 23716 4564 23722 4616
rect 23753 4607 23811 4613
rect 23753 4573 23765 4607
rect 23799 4604 23811 4607
rect 24210 4604 24216 4616
rect 23799 4576 24216 4604
rect 23799 4573 23811 4576
rect 23753 4567 23811 4573
rect 24210 4564 24216 4576
rect 24268 4564 24274 4616
rect 24302 4564 24308 4616
rect 24360 4604 24366 4616
rect 24397 4607 24455 4613
rect 24397 4604 24409 4607
rect 24360 4576 24409 4604
rect 24360 4564 24366 4576
rect 24397 4573 24409 4576
rect 24443 4573 24455 4607
rect 24397 4567 24455 4573
rect 24486 4564 24492 4616
rect 24544 4604 24550 4616
rect 24670 4604 24676 4616
rect 24544 4576 24589 4604
rect 24631 4576 24676 4604
rect 24544 4564 24550 4576
rect 24670 4564 24676 4576
rect 24728 4564 24734 4616
rect 24780 4613 24808 4644
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 25593 4607 25651 4613
rect 25593 4573 25605 4607
rect 25639 4573 25651 4607
rect 25593 4567 25651 4573
rect 25608 4536 25636 4567
rect 23492 4508 25636 4536
rect 18782 4468 18788 4480
rect 14200 4440 18788 4468
rect 14093 4431 14151 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 23658 4428 23664 4480
rect 23716 4468 23722 4480
rect 25792 4468 25820 4700
rect 28445 4675 28503 4681
rect 28445 4641 28457 4675
rect 28491 4672 28503 4675
rect 29178 4672 29184 4684
rect 28491 4644 29184 4672
rect 28491 4641 28503 4644
rect 28445 4635 28503 4641
rect 29178 4632 29184 4644
rect 29236 4632 29242 4684
rect 31294 4632 31300 4684
rect 31352 4672 31358 4684
rect 31389 4675 31447 4681
rect 31389 4672 31401 4675
rect 31352 4644 31401 4672
rect 31352 4632 31358 4644
rect 31389 4641 31401 4644
rect 31435 4672 31447 4675
rect 32309 4675 32367 4681
rect 32309 4672 32321 4675
rect 31435 4644 32321 4672
rect 31435 4641 31447 4644
rect 31389 4635 31447 4641
rect 32309 4641 32321 4644
rect 32355 4641 32367 4675
rect 32309 4635 32367 4641
rect 33597 4675 33655 4681
rect 33597 4641 33609 4675
rect 33643 4672 33655 4675
rect 33870 4672 33876 4684
rect 33643 4644 33876 4672
rect 33643 4641 33655 4644
rect 33597 4635 33655 4641
rect 33870 4632 33876 4644
rect 33928 4672 33934 4684
rect 34330 4672 34336 4684
rect 33928 4644 34336 4672
rect 33928 4632 33934 4644
rect 34330 4632 34336 4644
rect 34388 4632 34394 4684
rect 34606 4632 34612 4684
rect 34664 4672 34670 4684
rect 35253 4675 35311 4681
rect 35253 4672 35265 4675
rect 34664 4644 35265 4672
rect 34664 4632 34670 4644
rect 35253 4641 35265 4644
rect 35299 4641 35311 4675
rect 35253 4635 35311 4641
rect 35894 4632 35900 4684
rect 35952 4672 35958 4684
rect 36354 4672 36360 4684
rect 35952 4644 36360 4672
rect 35952 4632 35958 4644
rect 36354 4632 36360 4644
rect 36412 4632 36418 4684
rect 25866 4564 25872 4616
rect 25924 4604 25930 4616
rect 26418 4604 26424 4616
rect 25924 4576 25969 4604
rect 26379 4576 26424 4604
rect 25924 4564 25930 4576
rect 26418 4564 26424 4576
rect 26476 4564 26482 4616
rect 27706 4564 27712 4616
rect 27764 4604 27770 4616
rect 27801 4607 27859 4613
rect 27801 4604 27813 4607
rect 27764 4576 27813 4604
rect 27764 4564 27770 4576
rect 27801 4573 27813 4576
rect 27847 4573 27859 4607
rect 28534 4604 28540 4616
rect 27801 4567 27859 4573
rect 28368 4576 28540 4604
rect 26605 4539 26663 4545
rect 26605 4505 26617 4539
rect 26651 4536 26663 4539
rect 27617 4539 27675 4545
rect 26651 4508 27568 4536
rect 26651 4505 26663 4508
rect 26605 4499 26663 4505
rect 23716 4440 25820 4468
rect 27540 4468 27568 4508
rect 27617 4505 27629 4539
rect 27663 4536 27675 4539
rect 28368 4536 28396 4576
rect 28534 4564 28540 4576
rect 28592 4564 28598 4616
rect 28626 4564 28632 4616
rect 28684 4604 28690 4616
rect 29546 4604 29552 4616
rect 28684 4576 28729 4604
rect 29507 4576 29552 4604
rect 28684 4564 28690 4576
rect 29546 4564 29552 4576
rect 29604 4564 29610 4616
rect 29816 4607 29874 4613
rect 29816 4573 29828 4607
rect 29862 4604 29874 4607
rect 30190 4604 30196 4616
rect 29862 4576 30196 4604
rect 29862 4573 29874 4576
rect 29816 4567 29874 4573
rect 30190 4564 30196 4576
rect 30248 4564 30254 4616
rect 32953 4607 33011 4613
rect 32953 4573 32965 4607
rect 32999 4604 33011 4607
rect 33410 4604 33416 4616
rect 32999 4576 33416 4604
rect 32999 4573 33011 4576
rect 32953 4567 33011 4573
rect 33410 4564 33416 4576
rect 33468 4564 33474 4616
rect 36262 4564 36268 4616
rect 36320 4604 36326 4616
rect 36613 4607 36671 4613
rect 36613 4604 36625 4607
rect 36320 4576 36625 4604
rect 36320 4564 36326 4576
rect 36613 4573 36625 4576
rect 36659 4573 36671 4607
rect 36613 4567 36671 4573
rect 30282 4536 30288 4548
rect 27663 4508 28396 4536
rect 28460 4508 30288 4536
rect 27663 4505 27675 4508
rect 27617 4499 27675 4505
rect 28460 4468 28488 4508
rect 30282 4496 30288 4508
rect 30340 4496 30346 4548
rect 34606 4536 34612 4548
rect 33888 4508 34612 4536
rect 27540 4440 28488 4468
rect 23716 4428 23722 4440
rect 28534 4428 28540 4480
rect 28592 4468 28598 4480
rect 28994 4468 29000 4480
rect 28592 4440 28637 4468
rect 28955 4440 29000 4468
rect 28592 4428 28598 4440
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 31849 4471 31907 4477
rect 31849 4437 31861 4471
rect 31895 4468 31907 4471
rect 32122 4468 32128 4480
rect 31895 4440 32128 4468
rect 31895 4437 31907 4440
rect 31849 4431 31907 4437
rect 32122 4428 32128 4440
rect 32180 4428 32186 4480
rect 33137 4471 33195 4477
rect 33137 4437 33149 4471
rect 33183 4468 33195 4471
rect 33888 4468 33916 4508
rect 34606 4496 34612 4508
rect 34664 4496 34670 4548
rect 33183 4440 33916 4468
rect 33183 4437 33195 4440
rect 33137 4431 33195 4437
rect 33962 4428 33968 4480
rect 34020 4468 34026 4480
rect 34057 4471 34115 4477
rect 34057 4468 34069 4471
rect 34020 4440 34069 4468
rect 34020 4428 34026 4440
rect 34057 4437 34069 4440
rect 34103 4437 34115 4471
rect 34057 4431 34115 4437
rect 34422 4428 34428 4480
rect 34480 4468 34486 4480
rect 35069 4471 35127 4477
rect 35069 4468 35081 4471
rect 34480 4440 35081 4468
rect 34480 4428 34486 4440
rect 35069 4437 35081 4440
rect 35115 4437 35127 4471
rect 35069 4431 35127 4437
rect 35161 4471 35219 4477
rect 35161 4437 35173 4471
rect 35207 4468 35219 4471
rect 36078 4468 36084 4480
rect 35207 4440 36084 4468
rect 35207 4437 35219 4440
rect 35161 4431 35219 4437
rect 36078 4428 36084 4440
rect 36136 4428 36142 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 6638 4224 6644 4276
rect 6696 4264 6702 4276
rect 10778 4264 10784 4276
rect 6696 4236 10784 4264
rect 6696 4224 6702 4236
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 10962 4224 10968 4276
rect 11020 4224 11026 4276
rect 13357 4267 13415 4273
rect 13357 4233 13369 4267
rect 13403 4264 13415 4267
rect 13538 4264 13544 4276
rect 13403 4236 13544 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 13630 4224 13636 4276
rect 13688 4264 13694 4276
rect 23106 4264 23112 4276
rect 13688 4236 23112 4264
rect 13688 4224 13694 4236
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 24302 4224 24308 4276
rect 24360 4224 24366 4276
rect 26329 4267 26387 4273
rect 26329 4233 26341 4267
rect 26375 4264 26387 4267
rect 26418 4264 26424 4276
rect 26375 4236 26424 4264
rect 26375 4233 26387 4236
rect 26329 4227 26387 4233
rect 26418 4224 26424 4236
rect 26476 4224 26482 4276
rect 27890 4224 27896 4276
rect 27948 4264 27954 4276
rect 28626 4264 28632 4276
rect 27948 4236 28632 4264
rect 27948 4224 27954 4236
rect 28626 4224 28632 4236
rect 28684 4224 28690 4276
rect 31113 4267 31171 4273
rect 31113 4233 31125 4267
rect 31159 4264 31171 4267
rect 31662 4264 31668 4276
rect 31159 4236 31668 4264
rect 31159 4233 31171 4236
rect 31113 4227 31171 4233
rect 31662 4224 31668 4236
rect 31720 4224 31726 4276
rect 35526 4224 35532 4276
rect 35584 4264 35590 4276
rect 35713 4267 35771 4273
rect 35713 4264 35725 4267
rect 35584 4236 35725 4264
rect 35584 4224 35590 4236
rect 35713 4233 35725 4236
rect 35759 4233 35771 4267
rect 35713 4227 35771 4233
rect 3320 4199 3378 4205
rect 3320 4165 3332 4199
rect 3366 4196 3378 4199
rect 3786 4196 3792 4208
rect 3366 4168 3792 4196
rect 3366 4165 3378 4168
rect 3320 4159 3378 4165
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 7098 4196 7104 4208
rect 4212 4168 7104 4196
rect 4212 4156 4218 4168
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 2314 4128 2320 4140
rect 1443 4100 2320 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2556 4100 2605 4128
rect 2556 4088 2562 4100
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 5074 4128 5080 4140
rect 2593 4091 2651 4097
rect 2746 4100 4108 4128
rect 5035 4100 5080 4128
rect 2130 4060 2136 4072
rect 2091 4032 2136 4060
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 2746 3992 2774 4100
rect 3050 4060 3056 4072
rect 3011 4032 3056 4060
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 4080 4060 4108 4100
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5276 4137 5304 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 7558 4196 7564 4208
rect 7208 4168 7564 4196
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7208 4137 7236 4168
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 10980 4196 11008 4224
rect 23382 4196 23388 4208
rect 10796 4168 11008 4196
rect 13464 4168 13676 4196
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6972 4100 7021 4128
rect 6972 4088 6978 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7193 4091 7251 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 5353 4063 5411 4069
rect 5353 4060 5365 4063
rect 4080 4032 5365 4060
rect 5353 4029 5365 4032
rect 5399 4060 5411 4063
rect 5399 4032 7144 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 1820 3964 2774 3992
rect 4433 3995 4491 4001
rect 1820 3952 1826 3964
rect 4433 3961 4445 3995
rect 4479 3992 4491 3995
rect 5442 3992 5448 4004
rect 4479 3964 5448 3992
rect 4479 3961 4491 3964
rect 4433 3955 4491 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 2958 3924 2964 3936
rect 2547 3896 2964 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 4890 3924 4896 3936
rect 4851 3896 4896 3924
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5776 3896 6377 3924
rect 5776 3884 5782 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 7116 3924 7144 4032
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 7668 4060 7696 4091
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 9217 4131 9275 4137
rect 9217 4128 9229 4131
rect 7892 4100 9229 4128
rect 7892 4088 7898 4100
rect 9217 4097 9229 4100
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10376 4100 10425 4128
rect 10376 4088 10382 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10796 4137 10824 4168
rect 10689 4131 10747 4137
rect 10560 4100 10605 4128
rect 10560 4088 10566 4100
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 11422 4128 11428 4140
rect 11011 4100 11428 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 10704 4060 10732 4091
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 13464 4128 13492 4168
rect 13648 4137 13676 4168
rect 16500 4168 17448 4196
rect 11532 4100 13492 4128
rect 13541 4131 13599 4137
rect 7432 4032 10732 4060
rect 7432 4020 7438 4032
rect 8202 3924 8208 3936
rect 7116 3896 8208 3924
rect 6365 3887 6423 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8352 3896 8677 3924
rect 8352 3884 8358 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 11532 3924 11560 4100
rect 13541 4097 13553 4131
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 13814 4128 13820 4140
rect 13775 4100 13820 4128
rect 13633 4091 13691 4097
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4060 11667 4063
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11655 4032 12081 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12342 4060 12348 4072
rect 12303 4032 12348 4060
rect 12069 4023 12127 4029
rect 8812 3896 11560 3924
rect 12084 3924 12112 4023
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 13556 3992 13584 4091
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 15286 4128 15292 4140
rect 13955 4100 15292 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 16500 4128 16528 4168
rect 16666 4128 16672 4140
rect 16132 4100 16528 4128
rect 16627 4100 16672 4128
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14240 4032 14381 4060
rect 14240 4020 14246 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 16132 4060 16160 4100
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16816 4100 16865 4128
rect 16816 4088 16822 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 17126 4128 17132 4140
rect 17087 4100 17132 4128
rect 16945 4091 17003 4097
rect 14884 4032 16160 4060
rect 14884 4020 14890 4032
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 16960 4060 16988 4091
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17420 4128 17448 4168
rect 23032 4168 23388 4196
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17276 4100 17321 4128
rect 17420 4100 17969 4128
rect 17276 4088 17282 4100
rect 17957 4097 17969 4100
rect 18003 4128 18015 4131
rect 19245 4131 19303 4137
rect 19245 4128 19257 4131
rect 18003 4100 19257 4128
rect 18003 4097 18015 4100
rect 17957 4091 18015 4097
rect 19245 4097 19257 4100
rect 19291 4097 19303 4131
rect 20622 4128 20628 4140
rect 19245 4091 19303 4097
rect 19720 4100 20628 4128
rect 18966 4060 18972 4072
rect 16448 4032 16988 4060
rect 18927 4032 18972 4060
rect 16448 4020 16454 4032
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 19058 4020 19064 4072
rect 19116 4060 19122 4072
rect 19720 4069 19748 4100
rect 20622 4088 20628 4100
rect 20680 4128 20686 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20680 4100 21005 4128
rect 20680 4088 20686 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 23032 4137 23060 4168
rect 23382 4156 23388 4168
rect 23440 4156 23446 4208
rect 24320 4196 24348 4224
rect 28353 4199 28411 4205
rect 24320 4168 24440 4196
rect 22833 4131 22891 4137
rect 22833 4128 22845 4131
rect 22796 4100 22845 4128
rect 22796 4088 22802 4100
rect 22833 4097 22845 4100
rect 22879 4097 22891 4131
rect 22833 4091 22891 4097
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 23293 4131 23351 4137
rect 23164 4100 23209 4128
rect 23164 4088 23170 4100
rect 23293 4097 23305 4131
rect 23339 4128 23351 4131
rect 23842 4128 23848 4140
rect 23339 4100 23704 4128
rect 23803 4100 23848 4128
rect 23339 4097 23351 4100
rect 23293 4091 23351 4097
rect 19705 4063 19763 4069
rect 19705 4060 19717 4063
rect 19116 4032 19717 4060
rect 19116 4020 19122 4032
rect 19705 4029 19717 4032
rect 19751 4029 19763 4063
rect 19978 4060 19984 4072
rect 19939 4032 19984 4060
rect 19705 4023 19763 4029
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 20088 4032 22385 4060
rect 14200 3992 14228 4020
rect 13556 3964 14228 3992
rect 14458 3952 14464 4004
rect 14516 3992 14522 4004
rect 20088 3992 20116 4032
rect 22373 4029 22385 4032
rect 22419 4060 22431 4063
rect 23198 4060 23204 4072
rect 22419 4032 23204 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 14516 3964 20116 3992
rect 14516 3952 14522 3964
rect 21542 3952 21548 4004
rect 21600 3992 21606 4004
rect 22554 3992 22560 4004
rect 21600 3964 22560 3992
rect 21600 3952 21606 3964
rect 22554 3952 22560 3964
rect 22612 3952 22618 4004
rect 14826 3924 14832 3936
rect 12084 3896 14832 3924
rect 8812 3884 8818 3896
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16942 3924 16948 3936
rect 16724 3896 16948 3924
rect 16724 3884 16730 3896
rect 16942 3884 16948 3896
rect 17000 3924 17006 3936
rect 17678 3924 17684 3936
rect 17000 3896 17684 3924
rect 17000 3884 17006 3896
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 23198 3924 23204 3936
rect 17828 3896 23204 3924
rect 17828 3884 17834 3896
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 23676 3924 23704 4100
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 24026 4128 24032 4140
rect 23987 4100 24032 4128
rect 24026 4088 24032 4100
rect 24084 4088 24090 4140
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 24412 4137 24440 4168
rect 28353 4165 28365 4199
rect 28399 4196 28411 4199
rect 29086 4196 29092 4208
rect 28399 4168 29092 4196
rect 28399 4165 28411 4168
rect 28353 4159 28411 4165
rect 29086 4156 29092 4168
rect 29144 4156 29150 4208
rect 29822 4156 29828 4208
rect 29880 4196 29886 4208
rect 30745 4199 30803 4205
rect 30745 4196 30757 4199
rect 29880 4168 30757 4196
rect 29880 4156 29886 4168
rect 30745 4165 30757 4168
rect 30791 4196 30803 4199
rect 34422 4196 34428 4208
rect 30791 4168 34428 4196
rect 30791 4165 30803 4168
rect 30745 4159 30803 4165
rect 34422 4156 34428 4168
rect 34480 4156 34486 4208
rect 24305 4131 24363 4137
rect 24176 4100 24221 4128
rect 24176 4088 24182 4100
rect 24305 4097 24317 4131
rect 24351 4097 24363 4131
rect 24305 4091 24363 4097
rect 24397 4131 24455 4137
rect 24397 4097 24409 4131
rect 24443 4097 24455 4131
rect 24854 4128 24860 4140
rect 24815 4100 24860 4128
rect 24397 4091 24455 4097
rect 24320 4060 24348 4091
rect 24854 4088 24860 4100
rect 24912 4088 24918 4140
rect 25038 4128 25044 4140
rect 24999 4100 25044 4128
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 28902 4128 28908 4140
rect 25363 4100 28908 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 29273 4131 29331 4137
rect 29273 4097 29285 4131
rect 29319 4097 29331 4131
rect 29273 4091 29331 4097
rect 25406 4060 25412 4072
rect 24320 4032 25412 4060
rect 25406 4020 25412 4032
rect 25464 4020 25470 4072
rect 28813 4063 28871 4069
rect 28813 4029 28825 4063
rect 28859 4060 28871 4063
rect 29288 4060 29316 4091
rect 30282 4088 30288 4140
rect 30340 4128 30346 4140
rect 30653 4131 30711 4137
rect 30653 4128 30665 4131
rect 30340 4100 30665 4128
rect 30340 4088 30346 4100
rect 30653 4097 30665 4100
rect 30699 4097 30711 4131
rect 32122 4128 32128 4140
rect 32083 4100 32128 4128
rect 30653 4091 30711 4097
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 32766 4088 32772 4140
rect 32824 4128 32830 4140
rect 34606 4137 34612 4140
rect 32861 4131 32919 4137
rect 32861 4128 32873 4131
rect 32824 4100 32873 4128
rect 32824 4088 32830 4100
rect 32861 4097 32873 4100
rect 32907 4128 32919 4131
rect 34333 4131 34391 4137
rect 34333 4128 34345 4131
rect 32907 4100 34345 4128
rect 32907 4097 32919 4100
rect 32861 4091 32919 4097
rect 34333 4097 34345 4100
rect 34379 4097 34391 4131
rect 34600 4128 34612 4137
rect 34567 4100 34612 4128
rect 34333 4091 34391 4097
rect 34600 4091 34612 4100
rect 34606 4088 34612 4091
rect 34664 4088 34670 4140
rect 35728 4128 35756 4227
rect 37826 4224 37832 4276
rect 37884 4224 37890 4276
rect 37734 4196 37740 4208
rect 37695 4168 37740 4196
rect 37734 4156 37740 4168
rect 37792 4156 37798 4208
rect 37844 4196 37872 4224
rect 37844 4168 38056 4196
rect 37550 4137 37556 4140
rect 36449 4131 36507 4137
rect 36449 4128 36461 4131
rect 35728 4100 36461 4128
rect 36449 4097 36461 4100
rect 36495 4097 36507 4131
rect 37548 4128 37556 4137
rect 37511 4100 37556 4128
rect 36449 4091 36507 4097
rect 37548 4091 37556 4100
rect 37550 4088 37556 4091
rect 37608 4088 37614 4140
rect 37645 4131 37703 4137
rect 37645 4097 37657 4131
rect 37691 4097 37703 4131
rect 37645 4091 37703 4097
rect 28859 4032 29316 4060
rect 28859 4029 28871 4032
rect 28813 4023 28871 4029
rect 30098 4020 30104 4072
rect 30156 4060 30162 4072
rect 30469 4063 30527 4069
rect 30469 4060 30481 4063
rect 30156 4032 30481 4060
rect 30156 4020 30162 4032
rect 30469 4029 30481 4032
rect 30515 4029 30527 4063
rect 33410 4060 33416 4072
rect 33371 4032 33416 4060
rect 30469 4023 30527 4029
rect 33410 4020 33416 4032
rect 33468 4020 33474 4072
rect 33870 4060 33876 4072
rect 33831 4032 33876 4060
rect 33870 4020 33876 4032
rect 33928 4020 33934 4072
rect 36078 4020 36084 4072
rect 36136 4060 36142 4072
rect 37660 4060 37688 4091
rect 37826 4088 37832 4140
rect 37884 4137 37890 4140
rect 38028 4137 38056 4168
rect 37884 4131 37923 4137
rect 37911 4097 37923 4131
rect 37884 4091 37923 4097
rect 38013 4131 38071 4137
rect 38013 4097 38025 4131
rect 38059 4097 38071 4131
rect 38013 4091 38071 4097
rect 37884 4088 37890 4091
rect 36136 4032 37688 4060
rect 36136 4020 36142 4032
rect 25130 3992 25136 4004
rect 25091 3964 25136 3992
rect 25130 3952 25136 3964
rect 25188 3952 25194 4004
rect 25222 3952 25228 4004
rect 25280 3992 25286 4004
rect 28721 3995 28779 4001
rect 25280 3964 25325 3992
rect 27724 3964 28672 3992
rect 25280 3952 25286 3964
rect 27724 3924 27752 3964
rect 27890 3924 27896 3936
rect 23676 3896 27752 3924
rect 27851 3896 27896 3924
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 28644 3924 28672 3964
rect 28721 3961 28733 3995
rect 28767 3992 28779 3995
rect 28994 3992 29000 4004
rect 28767 3964 29000 3992
rect 28767 3961 28779 3964
rect 28721 3955 28779 3961
rect 28994 3952 29000 3964
rect 29052 3952 29058 4004
rect 31202 3992 31208 4004
rect 29288 3964 31208 3992
rect 29288 3924 29316 3964
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 33594 3992 33600 4004
rect 33555 3964 33600 3992
rect 33594 3952 33600 3964
rect 33652 3952 33658 4004
rect 37366 3992 37372 4004
rect 37327 3964 37372 3992
rect 37366 3952 37372 3964
rect 37424 3952 37430 4004
rect 29454 3924 29460 3936
rect 28644 3896 29316 3924
rect 29415 3896 29460 3924
rect 29454 3884 29460 3896
rect 29512 3884 29518 3936
rect 32306 3924 32312 3936
rect 32267 3896 32312 3924
rect 32306 3884 32312 3896
rect 32364 3884 32370 3936
rect 32858 3884 32864 3936
rect 32916 3924 32922 3936
rect 35710 3924 35716 3936
rect 32916 3896 35716 3924
rect 32916 3884 32922 3896
rect 35710 3884 35716 3896
rect 35768 3884 35774 3936
rect 36630 3924 36636 3936
rect 36591 3896 36636 3924
rect 36630 3884 36636 3896
rect 36688 3884 36694 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1762 3720 1768 3732
rect 1723 3692 1768 3720
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3418 3720 3424 3732
rect 2823 3692 3424 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5534 3720 5540 3732
rect 5215 3692 5540 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5534 3680 5540 3692
rect 5592 3720 5598 3732
rect 6638 3720 6644 3732
rect 5592 3692 6644 3720
rect 5592 3680 5598 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7374 3720 7380 3732
rect 7335 3692 7380 3720
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10410 3720 10416 3732
rect 9907 3692 10416 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10744 3692 10885 3720
rect 10744 3680 10750 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 12894 3720 12900 3732
rect 12855 3692 12900 3720
rect 10873 3683 10931 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 15197 3723 15255 3729
rect 15197 3689 15209 3723
rect 15243 3720 15255 3723
rect 15470 3720 15476 3732
rect 15243 3692 15476 3720
rect 15243 3689 15255 3692
rect 15197 3683 15255 3689
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 16666 3720 16672 3732
rect 16627 3692 16672 3720
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 17092 3692 17141 3720
rect 17092 3680 17098 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18104 3692 18153 3720
rect 18104 3680 18110 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 22189 3723 22247 3729
rect 22189 3720 22201 3723
rect 22152 3692 22201 3720
rect 22152 3680 22158 3692
rect 22189 3689 22201 3692
rect 22235 3689 22247 3723
rect 22189 3683 22247 3689
rect 23106 3680 23112 3732
rect 23164 3720 23170 3732
rect 23293 3723 23351 3729
rect 23293 3720 23305 3723
rect 23164 3692 23305 3720
rect 23164 3680 23170 3692
rect 23293 3689 23305 3692
rect 23339 3689 23351 3723
rect 23293 3683 23351 3689
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 23716 3692 23765 3720
rect 23716 3680 23722 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 23753 3683 23811 3689
rect 24486 3680 24492 3732
rect 24544 3720 24550 3732
rect 24949 3723 25007 3729
rect 24949 3720 24961 3723
rect 24544 3692 24961 3720
rect 24544 3680 24550 3692
rect 24949 3689 24961 3692
rect 24995 3689 25007 3723
rect 25406 3720 25412 3732
rect 25367 3692 25412 3720
rect 24949 3683 25007 3689
rect 25406 3680 25412 3692
rect 25464 3680 25470 3732
rect 29362 3680 29368 3732
rect 29420 3720 29426 3732
rect 29549 3723 29607 3729
rect 29549 3720 29561 3723
rect 29420 3692 29561 3720
rect 29420 3680 29426 3692
rect 29549 3689 29561 3692
rect 29595 3689 29607 3723
rect 29549 3683 29607 3689
rect 29822 3680 29828 3732
rect 29880 3720 29886 3732
rect 30193 3723 30251 3729
rect 30193 3720 30205 3723
rect 29880 3692 30205 3720
rect 29880 3680 29886 3692
rect 30193 3689 30205 3692
rect 30239 3689 30251 3723
rect 30193 3683 30251 3689
rect 30282 3680 30288 3732
rect 30340 3720 30346 3732
rect 31021 3723 31079 3729
rect 31021 3720 31033 3723
rect 30340 3692 31033 3720
rect 30340 3680 30346 3692
rect 31021 3689 31033 3692
rect 31067 3689 31079 3723
rect 31021 3683 31079 3689
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 10318 3652 10324 3664
rect 8260 3624 10324 3652
rect 8260 3612 8266 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 10597 3655 10655 3661
rect 10597 3621 10609 3655
rect 10643 3652 10655 3655
rect 22554 3652 22560 3664
rect 10643 3624 10732 3652
rect 22515 3624 22560 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 5994 3584 6000 3596
rect 5955 3556 6000 3584
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 10505 3587 10563 3593
rect 7064 3556 10456 3584
rect 7064 3544 7070 3556
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2498 3516 2504 3528
rect 2363 3488 2504 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 2958 3516 2964 3528
rect 2871 3488 2964 3516
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3108 3488 3801 3516
rect 3108 3476 3114 3488
rect 3789 3485 3801 3488
rect 3835 3516 3847 3519
rect 6012 3516 6040 3544
rect 6270 3525 6276 3528
rect 6264 3516 6276 3525
rect 3835 3488 6040 3516
rect 6231 3488 6276 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 6264 3479 6276 3488
rect 6270 3476 6276 3479
rect 6328 3476 6334 3528
rect 7834 3516 7840 3528
rect 6380 3488 7840 3516
rect 1394 3408 1400 3460
rect 1452 3448 1458 3460
rect 1489 3451 1547 3457
rect 1489 3448 1501 3451
rect 1452 3420 1501 3448
rect 1452 3408 1458 3420
rect 1489 3417 1501 3420
rect 1535 3448 1547 3451
rect 2976 3448 3004 3476
rect 6380 3460 6408 3488
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 8036 3488 9413 3516
rect 3878 3448 3884 3460
rect 1535 3420 2774 3448
rect 2976 3420 3884 3448
rect 1535 3417 1547 3420
rect 1489 3411 1547 3417
rect 2746 3380 2774 3420
rect 3878 3408 3884 3420
rect 3936 3408 3942 3460
rect 4056 3451 4114 3457
rect 4056 3417 4068 3451
rect 4102 3448 4114 3451
rect 4890 3448 4896 3460
rect 4102 3420 4896 3448
rect 4102 3417 4114 3420
rect 4056 3411 4114 3417
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 6362 3408 6368 3460
rect 6420 3408 6426 3460
rect 4706 3380 4712 3392
rect 2746 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 8036 3389 8064 3488
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3349 8079 3383
rect 9508 3380 9536 3479
rect 9600 3448 9628 3479
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 10428 3525 10456 3556
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10704 3584 10732 3624
rect 22554 3612 22560 3624
rect 22612 3652 22618 3664
rect 24581 3655 24639 3661
rect 24581 3652 24593 3655
rect 22612 3624 24593 3652
rect 22612 3612 22618 3624
rect 24581 3621 24593 3624
rect 24627 3652 24639 3655
rect 25222 3652 25228 3664
rect 24627 3624 25228 3652
rect 24627 3621 24639 3624
rect 24581 3615 24639 3621
rect 25222 3612 25228 3624
rect 25280 3612 25286 3664
rect 25774 3612 25780 3664
rect 25832 3652 25838 3664
rect 26973 3655 27031 3661
rect 26973 3652 26985 3655
rect 25832 3624 26985 3652
rect 25832 3612 25838 3624
rect 26973 3621 26985 3624
rect 27019 3621 27031 3655
rect 26973 3615 27031 3621
rect 10962 3584 10968 3596
rect 10704 3556 10968 3584
rect 10505 3547 10563 3553
rect 10413 3519 10471 3525
rect 9732 3488 9777 3516
rect 9732 3476 9738 3488
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10318 3448 10324 3460
rect 9600 3420 10324 3448
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 10520 3380 10548 3547
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3584 11575 3587
rect 12894 3584 12900 3596
rect 11563 3556 12900 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 17402 3584 17408 3596
rect 17363 3556 17408 3584
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 18509 3587 18567 3593
rect 18509 3584 18521 3587
rect 17512 3556 18521 3584
rect 10778 3525 10784 3528
rect 10721 3519 10784 3525
rect 10721 3485 10733 3519
rect 10767 3485 10784 3519
rect 10721 3479 10784 3485
rect 10778 3476 10784 3479
rect 10836 3476 10842 3528
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 17512 3525 17540 3556
rect 18509 3553 18521 3556
rect 18555 3584 18567 3587
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 18555 3556 19533 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 19521 3547 19579 3553
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 20947 3556 22477 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 22465 3553 22477 3556
rect 22511 3584 22523 3587
rect 24673 3587 24731 3593
rect 24673 3584 24685 3587
rect 22511 3556 24685 3584
rect 22511 3553 22523 3556
rect 22465 3547 22523 3553
rect 24673 3553 24685 3556
rect 24719 3584 24731 3587
rect 25130 3584 25136 3596
rect 24719 3556 25136 3584
rect 24719 3553 24731 3556
rect 24673 3547 24731 3553
rect 25130 3544 25136 3556
rect 25188 3584 25194 3596
rect 25685 3587 25743 3593
rect 25685 3584 25697 3587
rect 25188 3556 25697 3584
rect 25188 3544 25194 3556
rect 25685 3553 25697 3556
rect 25731 3553 25743 3587
rect 25685 3547 25743 3553
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3516 17371 3519
rect 17497 3519 17555 3525
rect 17359 3488 17448 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 12492 3420 13216 3448
rect 12492 3408 12498 3420
rect 13188 3392 13216 3420
rect 17420 3392 17448 3488
rect 17497 3485 17509 3519
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17512 3448 17540 3479
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 18325 3519 18383 3525
rect 17644 3488 17689 3516
rect 17644 3476 17650 3488
rect 18325 3485 18337 3519
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 17678 3448 17684 3460
rect 17512 3420 17684 3448
rect 17678 3408 17684 3420
rect 17736 3408 17742 3460
rect 18340 3448 18368 3479
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18472 3488 18517 3516
rect 18472 3476 18478 3488
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 18656 3488 18701 3516
rect 18656 3476 18662 3488
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 18840 3488 19257 3516
rect 18840 3476 18846 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 22370 3516 22376 3528
rect 22331 3488 22376 3516
rect 19245 3479 19303 3485
rect 22370 3476 22376 3488
rect 22428 3476 22434 3528
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3516 22707 3519
rect 22738 3516 22744 3528
rect 22695 3488 22744 3516
rect 22695 3485 22707 3488
rect 22649 3479 22707 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24489 3519 24547 3525
rect 24489 3516 24501 3519
rect 24268 3488 24501 3516
rect 24268 3476 24274 3488
rect 24489 3485 24501 3488
rect 24535 3485 24547 3519
rect 24489 3479 24547 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 25038 3516 25044 3528
rect 24811 3488 25044 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 18966 3448 18972 3460
rect 18340 3420 18972 3448
rect 10686 3380 10692 3392
rect 9508 3352 10692 3380
rect 8021 3343 8079 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 13228 3352 13369 3380
rect 13228 3340 13234 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 18340 3380 18368 3420
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 22388 3448 22416 3476
rect 24780 3448 24808 3479
rect 25038 3476 25044 3488
rect 25096 3516 25102 3528
rect 25593 3519 25651 3525
rect 25593 3516 25605 3519
rect 25096 3488 25605 3516
rect 25096 3476 25102 3488
rect 25593 3485 25605 3488
rect 25639 3485 25651 3519
rect 25593 3479 25651 3485
rect 25777 3519 25835 3525
rect 25777 3485 25789 3519
rect 25823 3485 25835 3519
rect 25777 3479 25835 3485
rect 25869 3519 25927 3525
rect 25869 3485 25881 3519
rect 25915 3516 25927 3519
rect 26970 3516 26976 3528
rect 25915 3488 26976 3516
rect 25915 3485 25927 3488
rect 25869 3479 25927 3485
rect 22388 3420 24808 3448
rect 25222 3408 25228 3460
rect 25280 3448 25286 3460
rect 25792 3448 25820 3479
rect 26970 3476 26976 3488
rect 27028 3476 27034 3528
rect 28353 3519 28411 3525
rect 28353 3485 28365 3519
rect 28399 3516 28411 3519
rect 28718 3516 28724 3528
rect 28399 3488 28724 3516
rect 28399 3485 28411 3488
rect 28353 3479 28411 3485
rect 28718 3476 28724 3488
rect 28776 3516 28782 3528
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 28776 3488 29009 3516
rect 28776 3476 28782 3488
rect 28997 3485 29009 3488
rect 29043 3485 29055 3519
rect 28997 3479 29055 3485
rect 27890 3448 27896 3460
rect 25280 3420 25820 3448
rect 26160 3420 27896 3448
rect 25280 3408 25286 3420
rect 17460 3352 18368 3380
rect 17460 3340 17466 3352
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 20622 3380 20628 3392
rect 18564 3352 20628 3380
rect 18564 3340 18570 3352
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 26160 3380 26188 3420
rect 27890 3408 27896 3420
rect 27948 3408 27954 3460
rect 23256 3352 26188 3380
rect 23256 3340 23262 3352
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 26421 3383 26479 3389
rect 26421 3380 26433 3383
rect 26292 3352 26433 3380
rect 26292 3340 26298 3352
rect 26421 3349 26433 3352
rect 26467 3349 26479 3383
rect 28810 3380 28816 3392
rect 28771 3352 28816 3380
rect 26421 3343 26479 3349
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 31036 3380 31064 3683
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 32861 3723 32919 3729
rect 32861 3720 32873 3723
rect 32824 3692 32873 3720
rect 32824 3680 32830 3692
rect 32861 3689 32873 3692
rect 32907 3720 32919 3723
rect 33413 3723 33471 3729
rect 33413 3720 33425 3723
rect 32907 3692 33425 3720
rect 32907 3689 32919 3692
rect 32861 3683 32919 3689
rect 33413 3689 33425 3692
rect 33459 3689 33471 3723
rect 36078 3720 36084 3732
rect 36039 3692 36084 3720
rect 33413 3683 33471 3689
rect 32401 3587 32459 3593
rect 32401 3553 32413 3587
rect 32447 3584 32459 3587
rect 32784 3584 32812 3680
rect 32447 3556 32812 3584
rect 33428 3584 33456 3683
rect 36078 3680 36084 3692
rect 36136 3680 36142 3732
rect 36354 3680 36360 3732
rect 36412 3720 36418 3732
rect 36541 3723 36599 3729
rect 36541 3720 36553 3723
rect 36412 3692 36553 3720
rect 36412 3680 36418 3692
rect 36541 3689 36553 3692
rect 36587 3689 36599 3723
rect 36541 3683 36599 3689
rect 34146 3652 34152 3664
rect 34107 3624 34152 3652
rect 34146 3612 34152 3624
rect 34204 3612 34210 3664
rect 34701 3587 34759 3593
rect 34701 3584 34713 3587
rect 33428 3556 34713 3584
rect 32447 3553 32459 3556
rect 32401 3547 32459 3553
rect 34701 3553 34713 3556
rect 34747 3553 34759 3587
rect 34701 3547 34759 3553
rect 32145 3519 32203 3525
rect 32145 3485 32157 3519
rect 32191 3516 32203 3519
rect 32306 3516 32312 3528
rect 32191 3488 32312 3516
rect 32191 3485 32203 3488
rect 32145 3479 32203 3485
rect 32306 3476 32312 3488
rect 32364 3476 32370 3528
rect 33962 3516 33968 3528
rect 33923 3488 33968 3516
rect 33962 3476 33968 3488
rect 34020 3476 34026 3528
rect 37093 3519 37151 3525
rect 37093 3516 37105 3519
rect 34072 3488 37105 3516
rect 31110 3408 31116 3460
rect 31168 3448 31174 3460
rect 34072 3448 34100 3488
rect 37093 3485 37105 3488
rect 37139 3485 37151 3519
rect 37093 3479 37151 3485
rect 37829 3519 37887 3525
rect 37829 3485 37841 3519
rect 37875 3485 37887 3519
rect 37829 3479 37887 3485
rect 31168 3420 34100 3448
rect 31168 3408 31174 3420
rect 34146 3408 34152 3460
rect 34204 3448 34210 3460
rect 34946 3451 35004 3457
rect 34946 3448 34958 3451
rect 34204 3420 34958 3448
rect 34204 3408 34210 3420
rect 34946 3417 34958 3420
rect 34992 3417 35004 3451
rect 37844 3448 37872 3479
rect 34946 3411 35004 3417
rect 35084 3420 37872 3448
rect 35084 3380 35112 3420
rect 37274 3380 37280 3392
rect 31036 3352 35112 3380
rect 37235 3352 37280 3380
rect 37274 3340 37280 3352
rect 37332 3340 37338 3392
rect 38010 3380 38016 3392
rect 37971 3352 38016 3380
rect 38010 3340 38016 3352
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 4614 3176 4620 3188
rect 3200 3148 4620 3176
rect 3200 3136 3206 3148
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 8021 3179 8079 3185
rect 4764 3148 7880 3176
rect 4764 3136 4770 3148
rect 1578 3068 1584 3120
rect 1636 3108 1642 3120
rect 7006 3108 7012 3120
rect 1636 3080 7012 3108
rect 1636 3068 1642 3080
rect 7006 3068 7012 3080
rect 7064 3068 7070 3120
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 3234 3040 3240 3052
rect 3195 3012 3240 3040
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 4249 3043 4307 3049
rect 3436 3012 3703 3040
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2774 2972 2780 2984
rect 2271 2944 2780 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2774 2932 2780 2944
rect 2832 2972 2838 2984
rect 3142 2972 3148 2984
rect 2832 2944 3148 2972
rect 2832 2932 2838 2944
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 1578 2864 1584 2916
rect 1636 2904 1642 2916
rect 3436 2904 3464 3012
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 3675 2972 3703 3012
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 5166 3040 5172 3052
rect 4295 3012 5172 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 5316 3012 5365 3040
rect 5316 3000 5322 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 6638 3040 6644 3052
rect 5500 3012 5672 3040
rect 6599 3012 6644 3040
rect 5500 3000 5506 3012
rect 5534 2972 5540 2984
rect 3568 2944 3613 2972
rect 3675 2944 5540 2972
rect 3568 2932 3574 2944
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5644 2972 5672 3012
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7852 3049 7880 3148
rect 8021 3145 8033 3179
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8036 3108 8064 3139
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10560 3148 10885 3176
rect 10560 3136 10566 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 10873 3139 10931 3145
rect 12069 3179 12127 3185
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 13262 3176 13268 3188
rect 12115 3148 13268 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 14737 3179 14795 3185
rect 14737 3145 14749 3179
rect 14783 3145 14795 3179
rect 14737 3139 14795 3145
rect 13817 3111 13875 3117
rect 13817 3108 13829 3111
rect 8036 3080 10088 3108
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8294 3040 8300 3052
rect 7883 3012 8300 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 8444 3012 8493 3040
rect 8444 3000 8450 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 8481 3003 8539 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 10060 3040 10088 3080
rect 10704 3080 11928 3108
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10060 3012 10425 3040
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10594 3040 10600 3052
rect 10555 3012 10600 3040
rect 10413 3003 10471 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10704 3049 10732 3080
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10778 3040 10784 3052
rect 10735 3012 10784 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11609 3043 11667 3049
rect 11609 3009 11621 3043
rect 11655 3009 11667 3043
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 11609 3003 11667 3009
rect 11624 2972 11652 3003
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11900 3049 11928 3080
rect 12728 3080 13829 3108
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12342 3040 12348 3052
rect 11931 3012 12348 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12728 3049 12756 3080
rect 13817 3077 13829 3080
rect 13863 3077 13875 3111
rect 14752 3108 14780 3139
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17221 3179 17279 3185
rect 17221 3176 17233 3179
rect 17184 3148 17233 3176
rect 17184 3136 17190 3148
rect 17221 3145 17233 3148
rect 17267 3145 17279 3179
rect 17221 3139 17279 3145
rect 18969 3179 19027 3185
rect 18969 3145 18981 3179
rect 19015 3176 19027 3179
rect 19334 3176 19340 3188
rect 19015 3148 19340 3176
rect 19015 3145 19027 3148
rect 18969 3139 19027 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 20441 3179 20499 3185
rect 20441 3145 20453 3179
rect 20487 3145 20499 3179
rect 20441 3139 20499 3145
rect 20456 3108 20484 3139
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 21085 3179 21143 3185
rect 21085 3176 21097 3179
rect 20772 3148 21097 3176
rect 20772 3136 20778 3148
rect 21085 3145 21097 3148
rect 21131 3145 21143 3179
rect 22738 3176 22744 3188
rect 22699 3148 22744 3176
rect 21085 3139 21143 3145
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 24210 3176 24216 3188
rect 24171 3148 24216 3176
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 24394 3136 24400 3188
rect 24452 3176 24458 3188
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 24452 3148 24685 3176
rect 24452 3136 24458 3148
rect 24673 3145 24685 3148
rect 24719 3145 24731 3179
rect 24673 3139 24731 3145
rect 24946 3136 24952 3188
rect 25004 3136 25010 3188
rect 25130 3176 25136 3188
rect 25056 3148 25136 3176
rect 20990 3108 20996 3120
rect 14752 3080 17724 3108
rect 13817 3071 13875 3077
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3009 12771 3043
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 12713 3003 12771 3009
rect 5644 2944 7328 2972
rect 11624 2944 12572 2972
rect 1636 2876 3464 2904
rect 1636 2864 1642 2876
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 3660 2876 5304 2904
rect 3660 2864 3666 2876
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 992 2808 4077 2836
rect 992 2796 998 2808
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4065 2799 4123 2805
rect 4982 2796 4988 2848
rect 5040 2836 5046 2848
rect 5169 2839 5227 2845
rect 5169 2836 5181 2839
rect 5040 2808 5181 2836
rect 5040 2796 5046 2808
rect 5169 2805 5181 2808
rect 5215 2805 5227 2839
rect 5276 2836 5304 2876
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 7193 2907 7251 2913
rect 7193 2904 7205 2907
rect 5684 2876 7205 2904
rect 5684 2864 5690 2876
rect 7193 2873 7205 2876
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 7300 2904 7328 2944
rect 8754 2904 8760 2916
rect 7300 2876 8760 2904
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 5276 2808 6469 2836
rect 5169 2799 5227 2805
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 6457 2799 6515 2805
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7300 2836 7328 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 10686 2904 10692 2916
rect 10551 2876 10692 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 10686 2864 10692 2876
rect 10744 2904 10750 2916
rect 11698 2904 11704 2916
rect 10744 2876 11704 2904
rect 10744 2864 10750 2876
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 12544 2913 12572 2944
rect 12529 2907 12587 2913
rect 12529 2873 12541 2907
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 6696 2808 7328 2836
rect 8665 2839 8723 2845
rect 6696 2796 6702 2808
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 9582 2836 9588 2848
rect 8711 2808 9588 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 12728 2836 12756 3003
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14516 3012 14565 3040
rect 14516 3000 14522 3012
rect 14553 3009 14565 3012
rect 14599 3040 14611 3043
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14599 3012 15209 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16390 3040 16396 3052
rect 16163 3012 16396 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17402 3040 17408 3052
rect 17363 3012 17408 3040
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 17696 3049 17724 3080
rect 18524 3080 20484 3108
rect 20548 3080 20996 3108
rect 18524 3049 18552 3080
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3040 18843 3043
rect 18966 3040 18972 3052
rect 18831 3012 18972 3040
rect 18831 3009 18843 3012
rect 18785 3003 18843 3009
rect 18966 3000 18972 3012
rect 19024 3040 19030 3052
rect 19426 3040 19432 3052
rect 19024 3012 19432 3040
rect 19024 3000 19030 3012
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 17310 2972 17316 2984
rect 13372 2944 17316 2972
rect 13372 2913 13400 2944
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 17604 2972 17632 3000
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 17604 2944 18613 2972
rect 18601 2941 18613 2944
rect 18647 2972 18659 2975
rect 19547 2972 19575 3003
rect 19702 3000 19708 3052
rect 19760 3040 19766 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19760 3012 19809 3040
rect 19760 3000 19766 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 20548 3040 20576 3080
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 24964 3108 24992 3136
rect 24872 3080 24992 3108
rect 20027 3012 20576 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 20680 3012 20725 3040
rect 20680 3000 20686 3012
rect 22646 3000 22652 3052
rect 22704 3040 22710 3052
rect 24872 3049 24900 3080
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 22704 3012 22937 3040
rect 22704 3000 22710 3012
rect 22925 3009 22937 3012
rect 22971 3040 22983 3043
rect 23385 3043 23443 3049
rect 23385 3040 23397 3043
rect 22971 3012 23397 3040
rect 22971 3009 22983 3012
rect 22925 3003 22983 3009
rect 23385 3009 23397 3012
rect 23431 3009 23443 3043
rect 23385 3003 23443 3009
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 24857 3043 24915 3049
rect 24857 3009 24869 3043
rect 24903 3009 24915 3043
rect 24857 3003 24915 3009
rect 24949 3043 25007 3049
rect 24949 3009 24961 3043
rect 24995 3040 25007 3043
rect 25056 3040 25084 3148
rect 25130 3136 25136 3148
rect 25188 3136 25194 3188
rect 26970 3176 26976 3188
rect 26931 3148 26976 3176
rect 26970 3136 26976 3148
rect 27028 3136 27034 3188
rect 28169 3179 28227 3185
rect 28169 3145 28181 3179
rect 28215 3176 28227 3179
rect 28534 3176 28540 3188
rect 28215 3148 28540 3176
rect 28215 3145 28227 3148
rect 28169 3139 28227 3145
rect 28534 3136 28540 3148
rect 28592 3176 28598 3188
rect 31110 3176 31116 3188
rect 28592 3148 31116 3176
rect 28592 3136 28598 3148
rect 31110 3136 31116 3148
rect 31168 3136 31174 3188
rect 31202 3136 31208 3188
rect 31260 3176 31266 3188
rect 33689 3179 33747 3185
rect 33689 3176 33701 3179
rect 31260 3148 33701 3176
rect 31260 3136 31266 3148
rect 33689 3145 33701 3148
rect 33735 3145 33747 3179
rect 33689 3139 33747 3145
rect 34517 3179 34575 3185
rect 34517 3145 34529 3179
rect 34563 3176 34575 3179
rect 35161 3179 35219 3185
rect 34563 3148 35112 3176
rect 34563 3145 34575 3148
rect 34517 3139 34575 3145
rect 28810 3108 28816 3120
rect 25148 3080 28816 3108
rect 25148 3049 25176 3080
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 29304 3111 29362 3117
rect 29304 3077 29316 3111
rect 29350 3108 29362 3111
rect 29454 3108 29460 3120
rect 29350 3080 29460 3108
rect 29350 3077 29362 3080
rect 29304 3071 29362 3077
rect 29454 3068 29460 3080
rect 29512 3068 29518 3120
rect 31573 3111 31631 3117
rect 31573 3077 31585 3111
rect 31619 3108 31631 3111
rect 34790 3108 34796 3120
rect 31619 3080 34796 3108
rect 31619 3077 31631 3080
rect 31573 3071 31631 3077
rect 24995 3012 25084 3040
rect 25133 3043 25191 3049
rect 24995 3009 25007 3012
rect 24949 3003 25007 3009
rect 25133 3009 25145 3043
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 20530 2972 20536 2984
rect 18647 2944 18828 2972
rect 19547 2944 20536 2972
rect 18647 2941 18659 2944
rect 18601 2935 18659 2941
rect 13357 2907 13415 2913
rect 13357 2873 13369 2907
rect 13403 2873 13415 2907
rect 13357 2867 13415 2873
rect 17218 2864 17224 2916
rect 17276 2904 17282 2916
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 17276 2876 17509 2904
rect 17276 2864 17282 2876
rect 17497 2873 17509 2876
rect 17543 2904 17555 2907
rect 18414 2904 18420 2916
rect 17543 2876 18420 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 18414 2864 18420 2876
rect 18472 2904 18478 2916
rect 18693 2907 18751 2913
rect 18693 2904 18705 2907
rect 18472 2876 18705 2904
rect 18472 2864 18478 2876
rect 18693 2873 18705 2876
rect 18739 2873 18751 2907
rect 18800 2904 18828 2944
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 24044 2972 24072 3003
rect 26694 3000 26700 3052
rect 26752 3040 26758 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26752 3012 27169 3040
rect 26752 3000 26758 3012
rect 27157 3009 27169 3012
rect 27203 3040 27215 3043
rect 27617 3043 27675 3049
rect 27617 3040 27629 3043
rect 27203 3012 27629 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 27617 3009 27629 3012
rect 27663 3009 27675 3043
rect 29546 3040 29552 3052
rect 29507 3012 29552 3040
rect 27617 3003 27675 3009
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 32401 3043 32459 3049
rect 32401 3009 32413 3043
rect 32447 3040 32459 3043
rect 32766 3040 32772 3052
rect 32447 3012 32772 3040
rect 32447 3009 32459 3012
rect 32401 3003 32459 3009
rect 32766 3000 32772 3012
rect 32824 3040 32830 3052
rect 33888 3049 33916 3080
rect 34790 3068 34796 3080
rect 34848 3068 34854 3120
rect 35084 3108 35112 3148
rect 35161 3145 35173 3179
rect 35207 3176 35219 3179
rect 38194 3176 38200 3188
rect 35207 3148 38200 3176
rect 35207 3145 35219 3148
rect 35161 3139 35219 3145
rect 38194 3136 38200 3148
rect 38252 3136 38258 3188
rect 37826 3108 37832 3120
rect 35084 3080 37832 3108
rect 37826 3068 37832 3080
rect 37884 3068 37890 3120
rect 33045 3043 33103 3049
rect 33045 3040 33057 3043
rect 32824 3012 33057 3040
rect 32824 3000 32830 3012
rect 33045 3009 33057 3012
rect 33091 3009 33103 3043
rect 33045 3003 33103 3009
rect 33873 3043 33931 3049
rect 33873 3009 33885 3043
rect 33919 3009 33931 3043
rect 33873 3003 33931 3009
rect 34333 3043 34391 3049
rect 34333 3009 34345 3043
rect 34379 3009 34391 3043
rect 34333 3003 34391 3009
rect 24670 2972 24676 2984
rect 24044 2944 24676 2972
rect 24670 2932 24676 2944
rect 24728 2972 24734 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 24728 2944 25697 2972
rect 24728 2932 24734 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 34348 2972 34376 3003
rect 34698 3000 34704 3052
rect 34756 3040 34762 3052
rect 34977 3043 35035 3049
rect 34977 3040 34989 3043
rect 34756 3012 34989 3040
rect 34756 3000 34762 3012
rect 34977 3009 34989 3012
rect 35023 3009 35035 3043
rect 35710 3040 35716 3052
rect 35671 3012 35716 3040
rect 34977 3003 35035 3009
rect 35710 3000 35716 3012
rect 35768 3000 35774 3052
rect 36170 3000 36176 3052
rect 36228 3040 36234 3052
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 36228 3012 36461 3040
rect 36228 3000 36234 3012
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 38105 3043 38163 3049
rect 38105 3040 38117 3043
rect 36449 3003 36507 3009
rect 37568 3012 38117 3040
rect 35066 2972 35072 2984
rect 25685 2935 25743 2941
rect 29564 2944 32904 2972
rect 34348 2944 35072 2972
rect 19613 2907 19671 2913
rect 19613 2904 19625 2907
rect 18800 2876 19625 2904
rect 18693 2867 18751 2873
rect 19613 2873 19625 2876
rect 19659 2873 19671 2907
rect 19613 2867 19671 2873
rect 19705 2907 19763 2913
rect 19705 2873 19717 2907
rect 19751 2904 19763 2907
rect 19978 2904 19984 2916
rect 19751 2876 19984 2904
rect 19751 2873 19763 2876
rect 19705 2867 19763 2873
rect 10468 2808 12756 2836
rect 10468 2796 10474 2808
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 15933 2839 15991 2845
rect 15933 2836 15945 2839
rect 15896 2808 15945 2836
rect 15896 2796 15902 2808
rect 15933 2805 15945 2808
rect 15979 2805 15991 2839
rect 15933 2799 15991 2805
rect 16761 2839 16819 2845
rect 16761 2805 16773 2839
rect 16807 2836 16819 2839
rect 18506 2836 18512 2848
rect 16807 2808 18512 2836
rect 16807 2805 16819 2808
rect 16761 2799 16819 2805
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 18708 2836 18736 2867
rect 19720 2836 19748 2867
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 21821 2907 21879 2913
rect 21821 2904 21833 2907
rect 20772 2876 21833 2904
rect 20772 2864 20778 2876
rect 21821 2873 21833 2876
rect 21867 2873 21879 2907
rect 21821 2867 21879 2873
rect 24118 2864 24124 2916
rect 24176 2864 24182 2916
rect 25041 2907 25099 2913
rect 25041 2873 25053 2907
rect 25087 2904 25099 2907
rect 25222 2904 25228 2916
rect 25087 2876 25228 2904
rect 25087 2873 25099 2876
rect 25041 2867 25099 2873
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 26602 2904 26608 2916
rect 25332 2876 26608 2904
rect 18708 2808 19748 2836
rect 24136 2836 24164 2864
rect 25332 2836 25360 2876
rect 26602 2864 26608 2876
rect 26660 2904 26666 2916
rect 26970 2904 26976 2916
rect 26660 2876 26976 2904
rect 26660 2864 26666 2876
rect 26970 2864 26976 2876
rect 27028 2864 27034 2916
rect 26234 2836 26240 2848
rect 24136 2808 25360 2836
rect 26195 2808 26240 2836
rect 26234 2796 26240 2808
rect 26292 2796 26298 2848
rect 27798 2796 27804 2848
rect 27856 2836 27862 2848
rect 29564 2836 29592 2944
rect 32876 2913 32904 2944
rect 35066 2932 35072 2944
rect 35124 2932 35130 2984
rect 35250 2932 35256 2984
rect 35308 2972 35314 2984
rect 37366 2972 37372 2984
rect 35308 2944 37372 2972
rect 35308 2932 35314 2944
rect 37366 2932 37372 2944
rect 37424 2932 37430 2984
rect 30377 2907 30435 2913
rect 30377 2873 30389 2907
rect 30423 2904 30435 2907
rect 32861 2907 32919 2913
rect 30423 2876 31754 2904
rect 30423 2873 30435 2876
rect 30377 2867 30435 2873
rect 27856 2808 29592 2836
rect 27856 2796 27862 2808
rect 30742 2796 30748 2848
rect 30800 2836 30806 2848
rect 30837 2839 30895 2845
rect 30837 2836 30849 2839
rect 30800 2808 30849 2836
rect 30800 2796 30806 2808
rect 30837 2805 30849 2808
rect 30883 2805 30895 2839
rect 31726 2836 31754 2876
rect 32861 2873 32873 2907
rect 32907 2873 32919 2907
rect 36633 2907 36691 2913
rect 32861 2867 32919 2873
rect 35820 2876 36584 2904
rect 35820 2836 35848 2876
rect 31726 2808 35848 2836
rect 35897 2839 35955 2845
rect 30837 2799 30895 2805
rect 35897 2805 35909 2839
rect 35943 2836 35955 2839
rect 36170 2836 36176 2848
rect 35943 2808 36176 2836
rect 35943 2805 35955 2808
rect 35897 2799 35955 2805
rect 36170 2796 36176 2808
rect 36228 2796 36234 2848
rect 36556 2836 36584 2876
rect 36633 2873 36645 2907
rect 36679 2904 36691 2907
rect 37458 2904 37464 2916
rect 36679 2876 37464 2904
rect 36679 2873 36691 2876
rect 36633 2867 36691 2873
rect 37458 2864 37464 2876
rect 37516 2864 37522 2916
rect 37568 2836 37596 3012
rect 38105 3009 38117 3012
rect 38151 3040 38163 3043
rect 39574 3040 39580 3052
rect 38151 3012 39580 3040
rect 38151 3009 38163 3012
rect 38105 3003 38163 3009
rect 39574 3000 39580 3012
rect 39632 3000 39638 3052
rect 37642 2864 37648 2916
rect 37700 2904 37706 2916
rect 37921 2907 37979 2913
rect 37921 2904 37933 2907
rect 37700 2876 37933 2904
rect 37700 2864 37706 2876
rect 37921 2873 37933 2876
rect 37967 2873 37979 2907
rect 37921 2867 37979 2873
rect 36556 2808 37596 2836
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 4062 2632 4068 2644
rect 3099 2604 4068 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 5592 2604 6469 2632
rect 5592 2592 5598 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10928 2604 10977 2632
rect 10928 2592 10934 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 14734 2632 14740 2644
rect 10965 2595 11023 2601
rect 11072 2604 14740 2632
rect 2866 2524 2872 2576
rect 2924 2564 2930 2576
rect 4798 2564 4804 2576
rect 2924 2536 4804 2564
rect 2924 2524 2930 2536
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 6886 2536 9812 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 6886 2496 6914 2536
rect 9674 2496 9680 2508
rect 1995 2468 6914 2496
rect 9416 2468 9680 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 290 2388 296 2440
rect 348 2428 354 2440
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 348 2400 2237 2428
rect 348 2388 354 2400
rect 2225 2397 2237 2400
rect 2271 2428 2283 2431
rect 2406 2428 2412 2440
rect 2271 2400 2412 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 2866 2428 2872 2440
rect 2823 2400 2872 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3804 2360 3832 2391
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3936 2400 4077 2428
rect 3936 2388 3942 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 5350 2428 5356 2440
rect 5311 2400 5356 2428
rect 4065 2391 4123 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 6638 2428 6644 2440
rect 6599 2400 6644 2428
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2428 7435 2431
rect 7742 2428 7748 2440
rect 7423 2400 7748 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8018 2388 8024 2440
rect 8076 2428 8082 2440
rect 9416 2437 9444 2468
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9784 2496 9812 2536
rect 10318 2524 10324 2576
rect 10376 2564 10382 2576
rect 10689 2567 10747 2573
rect 10689 2564 10701 2567
rect 10376 2536 10701 2564
rect 10376 2524 10382 2536
rect 10689 2533 10701 2536
rect 10735 2533 10747 2567
rect 10689 2527 10747 2533
rect 11072 2496 11100 2604
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 16853 2635 16911 2641
rect 16853 2601 16865 2635
rect 16899 2632 16911 2635
rect 18598 2632 18604 2644
rect 16899 2604 18604 2632
rect 16899 2601 16911 2604
rect 16853 2595 16911 2601
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 25774 2632 25780 2644
rect 20496 2604 25780 2632
rect 20496 2592 20502 2604
rect 25774 2592 25780 2604
rect 25832 2592 25838 2644
rect 26050 2592 26056 2644
rect 26108 2632 26114 2644
rect 26108 2604 34744 2632
rect 26108 2592 26114 2604
rect 20530 2524 20536 2576
rect 20588 2564 20594 2576
rect 20809 2567 20867 2573
rect 20809 2564 20821 2567
rect 20588 2536 20821 2564
rect 20588 2524 20594 2536
rect 20809 2533 20821 2536
rect 20855 2533 20867 2567
rect 20809 2527 20867 2533
rect 24118 2524 24124 2576
rect 24176 2564 24182 2576
rect 24176 2536 30328 2564
rect 24176 2524 24182 2536
rect 15746 2496 15752 2508
rect 9784 2468 11100 2496
rect 12544 2468 15752 2496
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 8076 2400 8125 2428
rect 8076 2388 8082 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 9640 2400 10517 2428
rect 9640 2388 9646 2400
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10686 2428 10692 2440
rect 10643 2400 10692 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10836 2400 10881 2428
rect 10836 2388 10842 2400
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 12544 2437 12572 2468
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 26234 2496 26240 2508
rect 16356 2468 21128 2496
rect 16356 2456 16362 2468
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11664 2400 11805 2428
rect 11664 2388 11670 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 13630 2428 13636 2440
rect 13587 2400 13636 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 15194 2428 15200 2440
rect 14415 2400 15200 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15378 2388 15384 2440
rect 15436 2428 15442 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15436 2400 15577 2428
rect 15436 2388 15442 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 16482 2428 16488 2440
rect 16163 2400 16488 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 16482 2388 16488 2400
rect 16540 2428 16546 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16540 2400 16681 2428
rect 16540 2388 16546 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17000 2400 17601 2428
rect 17000 2388 17006 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 17920 2400 18337 2428
rect 17920 2388 17926 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 18748 2400 19349 2428
rect 18748 2388 18754 2400
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 19337 2391 19395 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 20772 2400 21005 2428
rect 20772 2388 20778 2400
rect 20993 2397 21005 2400
rect 21039 2397 21051 2431
rect 21100 2428 21128 2468
rect 22112 2468 26240 2496
rect 22112 2437 22140 2468
rect 26234 2456 26240 2468
rect 26292 2456 26298 2508
rect 28905 2499 28963 2505
rect 28905 2496 28917 2499
rect 27724 2468 28917 2496
rect 27724 2440 27752 2468
rect 28905 2465 28917 2468
rect 28951 2465 28963 2499
rect 28905 2459 28963 2465
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21100 2400 22109 2428
rect 20993 2391 21051 2397
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2397 22615 2431
rect 23658 2428 23664 2440
rect 23619 2400 23664 2428
rect 22557 2391 22615 2397
rect 3970 2360 3976 2372
rect 3804 2332 3976 2360
rect 3970 2320 3976 2332
rect 4028 2320 4034 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 8444 2332 9873 2360
rect 8444 2320 8450 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 9861 2323 9919 2329
rect 20806 2320 20812 2372
rect 20864 2360 20870 2372
rect 22572 2360 22600 2391
rect 23658 2388 23664 2400
rect 23716 2388 23722 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 25685 2431 25743 2437
rect 25685 2397 25697 2431
rect 25731 2428 25743 2431
rect 25774 2428 25780 2440
rect 25731 2400 25780 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 20864 2332 22600 2360
rect 20864 2320 20870 2332
rect 22830 2320 22836 2372
rect 22888 2360 22894 2372
rect 24412 2360 24440 2391
rect 25774 2388 25780 2400
rect 25832 2388 25838 2440
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2397 26203 2431
rect 27706 2428 27712 2440
rect 27619 2400 27712 2428
rect 26145 2391 26203 2397
rect 22888 2332 24440 2360
rect 22888 2320 22894 2332
rect 24762 2320 24768 2372
rect 24820 2360 24826 2372
rect 26160 2360 26188 2391
rect 27706 2388 27712 2400
rect 27764 2388 27770 2440
rect 28169 2431 28227 2437
rect 28169 2397 28181 2431
rect 28215 2397 28227 2431
rect 28169 2391 28227 2397
rect 24820 2332 26188 2360
rect 24820 2320 24826 2332
rect 26970 2320 26976 2372
rect 27028 2360 27034 2372
rect 28184 2360 28212 2391
rect 29362 2388 29368 2440
rect 29420 2428 29426 2440
rect 30300 2437 30328 2536
rect 32122 2524 32128 2576
rect 32180 2564 32186 2576
rect 33045 2567 33103 2573
rect 33045 2564 33057 2567
rect 32180 2536 33057 2564
rect 32180 2524 32186 2536
rect 33045 2533 33057 2536
rect 33091 2533 33103 2567
rect 33045 2527 33103 2533
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29420 2400 29561 2428
rect 29420 2388 29426 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 30800 2400 31217 2428
rect 30800 2388 30806 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 32125 2431 32183 2437
rect 32125 2397 32137 2431
rect 32171 2428 32183 2431
rect 32214 2428 32220 2440
rect 32171 2400 32220 2428
rect 32171 2397 32183 2400
rect 32125 2391 32183 2397
rect 32214 2388 32220 2400
rect 32272 2388 32278 2440
rect 32858 2428 32864 2440
rect 32819 2400 32864 2428
rect 32858 2388 32864 2400
rect 32916 2388 32922 2440
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 34716 2437 34744 2604
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 37182 2496 37188 2508
rect 36964 2468 37188 2496
rect 36964 2456 36970 2468
rect 37182 2456 37188 2468
rect 37240 2496 37246 2508
rect 37277 2499 37335 2505
rect 37277 2496 37289 2499
rect 37240 2468 37289 2496
rect 37240 2456 37246 2468
rect 37277 2465 37289 2468
rect 37323 2465 37335 2499
rect 37277 2459 37335 2465
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33560 2400 33609 2428
rect 33560 2388 33566 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 34701 2431 34759 2437
rect 34701 2397 34713 2431
rect 34747 2397 34759 2431
rect 35618 2428 35624 2440
rect 35579 2400 35624 2428
rect 34701 2391 34759 2397
rect 35618 2388 35624 2400
rect 35676 2388 35682 2440
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 36136 2400 36461 2428
rect 36136 2388 36142 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 37550 2428 37556 2440
rect 37511 2400 37556 2428
rect 36449 2391 36507 2397
rect 37550 2388 37556 2400
rect 37608 2388 37614 2440
rect 27028 2332 28212 2360
rect 27028 2320 27034 2332
rect 28902 2320 28908 2372
rect 28960 2360 28966 2372
rect 28960 2332 31064 2360
rect 28960 2320 28966 2332
rect 2958 2252 2964 2304
rect 3016 2292 3022 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 3016 2264 5181 2292
rect 3016 2252 3022 2264
rect 5169 2261 5181 2264
rect 5215 2261 5227 2295
rect 5169 2255 5227 2261
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7193 2295 7251 2301
rect 7193 2292 7205 2295
rect 7064 2264 7205 2292
rect 7064 2252 7070 2264
rect 7193 2261 7205 2264
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9088 2264 9229 2292
rect 9088 2252 9094 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11609 2295 11667 2301
rect 11609 2292 11621 2295
rect 11112 2264 11621 2292
rect 11112 2252 11118 2264
rect 11609 2261 11621 2264
rect 11655 2261 11667 2295
rect 11609 2255 11667 2261
rect 11790 2252 11796 2304
rect 11848 2292 11854 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 11848 2264 12357 2292
rect 11848 2252 11854 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13228 2264 13369 2292
rect 13228 2252 13234 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 14185 2295 14243 2301
rect 14185 2292 14197 2295
rect 13872 2264 14197 2292
rect 13872 2252 13878 2264
rect 14185 2261 14197 2264
rect 14231 2261 14243 2295
rect 14185 2255 14243 2261
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 15252 2264 15393 2292
rect 15252 2252 15258 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17405 2295 17463 2301
rect 17405 2292 17417 2295
rect 17276 2264 17417 2292
rect 17276 2252 17282 2264
rect 17405 2261 17417 2264
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 18141 2295 18199 2301
rect 18141 2292 18153 2295
rect 17920 2264 18153 2292
rect 17920 2252 17926 2264
rect 18141 2261 18153 2264
rect 18187 2261 18199 2295
rect 18141 2255 18199 2261
rect 19242 2252 19248 2304
rect 19300 2292 19306 2304
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 19300 2264 19533 2292
rect 19300 2252 19306 2264
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19521 2255 19579 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21913 2295 21971 2301
rect 21913 2292 21925 2295
rect 21324 2264 21925 2292
rect 21324 2252 21330 2264
rect 21913 2261 21925 2264
rect 21959 2261 21971 2295
rect 21913 2255 21971 2261
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22060 2264 22753 2292
rect 22060 2252 22066 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23348 2264 23489 2292
rect 23348 2252 23354 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24084 2264 24593 2292
rect 24084 2252 24090 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 25314 2252 25320 2304
rect 25372 2292 25378 2304
rect 25501 2295 25559 2301
rect 25501 2292 25513 2295
rect 25372 2264 25513 2292
rect 25372 2252 25378 2264
rect 25501 2261 25513 2264
rect 25547 2261 25559 2295
rect 25501 2255 25559 2261
rect 26050 2252 26056 2304
rect 26108 2292 26114 2304
rect 26329 2295 26387 2301
rect 26329 2292 26341 2295
rect 26108 2264 26341 2292
rect 26108 2252 26114 2264
rect 26329 2261 26341 2264
rect 26375 2261 26387 2295
rect 26329 2255 26387 2261
rect 27338 2252 27344 2304
rect 27396 2292 27402 2304
rect 27525 2295 27583 2301
rect 27525 2292 27537 2295
rect 27396 2264 27537 2292
rect 27396 2252 27402 2264
rect 27525 2261 27537 2264
rect 27571 2261 27583 2295
rect 27525 2255 27583 2261
rect 28074 2252 28080 2304
rect 28132 2292 28138 2304
rect 28353 2295 28411 2301
rect 28353 2292 28365 2295
rect 28132 2264 28365 2292
rect 28132 2252 28138 2264
rect 28353 2261 28365 2264
rect 28399 2261 28411 2295
rect 28353 2255 28411 2261
rect 29454 2252 29460 2304
rect 29512 2292 29518 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 29512 2264 29745 2292
rect 29512 2252 29518 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 30098 2252 30104 2304
rect 30156 2292 30162 2304
rect 31036 2301 31064 2332
rect 30469 2295 30527 2301
rect 30469 2292 30481 2295
rect 30156 2264 30481 2292
rect 30156 2252 30162 2264
rect 30469 2261 30481 2264
rect 30515 2261 30527 2295
rect 30469 2255 30527 2261
rect 31021 2295 31079 2301
rect 31021 2261 31033 2295
rect 31067 2261 31079 2295
rect 31021 2255 31079 2261
rect 31478 2252 31484 2304
rect 31536 2292 31542 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 31536 2264 32321 2292
rect 31536 2252 31542 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 33560 2264 33793 2292
rect 33560 2252 33566 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 34204 2264 34897 2292
rect 34204 2252 34210 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 35526 2252 35532 2304
rect 35584 2292 35590 2304
rect 35805 2295 35863 2301
rect 35805 2292 35817 2295
rect 35584 2264 35817 2292
rect 35584 2252 35590 2264
rect 35805 2261 35817 2264
rect 35851 2261 35863 2295
rect 36630 2292 36636 2304
rect 36591 2264 36636 2292
rect 35805 2255 35863 2261
rect 36630 2252 36636 2264
rect 36688 2252 36694 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 20254 2048 20260 2100
rect 20312 2088 20318 2100
rect 23658 2088 23664 2100
rect 20312 2060 23664 2088
rect 20312 2048 20318 2060
rect 23658 2048 23664 2060
rect 23716 2048 23722 2100
rect 25866 2048 25872 2100
rect 25924 2088 25930 2100
rect 37550 2088 37556 2100
rect 25924 2060 37556 2088
rect 25924 2048 25930 2060
rect 37550 2048 37556 2060
rect 37608 2048 37614 2100
rect 20162 1980 20168 2032
rect 20220 2020 20226 2032
rect 27706 2020 27712 2032
rect 20220 1992 27712 2020
rect 20220 1980 20226 1992
rect 27706 1980 27712 1992
rect 27764 1980 27770 2032
rect 23658 1912 23664 1964
rect 23716 1952 23722 1964
rect 26142 1952 26148 1964
rect 23716 1924 26148 1952
rect 23716 1912 23722 1924
rect 26142 1912 26148 1924
rect 26200 1912 26206 1964
rect 27522 1912 27528 1964
rect 27580 1952 27586 1964
rect 32858 1952 32864 1964
rect 27580 1924 32864 1952
rect 27580 1912 27586 1924
rect 32858 1912 32864 1924
rect 32916 1912 32922 1964
rect 3970 212 3976 264
rect 4028 252 4034 264
rect 5718 252 5724 264
rect 4028 224 5724 252
rect 4028 212 4034 224
rect 5718 212 5724 224
rect 5776 212 5782 264
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2780 37408 2832 37460
rect 2872 37340 2924 37392
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 19432 37204 19484 37256
rect 35808 37247 35860 37256
rect 35808 37213 35817 37247
rect 35817 37213 35851 37247
rect 35851 37213 35860 37247
rect 35808 37204 35860 37213
rect 36084 37204 36136 37256
rect 35716 37136 35768 37188
rect 19984 37068 20036 37120
rect 35992 37111 36044 37120
rect 35992 37077 36001 37111
rect 36001 37077 36035 37111
rect 36035 37077 36044 37111
rect 35992 37068 36044 37077
rect 37280 37111 37332 37120
rect 37280 37077 37289 37111
rect 37289 37077 37323 37111
rect 37323 37077 37332 37111
rect 37280 37068 37332 37077
rect 38016 37111 38068 37120
rect 38016 37077 38025 37111
rect 38025 37077 38059 37111
rect 38059 37077 38068 37111
rect 38016 37068 38068 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 35808 36864 35860 36916
rect 38200 36864 38252 36916
rect 1492 36728 1544 36780
rect 38200 36728 38252 36780
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19432 36363 19484 36372
rect 19432 36329 19441 36363
rect 19441 36329 19475 36363
rect 19475 36329 19484 36363
rect 19432 36320 19484 36329
rect 38108 36320 38160 36372
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 18972 36116 19024 36168
rect 37372 36159 37424 36168
rect 37372 36125 37381 36159
rect 37381 36125 37415 36159
rect 37415 36125 37424 36159
rect 37372 36116 37424 36125
rect 32128 36048 32180 36100
rect 36912 35980 36964 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 37004 35640 37056 35692
rect 1400 35479 1452 35488
rect 1400 35445 1409 35479
rect 1409 35445 1443 35479
rect 1443 35445 1452 35479
rect 1400 35436 1452 35445
rect 38016 35479 38068 35488
rect 38016 35445 38025 35479
rect 38025 35445 38059 35479
rect 38059 35445 38068 35479
rect 38016 35436 38068 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 25780 34892 25832 34944
rect 38016 34935 38068 34944
rect 38016 34901 38025 34935
rect 38025 34901 38059 34935
rect 38059 34901 38068 34935
rect 38016 34892 38068 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1400 34459 1452 34468
rect 1400 34425 1409 34459
rect 1409 34425 1443 34459
rect 1443 34425 1452 34459
rect 1400 34416 1452 34425
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 38108 33983 38160 33992
rect 38108 33949 38117 33983
rect 38117 33949 38151 33983
rect 38151 33949 38160 33983
rect 38108 33940 38160 33949
rect 38292 33804 38344 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 37556 33464 37608 33516
rect 38016 33303 38068 33312
rect 38016 33269 38025 33303
rect 38025 33269 38059 33303
rect 38059 33269 38068 33303
rect 38016 33260 38068 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 28356 32852 28408 32904
rect 38016 32759 38068 32768
rect 38016 32725 38025 32759
rect 38025 32725 38059 32759
rect 38059 32725 38068 32759
rect 38016 32716 38068 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 38108 32419 38160 32428
rect 38108 32385 38117 32419
rect 38117 32385 38151 32419
rect 38151 32385 38160 32419
rect 38108 32376 38160 32385
rect 37924 32215 37976 32224
rect 37924 32181 37933 32215
rect 37933 32181 37967 32215
rect 37967 32181 37976 32215
rect 37924 32172 37976 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 35992 31764 36044 31816
rect 38200 31764 38252 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1492 31288 1544 31340
rect 37832 31331 37884 31340
rect 37832 31297 37841 31331
rect 37841 31297 37875 31331
rect 37875 31297 37884 31331
rect 37832 31288 37884 31297
rect 2596 31084 2648 31136
rect 38016 31127 38068 31136
rect 38016 31093 38025 31127
rect 38025 31093 38059 31127
rect 38059 31093 38068 31127
rect 38016 31084 38068 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 2504 30540 2556 30592
rect 28448 30540 28500 30592
rect 38016 30583 38068 30592
rect 38016 30549 38025 30583
rect 38025 30549 38059 30583
rect 38059 30549 38068 30583
rect 38016 30540 38068 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 38108 30243 38160 30252
rect 38108 30209 38117 30243
rect 38117 30209 38151 30243
rect 38151 30209 38160 30243
rect 38108 30200 38160 30209
rect 1400 30039 1452 30048
rect 1400 30005 1409 30039
rect 1409 30005 1443 30039
rect 1443 30005 1452 30039
rect 1400 29996 1452 30005
rect 37740 29996 37792 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 1584 29495 1636 29504
rect 1584 29461 1593 29495
rect 1593 29461 1627 29495
rect 1627 29461 1636 29495
rect 1584 29452 1636 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1584 29180 1636 29232
rect 2504 29155 2556 29164
rect 2504 29121 2513 29155
rect 2513 29121 2547 29155
rect 2547 29121 2556 29155
rect 2504 29112 2556 29121
rect 38200 29112 38252 29164
rect 2596 29087 2648 29096
rect 2596 29053 2605 29087
rect 2605 29053 2639 29087
rect 2639 29053 2648 29087
rect 2596 29044 2648 29053
rect 1400 29019 1452 29028
rect 1400 28985 1409 29019
rect 1409 28985 1443 29019
rect 1443 28985 1452 29019
rect 1400 28976 1452 28985
rect 3516 28976 3568 29028
rect 38016 29019 38068 29028
rect 38016 28985 38025 29019
rect 38025 28985 38059 29019
rect 38059 28985 38068 29019
rect 38016 28976 38068 28985
rect 1584 28908 1636 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 27620 28364 27672 28416
rect 38016 28407 38068 28416
rect 38016 28373 38025 28407
rect 38025 28373 38059 28407
rect 38059 28373 38068 28407
rect 38016 28364 38068 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1584 28203 1636 28212
rect 1584 28169 1593 28203
rect 1593 28169 1627 28203
rect 1627 28169 1636 28203
rect 1584 28160 1636 28169
rect 32128 28203 32180 28212
rect 32128 28169 32137 28203
rect 32137 28169 32171 28203
rect 32171 28169 32180 28203
rect 32128 28160 32180 28169
rect 32864 28160 32916 28212
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 33232 28067 33284 28076
rect 33232 28033 33250 28067
rect 33250 28033 33284 28067
rect 33232 28024 33284 28033
rect 38108 28067 38160 28076
rect 38108 28033 38117 28067
rect 38117 28033 38151 28067
rect 38151 28033 38160 28067
rect 38108 28024 38160 28033
rect 33508 27999 33560 28008
rect 33508 27965 33517 27999
rect 33517 27965 33551 27999
rect 33551 27965 33560 27999
rect 33508 27956 33560 27965
rect 37648 27820 37700 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 25780 27591 25832 27600
rect 25780 27557 25789 27591
rect 25789 27557 25823 27591
rect 25823 27557 25832 27591
rect 25780 27548 25832 27557
rect 33232 27548 33284 27600
rect 36084 27591 36136 27600
rect 36084 27557 36093 27591
rect 36093 27557 36127 27591
rect 36127 27557 36136 27591
rect 36084 27548 36136 27557
rect 32036 27480 32088 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 22928 27412 22980 27464
rect 26976 27412 27028 27464
rect 22376 27344 22428 27396
rect 24860 27344 24912 27396
rect 30564 27344 30616 27396
rect 33508 27412 33560 27464
rect 35348 27412 35400 27464
rect 37280 27412 37332 27464
rect 34152 27344 34204 27396
rect 23664 27319 23716 27328
rect 23664 27285 23673 27319
rect 23673 27285 23707 27319
rect 23707 27285 23716 27319
rect 23664 27276 23716 27285
rect 32956 27276 33008 27328
rect 33600 27319 33652 27328
rect 33600 27285 33609 27319
rect 33609 27285 33643 27319
rect 33643 27285 33652 27319
rect 33600 27276 33652 27285
rect 33692 27276 33744 27328
rect 37464 27344 37516 27396
rect 37188 27276 37240 27328
rect 38016 27319 38068 27328
rect 38016 27285 38025 27319
rect 38025 27285 38059 27319
rect 38059 27285 38068 27319
rect 38016 27276 38068 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 24860 27115 24912 27124
rect 24860 27081 24869 27115
rect 24869 27081 24903 27115
rect 24903 27081 24912 27115
rect 24860 27072 24912 27081
rect 28356 27115 28408 27124
rect 28356 27081 28365 27115
rect 28365 27081 28399 27115
rect 28399 27081 28408 27115
rect 28356 27072 28408 27081
rect 30564 27115 30616 27124
rect 30564 27081 30573 27115
rect 30573 27081 30607 27115
rect 30607 27081 30616 27115
rect 30564 27072 30616 27081
rect 27528 27004 27580 27056
rect 31300 27072 31352 27124
rect 33600 27072 33652 27124
rect 34152 27115 34204 27124
rect 34152 27081 34161 27115
rect 34161 27081 34195 27115
rect 34195 27081 34204 27115
rect 34152 27072 34204 27081
rect 36636 27072 36688 27124
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 22284 26979 22336 26988
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 22928 26979 22980 26988
rect 22928 26945 22937 26979
rect 22937 26945 22971 26979
rect 22971 26945 22980 26979
rect 22928 26936 22980 26945
rect 23480 26936 23532 26988
rect 26976 26979 27028 26988
rect 26976 26945 26985 26979
rect 26985 26945 27019 26979
rect 27019 26945 27028 26979
rect 26976 26936 27028 26945
rect 27068 26936 27120 26988
rect 30840 26936 30892 26988
rect 33508 27004 33560 27056
rect 35992 27004 36044 27056
rect 38384 27004 38436 27056
rect 32220 26936 32272 26988
rect 34152 26936 34204 26988
rect 37188 26936 37240 26988
rect 31392 26843 31444 26852
rect 2872 26732 2924 26784
rect 23572 26732 23624 26784
rect 31392 26809 31401 26843
rect 31401 26809 31435 26843
rect 31435 26809 31444 26843
rect 31392 26800 31444 26809
rect 31760 26732 31812 26784
rect 33508 26868 33560 26920
rect 37004 26868 37056 26920
rect 37372 26868 37424 26920
rect 33508 26775 33560 26784
rect 33508 26741 33517 26775
rect 33517 26741 33551 26775
rect 33551 26741 33560 26775
rect 33508 26732 33560 26741
rect 37096 26732 37148 26784
rect 37372 26732 37424 26784
rect 38384 26732 38436 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 22376 26571 22428 26580
rect 22376 26537 22385 26571
rect 22385 26537 22419 26571
rect 22419 26537 22428 26571
rect 22376 26528 22428 26537
rect 23480 26571 23532 26580
rect 23480 26537 23489 26571
rect 23489 26537 23523 26571
rect 23523 26537 23532 26571
rect 23480 26528 23532 26537
rect 27068 26528 27120 26580
rect 30840 26571 30892 26580
rect 23388 26503 23440 26512
rect 23388 26469 23397 26503
rect 23397 26469 23431 26503
rect 23431 26469 23440 26503
rect 23388 26460 23440 26469
rect 24676 26460 24728 26512
rect 30288 26503 30340 26512
rect 30288 26469 30297 26503
rect 30297 26469 30331 26503
rect 30331 26469 30340 26503
rect 30288 26460 30340 26469
rect 30840 26537 30849 26571
rect 30849 26537 30883 26571
rect 30883 26537 30892 26571
rect 30840 26528 30892 26537
rect 32220 26528 32272 26580
rect 30932 26503 30984 26512
rect 30932 26469 30941 26503
rect 30941 26469 30975 26503
rect 30975 26469 30984 26503
rect 30932 26460 30984 26469
rect 34152 26528 34204 26580
rect 35992 26528 36044 26580
rect 36268 26571 36320 26580
rect 36268 26537 36277 26571
rect 36277 26537 36311 26571
rect 36311 26537 36320 26571
rect 36268 26528 36320 26537
rect 37372 26528 37424 26580
rect 37096 26460 37148 26512
rect 38016 26503 38068 26512
rect 32588 26435 32640 26444
rect 22652 26324 22704 26376
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 27528 26324 27580 26376
rect 32588 26401 32597 26435
rect 32597 26401 32631 26435
rect 32631 26401 32640 26435
rect 32588 26392 32640 26401
rect 36084 26392 36136 26444
rect 36544 26392 36596 26444
rect 31760 26367 31812 26376
rect 2228 26299 2280 26308
rect 2228 26265 2237 26299
rect 2237 26265 2271 26299
rect 2271 26265 2280 26299
rect 2228 26256 2280 26265
rect 22928 26256 22980 26308
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 23756 26188 23808 26240
rect 24676 26188 24728 26240
rect 27620 26256 27672 26308
rect 27896 26256 27948 26308
rect 31300 26299 31352 26308
rect 31300 26265 31309 26299
rect 31309 26265 31343 26299
rect 31343 26265 31352 26299
rect 31300 26256 31352 26265
rect 31760 26333 31769 26367
rect 31769 26333 31803 26367
rect 31803 26333 31812 26367
rect 31760 26324 31812 26333
rect 33600 26367 33652 26376
rect 33600 26333 33609 26367
rect 33609 26333 33643 26367
rect 33643 26333 33652 26367
rect 33600 26324 33652 26333
rect 36268 26324 36320 26376
rect 37004 26367 37056 26376
rect 37004 26333 37013 26367
rect 37013 26333 37047 26367
rect 37047 26333 37056 26367
rect 37004 26324 37056 26333
rect 38016 26469 38025 26503
rect 38025 26469 38059 26503
rect 38059 26469 38068 26503
rect 38016 26460 38068 26469
rect 32036 26256 32088 26308
rect 33140 26256 33192 26308
rect 32588 26188 32640 26240
rect 37464 26324 37516 26376
rect 38292 26324 38344 26376
rect 36728 26231 36780 26240
rect 36728 26197 36737 26231
rect 36737 26197 36771 26231
rect 36771 26197 36780 26231
rect 36728 26188 36780 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 22284 25984 22336 26036
rect 26240 25984 26292 26036
rect 27896 26027 27948 26036
rect 27896 25993 27905 26027
rect 27905 25993 27939 26027
rect 27939 25993 27948 26027
rect 27896 25984 27948 25993
rect 30932 25984 30984 26036
rect 31392 25984 31444 26036
rect 33508 25984 33560 26036
rect 32956 25916 33008 25968
rect 37556 25984 37608 26036
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 21180 25848 21232 25900
rect 28080 25891 28132 25900
rect 22468 25780 22520 25832
rect 22928 25780 22980 25832
rect 23664 25780 23716 25832
rect 26240 25780 26292 25832
rect 27436 25823 27488 25832
rect 27436 25789 27445 25823
rect 27445 25789 27479 25823
rect 27479 25789 27488 25823
rect 27436 25780 27488 25789
rect 23020 25712 23072 25764
rect 27068 25755 27120 25764
rect 27068 25721 27077 25755
rect 27077 25721 27111 25755
rect 27111 25721 27120 25755
rect 27068 25712 27120 25721
rect 28080 25857 28089 25891
rect 28089 25857 28123 25891
rect 28123 25857 28132 25891
rect 28080 25848 28132 25857
rect 30380 25891 30432 25900
rect 30380 25857 30389 25891
rect 30389 25857 30423 25891
rect 30423 25857 30432 25891
rect 30380 25848 30432 25857
rect 32772 25848 32824 25900
rect 36268 25891 36320 25900
rect 36268 25857 36272 25891
rect 36272 25857 36306 25891
rect 36306 25857 36320 25891
rect 36268 25848 36320 25857
rect 32588 25780 32640 25832
rect 32864 25780 32916 25832
rect 36544 25848 36596 25900
rect 36912 25916 36964 25968
rect 37832 25916 37884 25968
rect 38200 25916 38252 25968
rect 33140 25712 33192 25764
rect 36268 25712 36320 25764
rect 37096 25848 37148 25900
rect 37556 25891 37608 25900
rect 37556 25857 37560 25891
rect 37560 25857 37594 25891
rect 37594 25857 37608 25891
rect 37556 25848 37608 25857
rect 37924 25891 37976 25900
rect 37004 25780 37056 25832
rect 37924 25857 37932 25891
rect 37932 25857 37966 25891
rect 37966 25857 37976 25891
rect 37924 25848 37976 25857
rect 21180 25687 21232 25696
rect 21180 25653 21189 25687
rect 21189 25653 21223 25687
rect 21223 25653 21232 25687
rect 21180 25644 21232 25653
rect 22560 25644 22612 25696
rect 24400 25687 24452 25696
rect 24400 25653 24409 25687
rect 24409 25653 24443 25687
rect 24443 25653 24452 25687
rect 24400 25644 24452 25653
rect 32588 25644 32640 25696
rect 36084 25687 36136 25696
rect 36084 25653 36093 25687
rect 36093 25653 36127 25687
rect 36127 25653 36136 25687
rect 36084 25644 36136 25653
rect 37372 25687 37424 25696
rect 37372 25653 37381 25687
rect 37381 25653 37415 25687
rect 37415 25653 37424 25687
rect 37372 25644 37424 25653
rect 37556 25712 37608 25764
rect 37832 25712 37884 25764
rect 38292 25712 38344 25764
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 22652 25483 22704 25492
rect 22652 25449 22661 25483
rect 22661 25449 22695 25483
rect 22695 25449 22704 25483
rect 22652 25440 22704 25449
rect 23020 25440 23072 25492
rect 23388 25440 23440 25492
rect 25780 25440 25832 25492
rect 28448 25483 28500 25492
rect 28448 25449 28457 25483
rect 28457 25449 28491 25483
rect 28491 25449 28500 25483
rect 28448 25440 28500 25449
rect 30288 25440 30340 25492
rect 36176 25440 36228 25492
rect 2780 25372 2832 25424
rect 22560 25415 22612 25424
rect 22560 25381 22569 25415
rect 22569 25381 22603 25415
rect 22603 25381 22612 25415
rect 22560 25372 22612 25381
rect 23572 25347 23624 25356
rect 23572 25313 23581 25347
rect 23581 25313 23615 25347
rect 23615 25313 23624 25347
rect 23572 25304 23624 25313
rect 26240 25304 26292 25356
rect 32588 25304 32640 25356
rect 35348 25304 35400 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 24492 25236 24544 25288
rect 25780 25236 25832 25288
rect 22468 25168 22520 25220
rect 2688 25143 2740 25152
rect 2688 25109 2697 25143
rect 2697 25109 2731 25143
rect 2731 25109 2740 25143
rect 2688 25100 2740 25109
rect 21640 25143 21692 25152
rect 21640 25109 21649 25143
rect 21649 25109 21683 25143
rect 21683 25109 21692 25143
rect 24676 25168 24728 25220
rect 21640 25100 21692 25109
rect 24400 25100 24452 25152
rect 25872 25100 25924 25152
rect 26240 25143 26292 25152
rect 26240 25109 26249 25143
rect 26249 25109 26283 25143
rect 26283 25109 26292 25143
rect 32864 25236 32916 25288
rect 37280 25372 37332 25424
rect 37188 25236 37240 25288
rect 37464 25279 37516 25288
rect 37464 25245 37474 25279
rect 37474 25245 37508 25279
rect 37508 25245 37516 25279
rect 37464 25236 37516 25245
rect 37832 25279 37884 25288
rect 37832 25245 37846 25279
rect 37846 25245 37880 25279
rect 37880 25245 37884 25279
rect 37832 25236 37884 25245
rect 27344 25211 27396 25220
rect 27344 25177 27356 25211
rect 27356 25177 27396 25211
rect 27344 25168 27396 25177
rect 27528 25168 27580 25220
rect 35532 25168 35584 25220
rect 35900 25168 35952 25220
rect 36544 25168 36596 25220
rect 37004 25168 37056 25220
rect 26240 25100 26292 25109
rect 30472 25100 30524 25152
rect 31300 25100 31352 25152
rect 32772 25143 32824 25152
rect 32772 25109 32781 25143
rect 32781 25109 32815 25143
rect 32815 25109 32824 25143
rect 32772 25100 32824 25109
rect 37280 25100 37332 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 27068 24896 27120 24948
rect 27712 24896 27764 24948
rect 28264 24896 28316 24948
rect 25872 24828 25924 24880
rect 32772 24828 32824 24880
rect 1860 24803 1912 24812
rect 1860 24769 1869 24803
rect 1869 24769 1903 24803
rect 1903 24769 1912 24803
rect 1860 24760 1912 24769
rect 23848 24760 23900 24812
rect 26240 24803 26292 24812
rect 26240 24769 26249 24803
rect 26249 24769 26283 24803
rect 26283 24769 26292 24803
rect 26240 24760 26292 24769
rect 23664 24692 23716 24744
rect 24860 24692 24912 24744
rect 28356 24760 28408 24812
rect 30472 24760 30524 24812
rect 35348 24803 35400 24812
rect 35348 24769 35357 24803
rect 35357 24769 35391 24803
rect 35391 24769 35400 24803
rect 35348 24760 35400 24769
rect 35992 24760 36044 24812
rect 37556 24760 37608 24812
rect 28264 24735 28316 24744
rect 21640 24624 21692 24676
rect 23020 24624 23072 24676
rect 26332 24624 26384 24676
rect 27160 24624 27212 24676
rect 28264 24701 28273 24735
rect 28273 24701 28307 24735
rect 28307 24701 28316 24735
rect 28264 24692 28316 24701
rect 30380 24692 30432 24744
rect 37464 24692 37516 24744
rect 38108 24692 38160 24744
rect 38016 24667 38068 24676
rect 38016 24633 38025 24667
rect 38025 24633 38059 24667
rect 38059 24633 38068 24667
rect 38016 24624 38068 24633
rect 22468 24556 22520 24608
rect 22836 24556 22888 24608
rect 23848 24556 23900 24608
rect 27344 24556 27396 24608
rect 32588 24556 32640 24608
rect 37188 24556 37240 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1492 24395 1544 24404
rect 1492 24361 1501 24395
rect 1501 24361 1535 24395
rect 1535 24361 1544 24395
rect 1492 24352 1544 24361
rect 24492 24395 24544 24404
rect 24492 24361 24501 24395
rect 24501 24361 24535 24395
rect 24535 24361 24544 24395
rect 24492 24352 24544 24361
rect 28080 24352 28132 24404
rect 35532 24395 35584 24404
rect 35532 24361 35541 24395
rect 35541 24361 35575 24395
rect 35575 24361 35584 24395
rect 35532 24352 35584 24361
rect 35992 24395 36044 24404
rect 35992 24361 36001 24395
rect 36001 24361 36035 24395
rect 36035 24361 36044 24395
rect 35992 24352 36044 24361
rect 36268 24352 36320 24404
rect 37188 24352 37240 24404
rect 2228 24284 2280 24336
rect 23572 24284 23624 24336
rect 27068 24327 27120 24336
rect 27068 24293 27077 24327
rect 27077 24293 27111 24327
rect 27111 24293 27120 24327
rect 27068 24284 27120 24293
rect 27896 24327 27948 24336
rect 27896 24293 27905 24327
rect 27905 24293 27939 24327
rect 27939 24293 27948 24327
rect 27896 24284 27948 24293
rect 28448 24284 28500 24336
rect 2688 24216 2740 24268
rect 22652 24216 22704 24268
rect 22836 24259 22888 24268
rect 22836 24225 22845 24259
rect 22845 24225 22879 24259
rect 22879 24225 22888 24259
rect 22836 24216 22888 24225
rect 27436 24216 27488 24268
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 21824 24080 21876 24132
rect 37280 24284 37332 24336
rect 37832 24284 37884 24336
rect 38292 24284 38344 24336
rect 23020 24080 23072 24132
rect 23848 24123 23900 24132
rect 2412 24012 2464 24064
rect 22560 24012 22612 24064
rect 23480 24055 23532 24064
rect 23480 24021 23489 24055
rect 23489 24021 23523 24055
rect 23523 24021 23532 24055
rect 23480 24012 23532 24021
rect 23848 24089 23857 24123
rect 23857 24089 23891 24123
rect 23891 24089 23900 24123
rect 23848 24080 23900 24089
rect 28908 24080 28960 24132
rect 36728 24216 36780 24268
rect 34520 24148 34572 24200
rect 36176 24191 36228 24200
rect 36176 24157 36185 24191
rect 36185 24157 36219 24191
rect 36219 24157 36228 24191
rect 36176 24148 36228 24157
rect 37372 24148 37424 24200
rect 24492 24012 24544 24064
rect 27160 24012 27212 24064
rect 28632 24012 28684 24064
rect 31392 24012 31444 24064
rect 38016 24055 38068 24064
rect 38016 24021 38025 24055
rect 38025 24021 38059 24055
rect 38059 24021 38068 24055
rect 38016 24012 38068 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 22652 23851 22704 23860
rect 22652 23817 22661 23851
rect 22661 23817 22695 23851
rect 22695 23817 22704 23851
rect 22652 23808 22704 23817
rect 24952 23808 25004 23860
rect 27896 23808 27948 23860
rect 29000 23808 29052 23860
rect 31392 23808 31444 23860
rect 36084 23740 36136 23792
rect 2412 23715 2464 23724
rect 2412 23681 2421 23715
rect 2421 23681 2455 23715
rect 2455 23681 2464 23715
rect 2412 23672 2464 23681
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2872 23715 2924 23724
rect 2504 23672 2556 23681
rect 2872 23681 2881 23715
rect 2881 23681 2915 23715
rect 2915 23681 2924 23715
rect 2872 23672 2924 23681
rect 22100 23672 22152 23724
rect 21640 23604 21692 23656
rect 23572 23672 23624 23724
rect 23848 23672 23900 23724
rect 25044 23672 25096 23724
rect 22652 23604 22704 23656
rect 16948 23536 17000 23588
rect 34152 23672 34204 23724
rect 38108 23715 38160 23724
rect 38108 23681 38117 23715
rect 38117 23681 38151 23715
rect 38151 23681 38160 23715
rect 38108 23672 38160 23681
rect 27344 23536 27396 23588
rect 28816 23604 28868 23656
rect 27620 23536 27672 23588
rect 1492 23511 1544 23520
rect 1492 23477 1501 23511
rect 1501 23477 1535 23511
rect 1535 23477 1544 23511
rect 1492 23468 1544 23477
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 2780 23468 2832 23477
rect 3332 23468 3384 23520
rect 3608 23511 3660 23520
rect 3608 23477 3617 23511
rect 3617 23477 3651 23511
rect 3651 23477 3660 23511
rect 3608 23468 3660 23477
rect 26884 23468 26936 23520
rect 28724 23511 28776 23520
rect 28724 23477 28733 23511
rect 28733 23477 28767 23511
rect 28767 23477 28776 23511
rect 28724 23468 28776 23477
rect 37832 23468 37884 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 24860 23264 24912 23316
rect 26240 23264 26292 23316
rect 29460 23264 29512 23316
rect 33692 23264 33744 23316
rect 36176 23264 36228 23316
rect 24400 23196 24452 23248
rect 26884 23239 26936 23248
rect 26884 23205 26893 23239
rect 26893 23205 26927 23239
rect 26927 23205 26936 23239
rect 26884 23196 26936 23205
rect 35072 23239 35124 23248
rect 35072 23205 35081 23239
rect 35081 23205 35115 23239
rect 35115 23205 35124 23239
rect 35072 23196 35124 23205
rect 23480 23128 23532 23180
rect 26240 23128 26292 23180
rect 27436 23128 27488 23180
rect 27620 23171 27672 23180
rect 27620 23137 27629 23171
rect 27629 23137 27663 23171
rect 27663 23137 27672 23171
rect 27620 23128 27672 23137
rect 22928 23103 22980 23112
rect 22928 23069 22937 23103
rect 22937 23069 22971 23103
rect 22971 23069 22980 23103
rect 22928 23060 22980 23069
rect 1860 23035 1912 23044
rect 1860 23001 1869 23035
rect 1869 23001 1903 23035
rect 1903 23001 1912 23035
rect 1860 22992 1912 23001
rect 3608 22992 3660 23044
rect 22652 23035 22704 23044
rect 22652 23001 22661 23035
rect 22661 23001 22695 23035
rect 22695 23001 22704 23035
rect 22652 22992 22704 23001
rect 23204 22992 23256 23044
rect 28908 23060 28960 23112
rect 31392 23103 31444 23112
rect 31392 23069 31401 23103
rect 31401 23069 31435 23103
rect 31435 23069 31444 23103
rect 31392 23060 31444 23069
rect 37924 23060 37976 23112
rect 27252 22992 27304 23044
rect 31484 22992 31536 23044
rect 34612 22992 34664 23044
rect 25044 22924 25096 22976
rect 26792 22924 26844 22976
rect 27620 22924 27672 22976
rect 32772 22967 32824 22976
rect 32772 22933 32781 22967
rect 32781 22933 32815 22967
rect 32815 22933 32824 22967
rect 32772 22924 32824 22933
rect 37556 22924 37608 22976
rect 38016 22967 38068 22976
rect 38016 22933 38025 22967
rect 38025 22933 38059 22967
rect 38059 22933 38068 22967
rect 38016 22924 38068 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2504 22720 2556 22772
rect 24952 22763 25004 22772
rect 24952 22729 24961 22763
rect 24961 22729 24995 22763
rect 24995 22729 25004 22763
rect 24952 22720 25004 22729
rect 27252 22720 27304 22772
rect 27620 22720 27672 22772
rect 29460 22763 29512 22772
rect 29460 22729 29469 22763
rect 29469 22729 29503 22763
rect 29503 22729 29512 22763
rect 29460 22720 29512 22729
rect 31484 22763 31536 22772
rect 31484 22729 31493 22763
rect 31493 22729 31527 22763
rect 31527 22729 31536 22763
rect 31484 22720 31536 22729
rect 34520 22720 34572 22772
rect 37464 22720 37516 22772
rect 38384 22720 38436 22772
rect 24860 22652 24912 22704
rect 2136 22627 2188 22636
rect 2136 22593 2145 22627
rect 2145 22593 2179 22627
rect 2179 22593 2188 22627
rect 2136 22584 2188 22593
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 28264 22652 28316 22704
rect 25228 22516 25280 22568
rect 26792 22516 26844 22568
rect 33968 22652 34020 22704
rect 37372 22652 37424 22704
rect 28908 22584 28960 22636
rect 27344 22516 27396 22568
rect 27620 22516 27672 22568
rect 28724 22559 28776 22568
rect 1492 22423 1544 22432
rect 1492 22389 1501 22423
rect 1501 22389 1535 22423
rect 1535 22389 1544 22423
rect 1492 22380 1544 22389
rect 3424 22423 3476 22432
rect 3424 22389 3433 22423
rect 3433 22389 3467 22423
rect 3467 22389 3476 22423
rect 3424 22380 3476 22389
rect 22100 22380 22152 22432
rect 24032 22423 24084 22432
rect 24032 22389 24041 22423
rect 24041 22389 24075 22423
rect 24075 22389 24084 22423
rect 24032 22380 24084 22389
rect 24308 22380 24360 22432
rect 25320 22380 25372 22432
rect 27068 22448 27120 22500
rect 28724 22525 28733 22559
rect 28733 22525 28767 22559
rect 28767 22525 28776 22559
rect 28724 22516 28776 22525
rect 34520 22584 34572 22636
rect 35808 22627 35860 22636
rect 35808 22593 35817 22627
rect 35817 22593 35851 22627
rect 35851 22593 35860 22627
rect 35808 22584 35860 22593
rect 37464 22627 37516 22636
rect 37464 22593 37468 22627
rect 37468 22593 37502 22627
rect 37502 22593 37516 22627
rect 37464 22584 37516 22593
rect 32496 22516 32548 22568
rect 34612 22516 34664 22568
rect 34796 22559 34848 22568
rect 34796 22525 34805 22559
rect 34805 22525 34839 22559
rect 34839 22525 34848 22559
rect 34796 22516 34848 22525
rect 37188 22516 37240 22568
rect 37740 22627 37792 22636
rect 37740 22593 37785 22627
rect 37785 22593 37792 22627
rect 37740 22584 37792 22593
rect 38108 22584 38160 22636
rect 38200 22516 38252 22568
rect 32220 22491 32272 22500
rect 32220 22457 32229 22491
rect 32229 22457 32263 22491
rect 32263 22457 32272 22491
rect 32220 22448 32272 22457
rect 34060 22491 34112 22500
rect 34060 22457 34069 22491
rect 34069 22457 34103 22491
rect 34103 22457 34112 22491
rect 34060 22448 34112 22457
rect 35072 22448 35124 22500
rect 27804 22423 27856 22432
rect 27804 22389 27813 22423
rect 27813 22389 27847 22423
rect 27847 22389 27856 22423
rect 27804 22380 27856 22389
rect 31024 22380 31076 22432
rect 36084 22380 36136 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 28908 22176 28960 22228
rect 34520 22176 34572 22228
rect 35808 22176 35860 22228
rect 35992 22176 36044 22228
rect 37188 22219 37240 22228
rect 37188 22185 37197 22219
rect 37197 22185 37231 22219
rect 37231 22185 37240 22219
rect 37188 22176 37240 22185
rect 26332 22108 26384 22160
rect 27804 22108 27856 22160
rect 34704 22108 34756 22160
rect 17224 22040 17276 22092
rect 22652 22040 22704 22092
rect 22560 22015 22612 22024
rect 22560 21981 22569 22015
rect 22569 21981 22603 22015
rect 22603 21981 22612 22015
rect 22560 21972 22612 21981
rect 23296 22040 23348 22092
rect 26148 22040 26200 22092
rect 27436 22040 27488 22092
rect 28080 22040 28132 22092
rect 28264 22083 28316 22092
rect 28264 22049 28273 22083
rect 28273 22049 28307 22083
rect 28307 22049 28316 22083
rect 28264 22040 28316 22049
rect 28448 22040 28500 22092
rect 28908 22040 28960 22092
rect 24032 21972 24084 22024
rect 24400 22015 24452 22024
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24400 21972 24452 21981
rect 24952 21972 25004 22024
rect 26240 21972 26292 22024
rect 27528 21972 27580 22024
rect 1860 21947 1912 21956
rect 1860 21913 1869 21947
rect 1869 21913 1903 21947
rect 1903 21913 1912 21947
rect 1860 21904 1912 21913
rect 22744 21947 22796 21956
rect 22744 21913 22761 21947
rect 22761 21913 22796 21947
rect 22744 21904 22796 21913
rect 3424 21836 3476 21888
rect 23756 21836 23808 21888
rect 25964 21879 26016 21888
rect 25964 21845 25973 21879
rect 25973 21845 26007 21879
rect 26007 21845 26016 21879
rect 25964 21836 26016 21845
rect 26516 21904 26568 21956
rect 28632 21972 28684 22024
rect 28080 21904 28132 21956
rect 29828 21904 29880 21956
rect 31392 21972 31444 22024
rect 35348 22040 35400 22092
rect 37648 22040 37700 22092
rect 38016 22040 38068 22092
rect 33508 22015 33560 22024
rect 33508 21981 33517 22015
rect 33517 21981 33551 22015
rect 33551 21981 33560 22015
rect 33508 21972 33560 21981
rect 34612 21972 34664 22024
rect 36084 22015 36136 22024
rect 36084 21981 36118 22015
rect 36118 21981 36136 22015
rect 36084 21972 36136 21981
rect 37924 21972 37976 22024
rect 27804 21879 27856 21888
rect 27804 21845 27813 21879
rect 27813 21845 27847 21879
rect 27847 21845 27856 21879
rect 27804 21836 27856 21845
rect 29000 21836 29052 21888
rect 30932 21879 30984 21888
rect 30932 21845 30941 21879
rect 30941 21845 30975 21879
rect 30975 21845 30984 21879
rect 30932 21836 30984 21845
rect 32404 21836 32456 21888
rect 38016 21879 38068 21888
rect 38016 21845 38025 21879
rect 38025 21845 38059 21879
rect 38059 21845 38068 21879
rect 38016 21836 38068 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 17224 21632 17276 21684
rect 22652 21632 22704 21684
rect 22744 21632 22796 21684
rect 24124 21632 24176 21684
rect 26516 21632 26568 21684
rect 13820 21607 13872 21616
rect 13820 21573 13829 21607
rect 13829 21573 13863 21607
rect 13863 21573 13872 21607
rect 13820 21564 13872 21573
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 14464 21539 14516 21548
rect 14464 21505 14473 21539
rect 14473 21505 14507 21539
rect 14507 21505 14516 21539
rect 14464 21496 14516 21505
rect 24308 21564 24360 21616
rect 24400 21564 24452 21616
rect 17408 21496 17460 21548
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 25964 21496 26016 21548
rect 3056 21292 3108 21344
rect 14280 21335 14332 21344
rect 14280 21301 14289 21335
rect 14289 21301 14323 21335
rect 14323 21301 14332 21335
rect 14280 21292 14332 21301
rect 14556 21292 14608 21344
rect 16488 21292 16540 21344
rect 23572 21428 23624 21480
rect 28264 21632 28316 21684
rect 29828 21675 29880 21684
rect 27528 21564 27580 21616
rect 29828 21641 29837 21675
rect 29837 21641 29871 21675
rect 29871 21641 29880 21675
rect 29828 21632 29880 21641
rect 32220 21632 32272 21684
rect 32772 21632 32824 21684
rect 34060 21632 34112 21684
rect 37372 21632 37424 21684
rect 27344 21539 27396 21548
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 29460 21496 29512 21548
rect 35900 21564 35952 21616
rect 33968 21496 34020 21548
rect 27160 21428 27212 21480
rect 22652 21360 22704 21412
rect 24768 21360 24820 21412
rect 26332 21360 26384 21412
rect 27620 21428 27672 21480
rect 32312 21428 32364 21480
rect 32956 21428 33008 21480
rect 34796 21428 34848 21480
rect 35348 21428 35400 21480
rect 27804 21360 27856 21412
rect 31944 21360 31996 21412
rect 36452 21539 36504 21548
rect 36452 21505 36461 21539
rect 36461 21505 36495 21539
rect 36495 21505 36504 21539
rect 36636 21539 36688 21548
rect 36452 21496 36504 21505
rect 36636 21505 36644 21539
rect 36644 21505 36678 21539
rect 36678 21505 36688 21539
rect 36636 21496 36688 21505
rect 36912 21496 36964 21548
rect 37004 21496 37056 21548
rect 37464 21496 37516 21548
rect 37556 21539 37608 21548
rect 37556 21505 37565 21539
rect 37565 21505 37599 21539
rect 37599 21505 37608 21539
rect 37832 21539 37884 21548
rect 37556 21496 37608 21505
rect 37832 21505 37840 21539
rect 37840 21505 37874 21539
rect 37874 21505 37884 21539
rect 37832 21496 37884 21505
rect 37924 21539 37976 21548
rect 37924 21505 37933 21539
rect 37933 21505 37967 21539
rect 37967 21505 37976 21539
rect 37924 21496 37976 21505
rect 38108 21496 38160 21548
rect 37004 21360 37056 21412
rect 18788 21292 18840 21344
rect 24308 21335 24360 21344
rect 24308 21301 24317 21335
rect 24317 21301 24351 21335
rect 24351 21301 24360 21335
rect 24308 21292 24360 21301
rect 24492 21292 24544 21344
rect 28724 21292 28776 21344
rect 33508 21292 33560 21344
rect 36084 21335 36136 21344
rect 36084 21301 36093 21335
rect 36093 21301 36127 21335
rect 36127 21301 36136 21335
rect 36084 21292 36136 21301
rect 37372 21292 37424 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2228 21088 2280 21140
rect 13820 21088 13872 21140
rect 14556 21020 14608 21072
rect 16672 21020 16724 21072
rect 15016 20952 15068 21004
rect 23572 21088 23624 21140
rect 23664 21088 23716 21140
rect 31024 21088 31076 21140
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 34152 21131 34204 21140
rect 34152 21097 34161 21131
rect 34161 21097 34195 21131
rect 34195 21097 34204 21131
rect 34152 21088 34204 21097
rect 21364 21020 21416 21072
rect 27344 21020 27396 21072
rect 36912 21088 36964 21140
rect 37832 21088 37884 21140
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 15660 20884 15712 20936
rect 17132 20884 17184 20936
rect 20076 20952 20128 21004
rect 32956 20952 33008 21004
rect 35348 20995 35400 21004
rect 18052 20927 18104 20936
rect 18052 20893 18061 20927
rect 18061 20893 18095 20927
rect 18095 20893 18104 20927
rect 18052 20884 18104 20893
rect 24400 20884 24452 20936
rect 32404 20927 32456 20936
rect 32404 20893 32413 20927
rect 32413 20893 32447 20927
rect 32447 20893 32456 20927
rect 32404 20884 32456 20893
rect 34152 20884 34204 20936
rect 35348 20961 35357 20995
rect 35357 20961 35391 20995
rect 35391 20961 35400 20995
rect 35348 20952 35400 20961
rect 36820 20884 36872 20936
rect 37004 20927 37056 20936
rect 37004 20893 37008 20927
rect 37008 20893 37042 20927
rect 37042 20893 37056 20927
rect 37004 20884 37056 20893
rect 37648 20952 37700 21004
rect 22928 20816 22980 20868
rect 27160 20816 27212 20868
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 1860 20748 1912 20800
rect 14372 20748 14424 20800
rect 15660 20791 15712 20800
rect 15660 20757 15669 20791
rect 15669 20757 15703 20791
rect 15703 20757 15712 20791
rect 15660 20748 15712 20757
rect 17132 20748 17184 20800
rect 18236 20791 18288 20800
rect 18236 20757 18245 20791
rect 18245 20757 18279 20791
rect 18279 20757 18288 20791
rect 18236 20748 18288 20757
rect 23572 20748 23624 20800
rect 24676 20748 24728 20800
rect 25136 20748 25188 20800
rect 31392 20791 31444 20800
rect 31392 20757 31401 20791
rect 31401 20757 31435 20791
rect 31435 20757 31444 20791
rect 37832 20884 37884 20936
rect 38108 20927 38160 20936
rect 38108 20893 38117 20927
rect 38117 20893 38151 20927
rect 38151 20893 38160 20927
rect 38108 20884 38160 20893
rect 34704 20791 34756 20800
rect 31392 20748 31444 20757
rect 34704 20757 34713 20791
rect 34713 20757 34747 20791
rect 34747 20757 34756 20791
rect 34704 20748 34756 20757
rect 35992 20748 36044 20800
rect 36176 20791 36228 20800
rect 36176 20757 36185 20791
rect 36185 20757 36219 20791
rect 36219 20757 36228 20791
rect 36176 20748 36228 20757
rect 36452 20748 36504 20800
rect 37648 20748 37700 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 13544 20587 13596 20596
rect 13544 20553 13553 20587
rect 13553 20553 13587 20587
rect 13587 20553 13596 20587
rect 13544 20544 13596 20553
rect 17408 20587 17460 20596
rect 14280 20519 14332 20528
rect 14280 20485 14314 20519
rect 14314 20485 14332 20519
rect 14280 20476 14332 20485
rect 17408 20553 17417 20587
rect 17417 20553 17451 20587
rect 17451 20553 17460 20587
rect 17408 20544 17460 20553
rect 18052 20544 18104 20596
rect 23480 20587 23532 20596
rect 23480 20553 23489 20587
rect 23489 20553 23523 20587
rect 23523 20553 23532 20587
rect 23480 20544 23532 20553
rect 23664 20544 23716 20596
rect 25228 20587 25280 20596
rect 25228 20553 25237 20587
rect 25237 20553 25271 20587
rect 25271 20553 25280 20587
rect 25228 20544 25280 20553
rect 27436 20544 27488 20596
rect 36728 20587 36780 20596
rect 36728 20553 36737 20587
rect 36737 20553 36771 20587
rect 36771 20553 36780 20587
rect 36728 20544 36780 20553
rect 37372 20544 37424 20596
rect 1860 20451 1912 20460
rect 1860 20417 1869 20451
rect 1869 20417 1903 20451
rect 1903 20417 1912 20451
rect 1860 20408 1912 20417
rect 2780 20408 2832 20460
rect 17224 20451 17276 20460
rect 13912 20340 13964 20392
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 18236 20476 18288 20528
rect 20536 20476 20588 20528
rect 22928 20519 22980 20528
rect 22928 20485 22937 20519
rect 22937 20485 22971 20519
rect 22971 20485 22980 20519
rect 22928 20476 22980 20485
rect 24400 20476 24452 20528
rect 18604 20408 18656 20460
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20260 20408 20312 20417
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 22192 20408 22244 20460
rect 23756 20408 23808 20460
rect 23388 20383 23440 20392
rect 16488 20272 16540 20324
rect 23388 20349 23414 20383
rect 23414 20349 23440 20383
rect 23388 20340 23440 20349
rect 22652 20272 22704 20324
rect 38384 20476 38436 20528
rect 27712 20408 27764 20460
rect 29736 20408 29788 20460
rect 32312 20408 32364 20460
rect 37372 20408 37424 20460
rect 37648 20451 37700 20460
rect 37648 20417 37657 20451
rect 37657 20417 37691 20451
rect 37691 20417 37700 20451
rect 37648 20408 37700 20417
rect 37740 20451 37792 20460
rect 37740 20417 37785 20451
rect 37785 20417 37792 20451
rect 37740 20408 37792 20417
rect 37924 20451 37976 20460
rect 37924 20417 37933 20451
rect 37933 20417 37967 20451
rect 37967 20417 37976 20451
rect 37924 20408 37976 20417
rect 30932 20383 30984 20392
rect 30932 20349 30941 20383
rect 30941 20349 30975 20383
rect 30975 20349 30984 20383
rect 30932 20340 30984 20349
rect 33048 20383 33100 20392
rect 33048 20349 33057 20383
rect 33057 20349 33091 20383
rect 33091 20349 33100 20383
rect 33048 20340 33100 20349
rect 27528 20272 27580 20324
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 16672 20204 16724 20256
rect 19984 20204 20036 20256
rect 23756 20204 23808 20256
rect 27712 20247 27764 20256
rect 27712 20213 27721 20247
rect 27721 20213 27755 20247
rect 27755 20213 27764 20247
rect 27712 20204 27764 20213
rect 38016 20272 38068 20324
rect 37280 20247 37332 20256
rect 37280 20213 37289 20247
rect 37289 20213 37323 20247
rect 37323 20213 37332 20247
rect 37280 20204 37332 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 14464 20000 14516 20052
rect 14924 20000 14976 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 17224 20000 17276 20052
rect 19432 20000 19484 20052
rect 24400 20000 24452 20052
rect 24676 20000 24728 20052
rect 29736 20043 29788 20052
rect 1860 19728 1912 19780
rect 10324 19796 10376 19848
rect 13452 19796 13504 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 15200 19728 15252 19780
rect 15936 19796 15988 19848
rect 16672 19796 16724 19848
rect 20260 19864 20312 19916
rect 22652 19932 22704 19984
rect 22928 19932 22980 19984
rect 29736 20009 29745 20043
rect 29745 20009 29779 20043
rect 29779 20009 29788 20043
rect 29736 20000 29788 20009
rect 32956 20043 33008 20052
rect 32956 20009 32965 20043
rect 32965 20009 32999 20043
rect 32999 20009 33008 20043
rect 32956 20000 33008 20009
rect 23572 19864 23624 19916
rect 23756 19907 23808 19916
rect 23756 19873 23765 19907
rect 23765 19873 23799 19907
rect 23799 19873 23808 19907
rect 23756 19864 23808 19873
rect 27620 19864 27672 19916
rect 37280 19932 37332 19984
rect 38016 19975 38068 19984
rect 38016 19941 38025 19975
rect 38025 19941 38059 19975
rect 38059 19941 38068 19975
rect 38016 19932 38068 19941
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 22744 19796 22796 19848
rect 24216 19796 24268 19848
rect 24860 19796 24912 19848
rect 27528 19796 27580 19848
rect 28816 19864 28868 19916
rect 28954 19864 29006 19916
rect 31392 19864 31444 19916
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 1952 19660 2004 19712
rect 3884 19703 3936 19712
rect 3884 19669 3893 19703
rect 3893 19669 3927 19703
rect 3927 19669 3936 19703
rect 3884 19660 3936 19669
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 18604 19728 18656 19780
rect 19340 19728 19392 19780
rect 22008 19771 22060 19780
rect 22008 19737 22017 19771
rect 22017 19737 22051 19771
rect 22051 19737 22060 19771
rect 22008 19728 22060 19737
rect 16488 19660 16540 19712
rect 19984 19660 20036 19712
rect 21272 19660 21324 19712
rect 29092 19796 29144 19848
rect 36084 19796 36136 19848
rect 36176 19796 36228 19848
rect 22376 19703 22428 19712
rect 22376 19669 22385 19703
rect 22385 19669 22419 19703
rect 22419 19669 22428 19703
rect 23572 19703 23624 19712
rect 22376 19660 22428 19669
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 28908 19660 28960 19712
rect 32404 19703 32456 19712
rect 32404 19669 32413 19703
rect 32413 19669 32447 19703
rect 32447 19669 32456 19703
rect 32404 19660 32456 19669
rect 36360 19660 36412 19712
rect 38108 19660 38160 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3700 19456 3752 19508
rect 15660 19456 15712 19508
rect 19248 19456 19300 19508
rect 20260 19456 20312 19508
rect 22376 19456 22428 19508
rect 23572 19456 23624 19508
rect 29092 19499 29144 19508
rect 29092 19465 29101 19499
rect 29101 19465 29135 19499
rect 29135 19465 29144 19499
rect 29092 19456 29144 19465
rect 3884 19388 3936 19440
rect 13728 19388 13780 19440
rect 16672 19388 16724 19440
rect 18880 19388 18932 19440
rect 22928 19388 22980 19440
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 2872 19320 2924 19372
rect 13912 19363 13964 19372
rect 2964 19252 3016 19304
rect 3056 19252 3108 19304
rect 13912 19329 13921 19363
rect 13921 19329 13955 19363
rect 13955 19329 13964 19363
rect 13912 19320 13964 19329
rect 14188 19363 14240 19372
rect 14188 19329 14222 19363
rect 14222 19329 14240 19363
rect 14188 19320 14240 19329
rect 20168 19320 20220 19372
rect 21088 19320 21140 19372
rect 24676 19388 24728 19440
rect 27620 19431 27672 19440
rect 27620 19397 27629 19431
rect 27629 19397 27663 19431
rect 27663 19397 27672 19431
rect 27620 19388 27672 19397
rect 36084 19388 36136 19440
rect 24308 19320 24360 19372
rect 19984 19252 20036 19304
rect 20628 19252 20680 19304
rect 9312 19184 9364 19236
rect 18696 19184 18748 19236
rect 20812 19227 20864 19236
rect 3056 19116 3108 19168
rect 3792 19116 3844 19168
rect 16488 19116 16540 19168
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 20812 19193 20821 19227
rect 20821 19193 20855 19227
rect 20855 19193 20864 19227
rect 20812 19184 20864 19193
rect 22928 19227 22980 19236
rect 22928 19193 22937 19227
rect 22937 19193 22971 19227
rect 22971 19193 22980 19227
rect 22928 19184 22980 19193
rect 23848 19184 23900 19236
rect 36452 19363 36504 19372
rect 36452 19329 36461 19363
rect 36461 19329 36495 19363
rect 36495 19329 36504 19363
rect 36452 19320 36504 19329
rect 28632 19295 28684 19304
rect 28632 19261 28641 19295
rect 28641 19261 28675 19295
rect 28675 19261 28684 19295
rect 28632 19252 28684 19261
rect 28908 19227 28960 19236
rect 28908 19193 28917 19227
rect 28917 19193 28951 19227
rect 28951 19193 28960 19227
rect 28908 19184 28960 19193
rect 22284 19116 22336 19168
rect 23388 19116 23440 19168
rect 23940 19116 23992 19168
rect 27620 19116 27672 19168
rect 34796 19159 34848 19168
rect 34796 19125 34805 19159
rect 34805 19125 34839 19159
rect 34839 19125 34848 19159
rect 34796 19116 34848 19125
rect 36360 19116 36412 19168
rect 37280 19159 37332 19168
rect 37280 19125 37289 19159
rect 37289 19125 37323 19159
rect 37323 19125 37332 19159
rect 37280 19116 37332 19125
rect 38016 19159 38068 19168
rect 38016 19125 38025 19159
rect 38025 19125 38059 19159
rect 38059 19125 38068 19159
rect 38016 19116 38068 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3056 18912 3108 18964
rect 3516 18912 3568 18964
rect 15936 18912 15988 18964
rect 20168 18955 20220 18964
rect 2872 18844 2924 18896
rect 4068 18844 4120 18896
rect 19340 18844 19392 18896
rect 20168 18921 20177 18955
rect 20177 18921 20211 18955
rect 20211 18921 20220 18955
rect 20168 18912 20220 18921
rect 22008 18912 22060 18964
rect 22192 18955 22244 18964
rect 22192 18921 22201 18955
rect 22201 18921 22235 18955
rect 22235 18921 22244 18955
rect 22192 18912 22244 18921
rect 20720 18844 20772 18896
rect 20904 18844 20956 18896
rect 3332 18776 3384 18828
rect 3976 18776 4028 18828
rect 19432 18776 19484 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 3056 18708 3108 18760
rect 3792 18751 3844 18760
rect 3792 18717 3801 18751
rect 3801 18717 3835 18751
rect 3835 18717 3844 18751
rect 3792 18708 3844 18717
rect 2964 18640 3016 18692
rect 14464 18708 14516 18760
rect 14924 18751 14976 18760
rect 7472 18640 7524 18692
rect 13360 18683 13412 18692
rect 3240 18572 3292 18624
rect 5448 18572 5500 18624
rect 11796 18572 11848 18624
rect 13360 18649 13369 18683
rect 13369 18649 13403 18683
rect 13403 18649 13412 18683
rect 13360 18640 13412 18649
rect 14556 18640 14608 18692
rect 14924 18717 14933 18751
rect 14933 18717 14967 18751
rect 14967 18717 14976 18751
rect 14924 18708 14976 18717
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15200 18708 15252 18717
rect 18236 18708 18288 18760
rect 20444 18776 20496 18828
rect 37832 18844 37884 18896
rect 37372 18776 37424 18828
rect 16304 18640 16356 18692
rect 19708 18683 19760 18692
rect 19708 18649 19717 18683
rect 19717 18649 19751 18683
rect 19751 18649 19760 18683
rect 19708 18640 19760 18649
rect 20168 18708 20220 18760
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 21732 18751 21784 18760
rect 20628 18640 20680 18692
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 21916 18751 21968 18760
rect 21916 18717 21925 18751
rect 21925 18717 21959 18751
rect 21959 18717 21968 18751
rect 21916 18708 21968 18717
rect 27712 18751 27764 18760
rect 27712 18717 27721 18751
rect 27721 18717 27755 18751
rect 27755 18717 27764 18751
rect 27712 18708 27764 18717
rect 28080 18708 28132 18760
rect 28632 18708 28684 18760
rect 30104 18708 30156 18760
rect 32404 18751 32456 18760
rect 24860 18683 24912 18692
rect 16672 18572 16724 18624
rect 17500 18572 17552 18624
rect 24860 18649 24869 18683
rect 24869 18649 24903 18683
rect 24903 18649 24912 18683
rect 24860 18640 24912 18649
rect 25044 18683 25096 18692
rect 25044 18649 25053 18683
rect 25053 18649 25087 18683
rect 25087 18649 25096 18683
rect 25044 18640 25096 18649
rect 25780 18640 25832 18692
rect 32404 18717 32413 18751
rect 32413 18717 32447 18751
rect 32447 18717 32456 18751
rect 32404 18708 32456 18717
rect 21088 18572 21140 18624
rect 27620 18572 27672 18624
rect 31852 18615 31904 18624
rect 31852 18581 31861 18615
rect 31861 18581 31895 18615
rect 31895 18581 31904 18615
rect 31852 18572 31904 18581
rect 32588 18615 32640 18624
rect 32588 18581 32597 18615
rect 32597 18581 32631 18615
rect 32631 18581 32640 18615
rect 32588 18572 32640 18581
rect 34796 18572 34848 18624
rect 35716 18572 35768 18624
rect 37280 18708 37332 18760
rect 38108 18751 38160 18760
rect 38108 18717 38117 18751
rect 38117 18717 38151 18751
rect 38151 18717 38160 18751
rect 38108 18708 38160 18717
rect 37372 18572 37424 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1400 18368 1452 18420
rect 2228 18343 2280 18352
rect 2228 18309 2237 18343
rect 2237 18309 2271 18343
rect 2271 18309 2280 18343
rect 2228 18300 2280 18309
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3516 18275 3568 18284
rect 3332 18232 3384 18241
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 10324 18368 10376 18420
rect 13452 18411 13504 18420
rect 13452 18377 13461 18411
rect 13461 18377 13495 18411
rect 13495 18377 13504 18411
rect 13452 18368 13504 18377
rect 14188 18411 14240 18420
rect 14188 18377 14197 18411
rect 14197 18377 14231 18411
rect 14231 18377 14240 18411
rect 14188 18368 14240 18377
rect 16948 18368 17000 18420
rect 19984 18368 20036 18420
rect 21272 18411 21324 18420
rect 9312 18300 9364 18352
rect 17132 18300 17184 18352
rect 19432 18300 19484 18352
rect 9496 18275 9548 18284
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 10048 18232 10100 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 13176 18232 13228 18284
rect 14372 18275 14424 18284
rect 9128 18028 9180 18080
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 13268 18096 13320 18148
rect 10048 18028 10100 18080
rect 10232 18028 10284 18080
rect 11796 18028 11848 18080
rect 12256 18028 12308 18080
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 19800 18275 19852 18284
rect 19800 18241 19809 18275
rect 19809 18241 19843 18275
rect 19843 18241 19852 18275
rect 20536 18300 20588 18352
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 21732 18368 21784 18420
rect 20996 18300 21048 18352
rect 27528 18300 27580 18352
rect 19800 18232 19852 18241
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 21456 18232 21508 18284
rect 22192 18232 22244 18284
rect 25964 18232 26016 18284
rect 27620 18232 27672 18284
rect 14188 18164 14240 18216
rect 19616 18164 19668 18216
rect 19892 18207 19944 18216
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 19892 18164 19944 18173
rect 20444 18164 20496 18216
rect 21916 18207 21968 18216
rect 21916 18173 21925 18207
rect 21925 18173 21959 18207
rect 21959 18173 21968 18207
rect 21916 18164 21968 18173
rect 13544 18096 13596 18148
rect 19340 18071 19392 18080
rect 19340 18037 19349 18071
rect 19349 18037 19383 18071
rect 19383 18037 19392 18071
rect 19800 18071 19852 18080
rect 19340 18028 19392 18037
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 20628 18096 20680 18148
rect 24952 18164 25004 18216
rect 27160 18164 27212 18216
rect 28264 18164 28316 18216
rect 30104 18164 30156 18216
rect 34520 18275 34572 18284
rect 34520 18241 34529 18275
rect 34529 18241 34563 18275
rect 34563 18241 34572 18275
rect 34520 18232 34572 18241
rect 35716 18275 35768 18284
rect 35716 18241 35725 18275
rect 35725 18241 35759 18275
rect 35759 18241 35768 18275
rect 35716 18232 35768 18241
rect 36360 18232 36412 18284
rect 32312 18164 32364 18216
rect 24216 18096 24268 18148
rect 25044 18096 25096 18148
rect 21732 18028 21784 18080
rect 22192 18028 22244 18080
rect 29276 18096 29328 18148
rect 30288 18139 30340 18148
rect 30288 18105 30297 18139
rect 30297 18105 30331 18139
rect 30331 18105 30340 18139
rect 30288 18096 30340 18105
rect 35808 18096 35860 18148
rect 36268 18096 36320 18148
rect 36636 18139 36688 18148
rect 36636 18105 36645 18139
rect 36645 18105 36679 18139
rect 36679 18105 36688 18139
rect 36636 18096 36688 18105
rect 27252 18028 27304 18080
rect 31116 18071 31168 18080
rect 31116 18037 31125 18071
rect 31125 18037 31159 18071
rect 31159 18037 31168 18071
rect 31116 18028 31168 18037
rect 34796 18028 34848 18080
rect 37280 18071 37332 18080
rect 37280 18037 37289 18071
rect 37289 18037 37323 18071
rect 37323 18037 37332 18071
rect 37280 18028 37332 18037
rect 38016 18071 38068 18080
rect 38016 18037 38025 18071
rect 38025 18037 38059 18071
rect 38059 18037 38068 18071
rect 38016 18028 38068 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1492 17867 1544 17876
rect 1492 17833 1501 17867
rect 1501 17833 1535 17867
rect 1535 17833 1544 17867
rect 1492 17824 1544 17833
rect 3056 17824 3108 17876
rect 3516 17824 3568 17876
rect 9588 17824 9640 17876
rect 3332 17756 3384 17808
rect 6368 17756 6420 17808
rect 11060 17756 11112 17808
rect 12072 17824 12124 17876
rect 12440 17824 12492 17876
rect 12624 17824 12676 17876
rect 13452 17824 13504 17876
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 19800 17824 19852 17876
rect 7380 17688 7432 17740
rect 10140 17688 10192 17740
rect 20720 17824 20772 17876
rect 22560 17824 22612 17876
rect 27620 17824 27672 17876
rect 13544 17688 13596 17740
rect 19892 17688 19944 17740
rect 20444 17731 20496 17740
rect 20444 17697 20453 17731
rect 20453 17697 20487 17731
rect 20487 17697 20496 17731
rect 20444 17688 20496 17697
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3700 17620 3752 17672
rect 5448 17620 5500 17672
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 7288 17620 7340 17672
rect 10324 17620 10376 17672
rect 10968 17620 11020 17672
rect 11152 17663 11204 17672
rect 11152 17629 11161 17663
rect 11161 17629 11195 17663
rect 11195 17629 11204 17663
rect 11152 17620 11204 17629
rect 3332 17552 3384 17604
rect 7564 17595 7616 17604
rect 6368 17527 6420 17536
rect 6368 17493 6377 17527
rect 6377 17493 6411 17527
rect 6411 17493 6420 17527
rect 6368 17484 6420 17493
rect 7564 17561 7573 17595
rect 7573 17561 7607 17595
rect 7607 17561 7616 17595
rect 7564 17552 7616 17561
rect 10784 17484 10836 17536
rect 11796 17484 11848 17536
rect 15936 17620 15988 17672
rect 18788 17620 18840 17672
rect 20076 17620 20128 17672
rect 20352 17663 20404 17672
rect 20352 17629 20361 17663
rect 20361 17629 20395 17663
rect 20395 17629 20404 17663
rect 20352 17620 20404 17629
rect 13176 17595 13228 17604
rect 13176 17561 13185 17595
rect 13185 17561 13219 17595
rect 13219 17561 13228 17595
rect 13176 17552 13228 17561
rect 13452 17552 13504 17604
rect 16396 17552 16448 17604
rect 19708 17552 19760 17604
rect 16304 17484 16356 17536
rect 16580 17484 16632 17536
rect 20444 17484 20496 17536
rect 20904 17756 20956 17808
rect 21916 17756 21968 17808
rect 23020 17756 23072 17808
rect 25964 17756 26016 17808
rect 20812 17688 20864 17740
rect 21088 17688 21140 17740
rect 20628 17663 20680 17672
rect 20628 17629 20637 17663
rect 20637 17629 20671 17663
rect 20671 17629 20680 17663
rect 20628 17620 20680 17629
rect 21272 17620 21324 17672
rect 22008 17688 22060 17740
rect 21456 17552 21508 17604
rect 24860 17620 24912 17672
rect 26148 17620 26200 17672
rect 30656 17824 30708 17876
rect 36176 17824 36228 17876
rect 36820 17824 36872 17876
rect 30472 17799 30524 17808
rect 30472 17765 30481 17799
rect 30481 17765 30515 17799
rect 30515 17765 30524 17799
rect 30472 17756 30524 17765
rect 36084 17799 36136 17808
rect 36084 17765 36093 17799
rect 36093 17765 36127 17799
rect 36127 17765 36136 17799
rect 36084 17756 36136 17765
rect 30380 17620 30432 17672
rect 30932 17620 30984 17672
rect 26424 17552 26476 17604
rect 29644 17595 29696 17604
rect 22376 17484 22428 17536
rect 25136 17527 25188 17536
rect 25136 17493 25145 17527
rect 25145 17493 25179 17527
rect 25179 17493 25188 17527
rect 25136 17484 25188 17493
rect 25596 17484 25648 17536
rect 29644 17561 29653 17595
rect 29653 17561 29687 17595
rect 29687 17561 29696 17595
rect 29644 17552 29696 17561
rect 30104 17595 30156 17604
rect 30104 17561 30113 17595
rect 30113 17561 30147 17595
rect 30147 17561 30156 17595
rect 30104 17552 30156 17561
rect 31116 17552 31168 17604
rect 31852 17552 31904 17604
rect 34428 17552 34480 17604
rect 34796 17552 34848 17604
rect 35900 17552 35952 17604
rect 27068 17484 27120 17536
rect 31576 17484 31628 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 3976 17280 4028 17332
rect 6552 17280 6604 17332
rect 12072 17280 12124 17332
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 14556 17280 14608 17332
rect 16580 17280 16632 17332
rect 18420 17280 18472 17332
rect 4068 17144 4120 17196
rect 6920 17144 6972 17196
rect 12348 17212 12400 17264
rect 8944 17144 8996 17196
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 11060 17144 11112 17196
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 12532 17144 12584 17196
rect 12716 17144 12768 17196
rect 18328 17212 18380 17264
rect 18512 17255 18564 17264
rect 18512 17221 18521 17255
rect 18521 17221 18555 17255
rect 18555 17221 18564 17255
rect 18512 17212 18564 17221
rect 18788 17255 18840 17264
rect 18788 17221 18797 17255
rect 18797 17221 18831 17255
rect 18831 17221 18840 17255
rect 18788 17212 18840 17221
rect 19432 17280 19484 17332
rect 20352 17280 20404 17332
rect 20444 17280 20496 17332
rect 21824 17323 21876 17332
rect 19248 17212 19300 17264
rect 20260 17212 20312 17264
rect 14372 17144 14424 17196
rect 6828 17076 6880 17128
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 8116 17076 8168 17128
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 10048 17008 10100 17060
rect 14924 17076 14976 17128
rect 19064 17134 19116 17186
rect 20904 17144 20956 17196
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 21272 17212 21324 17264
rect 21456 17144 21508 17196
rect 21824 17144 21876 17196
rect 22284 17187 22336 17196
rect 22284 17153 22293 17187
rect 22293 17153 22327 17187
rect 22327 17153 22336 17187
rect 22284 17144 22336 17153
rect 22652 17144 22704 17196
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 26976 17280 27028 17332
rect 30288 17280 30340 17332
rect 34520 17280 34572 17332
rect 35348 17323 35400 17332
rect 35348 17289 35357 17323
rect 35357 17289 35391 17323
rect 35391 17289 35400 17323
rect 35348 17280 35400 17289
rect 30656 17255 30708 17264
rect 30656 17221 30665 17255
rect 30665 17221 30699 17255
rect 30699 17221 30708 17255
rect 30656 17212 30708 17221
rect 30748 17212 30800 17264
rect 33968 17212 34020 17264
rect 24860 17187 24912 17196
rect 24860 17153 24869 17187
rect 24869 17153 24903 17187
rect 24903 17153 24912 17187
rect 24860 17144 24912 17153
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 13544 16983 13596 16992
rect 12900 16940 12952 16949
rect 13544 16949 13553 16983
rect 13553 16949 13587 16983
rect 13587 16949 13596 16983
rect 13544 16940 13596 16949
rect 17500 17008 17552 17060
rect 16120 16940 16172 16992
rect 19248 17076 19300 17128
rect 25596 17144 25648 17196
rect 25964 17187 26016 17196
rect 25964 17153 25973 17187
rect 25973 17153 26007 17187
rect 26007 17153 26016 17187
rect 25964 17144 26016 17153
rect 27712 17187 27764 17196
rect 27712 17153 27721 17187
rect 27721 17153 27755 17187
rect 27755 17153 27764 17187
rect 27712 17144 27764 17153
rect 29644 17144 29696 17196
rect 31576 17187 31628 17196
rect 18972 17008 19024 17060
rect 19708 17008 19760 17060
rect 20444 17008 20496 17060
rect 25136 17119 25188 17128
rect 25136 17085 25145 17119
rect 25145 17085 25179 17119
rect 25179 17085 25188 17119
rect 25136 17076 25188 17085
rect 27344 17076 27396 17128
rect 27988 17076 28040 17128
rect 30380 17076 30432 17128
rect 31576 17153 31585 17187
rect 31585 17153 31619 17187
rect 31619 17153 31628 17187
rect 31576 17144 31628 17153
rect 36084 17212 36136 17264
rect 37096 17212 37148 17264
rect 38292 17212 38344 17264
rect 37188 17144 37240 17196
rect 37280 17144 37332 17196
rect 33140 17076 33192 17128
rect 33232 17119 33284 17128
rect 33232 17085 33241 17119
rect 33241 17085 33275 17119
rect 33275 17085 33284 17119
rect 33232 17076 33284 17085
rect 20996 17008 21048 17060
rect 21916 17008 21968 17060
rect 22376 17008 22428 17060
rect 22468 17008 22520 17060
rect 23020 17008 23072 17060
rect 23664 17008 23716 17060
rect 21088 16940 21140 16992
rect 21732 16940 21784 16992
rect 24768 16940 24820 16992
rect 24952 16940 25004 16992
rect 25228 16940 25280 16992
rect 28540 17008 28592 17060
rect 34428 17008 34480 17060
rect 35348 17076 35400 17128
rect 36360 17076 36412 17128
rect 27804 16940 27856 16992
rect 29736 16940 29788 16992
rect 30748 16940 30800 16992
rect 31208 16940 31260 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 6276 16736 6328 16788
rect 6828 16736 6880 16788
rect 13084 16736 13136 16788
rect 16212 16779 16264 16788
rect 6552 16711 6604 16720
rect 6552 16677 6561 16711
rect 6561 16677 6595 16711
rect 6595 16677 6604 16711
rect 6552 16668 6604 16677
rect 7380 16600 7432 16652
rect 12256 16600 12308 16652
rect 12440 16668 12492 16720
rect 13360 16668 13412 16720
rect 15936 16668 15988 16720
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 19248 16736 19300 16788
rect 19708 16668 19760 16720
rect 22836 16736 22888 16788
rect 22376 16668 22428 16720
rect 13268 16600 13320 16652
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 1860 16507 1912 16516
rect 1860 16473 1869 16507
rect 1869 16473 1903 16507
rect 1903 16473 1912 16507
rect 1860 16464 1912 16473
rect 6276 16507 6328 16516
rect 6276 16473 6285 16507
rect 6285 16473 6319 16507
rect 6319 16473 6328 16507
rect 6276 16464 6328 16473
rect 7012 16507 7064 16516
rect 7012 16473 7021 16507
rect 7021 16473 7055 16507
rect 7055 16473 7064 16507
rect 7012 16464 7064 16473
rect 9496 16532 9548 16584
rect 9956 16532 10008 16584
rect 10784 16532 10836 16584
rect 12532 16532 12584 16584
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 16028 16600 16080 16652
rect 16948 16600 17000 16652
rect 18236 16600 18288 16652
rect 20260 16600 20312 16652
rect 20720 16600 20772 16652
rect 23296 16600 23348 16652
rect 26240 16736 26292 16788
rect 30472 16779 30524 16788
rect 30472 16745 30481 16779
rect 30481 16745 30515 16779
rect 30515 16745 30524 16779
rect 30472 16736 30524 16745
rect 16396 16532 16448 16584
rect 8300 16396 8352 16448
rect 10324 16464 10376 16516
rect 16304 16464 16356 16516
rect 16672 16532 16724 16584
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 17592 16532 17644 16584
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 21916 16575 21968 16584
rect 21916 16541 21925 16575
rect 21925 16541 21959 16575
rect 21959 16541 21968 16575
rect 21916 16532 21968 16541
rect 24768 16575 24820 16584
rect 24768 16541 24802 16575
rect 24802 16541 24820 16575
rect 21824 16464 21876 16516
rect 24768 16532 24820 16541
rect 26884 16575 26936 16584
rect 10692 16396 10744 16448
rect 12808 16396 12860 16448
rect 18144 16396 18196 16448
rect 18788 16396 18840 16448
rect 24952 16464 25004 16516
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 27068 16575 27120 16584
rect 27068 16541 27077 16575
rect 27077 16541 27111 16575
rect 27111 16541 27120 16575
rect 27068 16532 27120 16541
rect 27804 16575 27856 16584
rect 27804 16541 27838 16575
rect 27838 16541 27856 16575
rect 27804 16532 27856 16541
rect 27436 16464 27488 16516
rect 22376 16396 22428 16448
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 25412 16396 25464 16448
rect 26240 16396 26292 16448
rect 28172 16396 28224 16448
rect 30380 16600 30432 16652
rect 29736 16532 29788 16584
rect 34060 16736 34112 16788
rect 32312 16711 32364 16720
rect 32312 16677 32321 16711
rect 32321 16677 32355 16711
rect 32355 16677 32364 16711
rect 32312 16668 32364 16677
rect 33140 16668 33192 16720
rect 33968 16711 34020 16720
rect 33968 16677 33977 16711
rect 33977 16677 34011 16711
rect 34011 16677 34020 16711
rect 33968 16668 34020 16677
rect 34428 16668 34480 16720
rect 31208 16575 31260 16584
rect 31208 16541 31242 16575
rect 31242 16541 31260 16575
rect 31208 16532 31260 16541
rect 36084 16532 36136 16584
rect 36820 16532 36872 16584
rect 37004 16575 37056 16584
rect 37004 16541 37008 16575
rect 37008 16541 37042 16575
rect 37042 16541 37056 16575
rect 37004 16532 37056 16541
rect 37188 16575 37240 16584
rect 37188 16541 37197 16575
rect 37197 16541 37231 16575
rect 37231 16541 37240 16575
rect 37188 16532 37240 16541
rect 37372 16575 37424 16584
rect 37372 16541 37380 16575
rect 37380 16541 37414 16575
rect 37414 16541 37424 16575
rect 37372 16532 37424 16541
rect 37464 16575 37516 16584
rect 37464 16541 37473 16575
rect 37473 16541 37507 16575
rect 37507 16541 37516 16575
rect 37464 16532 37516 16541
rect 37648 16532 37700 16584
rect 38108 16575 38160 16584
rect 38108 16541 38117 16575
rect 38117 16541 38151 16575
rect 38151 16541 38160 16575
rect 38108 16532 38160 16541
rect 30012 16439 30064 16448
rect 30012 16405 30021 16439
rect 30021 16405 30055 16439
rect 30055 16405 30064 16439
rect 30012 16396 30064 16405
rect 32220 16464 32272 16516
rect 32312 16396 32364 16448
rect 34796 16396 34848 16448
rect 36176 16439 36228 16448
rect 36176 16405 36185 16439
rect 36185 16405 36219 16439
rect 36219 16405 36228 16439
rect 36176 16396 36228 16405
rect 36820 16439 36872 16448
rect 36820 16405 36829 16439
rect 36829 16405 36863 16439
rect 36863 16405 36872 16439
rect 36820 16396 36872 16405
rect 37372 16396 37424 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 6276 16056 6328 16108
rect 8116 16124 8168 16176
rect 13912 16192 13964 16244
rect 16764 16192 16816 16244
rect 18972 16192 19024 16244
rect 21640 16192 21692 16244
rect 22836 16192 22888 16244
rect 24860 16192 24912 16244
rect 26424 16235 26476 16244
rect 26424 16201 26433 16235
rect 26433 16201 26467 16235
rect 26467 16201 26476 16235
rect 26424 16192 26476 16201
rect 27712 16192 27764 16244
rect 28172 16235 28224 16244
rect 28172 16201 28181 16235
rect 28181 16201 28215 16235
rect 28215 16201 28224 16235
rect 28172 16192 28224 16201
rect 14372 16167 14424 16176
rect 14372 16133 14381 16167
rect 14381 16133 14415 16167
rect 14415 16133 14424 16167
rect 14372 16124 14424 16133
rect 8300 16099 8352 16108
rect 8300 16065 8334 16099
rect 8334 16065 8352 16099
rect 8300 16056 8352 16065
rect 10784 16099 10836 16108
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 13544 16056 13596 16108
rect 21548 16124 21600 16176
rect 22652 16124 22704 16176
rect 29460 16167 29512 16176
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 6920 15988 6972 16040
rect 7932 15988 7984 16040
rect 12440 15988 12492 16040
rect 17592 16056 17644 16108
rect 18144 16056 18196 16108
rect 21456 16056 21508 16108
rect 21824 16056 21876 16108
rect 22468 16056 22520 16108
rect 24952 16099 25004 16108
rect 16764 16031 16816 16040
rect 11888 15920 11940 15972
rect 12624 15920 12676 15972
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 16948 15988 17000 16040
rect 18788 16031 18840 16040
rect 18788 15997 18797 16031
rect 18797 15997 18831 16031
rect 18831 15997 18840 16031
rect 18788 15988 18840 15997
rect 19248 15988 19300 16040
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 2596 15852 2648 15904
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10876 15895 10928 15904
rect 10876 15861 10885 15895
rect 10885 15861 10919 15895
rect 10919 15861 10928 15895
rect 10876 15852 10928 15861
rect 10968 15852 11020 15904
rect 14280 15852 14332 15904
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 16028 15852 16080 15904
rect 20812 15920 20864 15972
rect 21916 15920 21968 15972
rect 22376 15920 22428 15972
rect 22928 16031 22980 16040
rect 22928 15997 22937 16031
rect 22937 15997 22971 16031
rect 22971 15997 22980 16031
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 22928 15988 22980 15997
rect 25872 16056 25924 16108
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 26976 16099 27028 16108
rect 26976 16065 26985 16099
rect 26985 16065 27019 16099
rect 27019 16065 27028 16099
rect 29460 16133 29469 16167
rect 29469 16133 29503 16167
rect 29503 16133 29512 16167
rect 29460 16124 29512 16133
rect 26976 16056 27028 16065
rect 27436 16099 27488 16108
rect 26884 15988 26936 16040
rect 27436 16065 27445 16099
rect 27445 16065 27479 16099
rect 27479 16065 27488 16099
rect 27436 16056 27488 16065
rect 33048 16056 33100 16108
rect 37004 16056 37056 16108
rect 33232 15988 33284 16040
rect 34244 15988 34296 16040
rect 35716 15988 35768 16040
rect 37280 16031 37332 16040
rect 34796 15963 34848 15972
rect 34796 15929 34805 15963
rect 34805 15929 34839 15963
rect 34839 15929 34848 15963
rect 34796 15920 34848 15929
rect 37280 15997 37289 16031
rect 37289 15997 37323 16031
rect 37323 15997 37332 16031
rect 37280 15988 37332 15997
rect 37464 15920 37516 15972
rect 21824 15852 21876 15904
rect 22468 15852 22520 15904
rect 22928 15852 22980 15904
rect 23296 15852 23348 15904
rect 25228 15852 25280 15904
rect 35624 15852 35676 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 7472 15648 7524 15700
rect 8944 15691 8996 15700
rect 8944 15657 8953 15691
rect 8953 15657 8987 15691
rect 8987 15657 8996 15691
rect 8944 15648 8996 15657
rect 9772 15648 9824 15700
rect 10692 15648 10744 15700
rect 11888 15691 11940 15700
rect 11888 15657 11897 15691
rect 11897 15657 11931 15691
rect 11931 15657 11940 15691
rect 11888 15648 11940 15657
rect 13084 15648 13136 15700
rect 14372 15648 14424 15700
rect 16212 15691 16264 15700
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 21824 15691 21876 15700
rect 13176 15623 13228 15632
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 13176 15589 13185 15623
rect 13185 15589 13219 15623
rect 13219 15589 13228 15623
rect 13176 15580 13228 15589
rect 14280 15580 14332 15632
rect 16856 15580 16908 15632
rect 17040 15580 17092 15632
rect 18236 15580 18288 15632
rect 1860 15419 1912 15428
rect 1860 15385 1869 15419
rect 1869 15385 1903 15419
rect 1903 15385 1912 15419
rect 1860 15376 1912 15385
rect 10876 15444 10928 15496
rect 12808 15512 12860 15564
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 16028 15555 16080 15564
rect 16028 15521 16037 15555
rect 16037 15521 16071 15555
rect 16071 15521 16080 15555
rect 16028 15512 16080 15521
rect 20720 15512 20772 15564
rect 20812 15555 20864 15564
rect 20812 15521 20821 15555
rect 20821 15521 20855 15555
rect 20855 15521 20864 15555
rect 20812 15512 20864 15521
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 11152 15308 11204 15360
rect 12256 15419 12308 15428
rect 12256 15385 12265 15419
rect 12265 15385 12299 15419
rect 12299 15385 12308 15419
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 14556 15487 14608 15496
rect 13268 15444 13320 15453
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 15200 15444 15252 15496
rect 12256 15376 12308 15385
rect 12900 15376 12952 15428
rect 13452 15376 13504 15428
rect 15660 15376 15712 15428
rect 16120 15444 16172 15496
rect 16396 15444 16448 15496
rect 18420 15444 18472 15496
rect 19064 15444 19116 15496
rect 19340 15444 19392 15496
rect 18512 15419 18564 15428
rect 18512 15385 18521 15419
rect 18521 15385 18555 15419
rect 18555 15385 18564 15419
rect 18512 15376 18564 15385
rect 16488 15308 16540 15360
rect 17500 15351 17552 15360
rect 17500 15317 17509 15351
rect 17509 15317 17543 15351
rect 17543 15317 17552 15351
rect 17500 15308 17552 15317
rect 21824 15657 21833 15691
rect 21833 15657 21867 15691
rect 21867 15657 21876 15691
rect 23296 15691 23348 15700
rect 21824 15648 21876 15657
rect 23296 15657 23305 15691
rect 23305 15657 23339 15691
rect 23339 15657 23348 15691
rect 23296 15648 23348 15657
rect 25228 15648 25280 15700
rect 35900 15648 35952 15700
rect 21732 15580 21784 15632
rect 22008 15512 22060 15564
rect 22468 15512 22520 15564
rect 21548 15444 21600 15496
rect 27068 15580 27120 15632
rect 30012 15444 30064 15496
rect 35624 15487 35676 15496
rect 35624 15453 35633 15487
rect 35633 15453 35667 15487
rect 35667 15453 35676 15487
rect 35624 15444 35676 15453
rect 37004 15487 37056 15496
rect 37004 15453 37008 15487
rect 37008 15453 37042 15487
rect 37042 15453 37056 15487
rect 37004 15444 37056 15453
rect 37188 15487 37240 15496
rect 37188 15453 37197 15487
rect 37197 15453 37231 15487
rect 37231 15453 37240 15487
rect 37188 15444 37240 15453
rect 37372 15487 37424 15496
rect 37372 15453 37380 15487
rect 37380 15453 37414 15487
rect 37414 15453 37424 15487
rect 37372 15444 37424 15453
rect 37464 15487 37516 15496
rect 37464 15453 37473 15487
rect 37473 15453 37507 15487
rect 37507 15453 37516 15487
rect 38108 15487 38160 15496
rect 37464 15444 37516 15453
rect 38108 15453 38117 15487
rect 38117 15453 38151 15487
rect 38151 15453 38160 15487
rect 38108 15444 38160 15453
rect 25964 15419 26016 15428
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 25964 15385 25973 15419
rect 25973 15385 26007 15419
rect 26007 15385 26016 15419
rect 25964 15376 26016 15385
rect 27068 15376 27120 15428
rect 33416 15376 33468 15428
rect 37096 15419 37148 15428
rect 26884 15351 26936 15360
rect 26884 15317 26893 15351
rect 26893 15317 26927 15351
rect 26927 15317 26936 15351
rect 26884 15308 26936 15317
rect 29000 15308 29052 15360
rect 37096 15385 37105 15419
rect 37105 15385 37139 15419
rect 37139 15385 37148 15419
rect 37096 15376 37148 15385
rect 37372 15308 37424 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2228 15104 2280 15156
rect 6276 15104 6328 15156
rect 9956 15104 10008 15156
rect 17316 15147 17368 15156
rect 11060 15036 11112 15088
rect 14372 15036 14424 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 14464 14968 14516 15020
rect 15292 14968 15344 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 18696 15104 18748 15156
rect 35716 15147 35768 15156
rect 17684 15036 17736 15088
rect 17960 15036 18012 15088
rect 18328 15036 18380 15088
rect 20536 15036 20588 15088
rect 22376 15036 22428 15088
rect 22652 15036 22704 15088
rect 25136 15036 25188 15088
rect 25504 15036 25556 15088
rect 25872 15036 25924 15088
rect 26884 15036 26936 15088
rect 35716 15113 35725 15147
rect 35725 15113 35759 15147
rect 35759 15113 35768 15147
rect 35716 15104 35768 15113
rect 37648 15104 37700 15156
rect 38016 15147 38068 15156
rect 38016 15113 38025 15147
rect 38025 15113 38059 15147
rect 38059 15113 38068 15147
rect 38016 15104 38068 15113
rect 37280 15079 37332 15088
rect 37280 15045 37289 15079
rect 37289 15045 37323 15079
rect 37323 15045 37332 15079
rect 37280 15036 37332 15045
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 15384 14900 15436 14952
rect 16028 14900 16080 14952
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 12992 14832 13044 14884
rect 13176 14875 13228 14884
rect 13176 14841 13185 14875
rect 13185 14841 13219 14875
rect 13219 14841 13228 14875
rect 13176 14832 13228 14841
rect 14740 14875 14792 14884
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 2504 14764 2556 14816
rect 12900 14764 12952 14816
rect 15660 14764 15712 14816
rect 16212 14832 16264 14884
rect 16856 14832 16908 14884
rect 16028 14764 16080 14816
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 17960 14832 18012 14884
rect 21548 14968 21600 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 28908 14968 28960 15020
rect 34704 15011 34756 15020
rect 34704 14977 34713 15011
rect 34713 14977 34747 15011
rect 34747 14977 34756 15011
rect 34704 14968 34756 14977
rect 18604 14900 18656 14952
rect 18788 14832 18840 14884
rect 18972 14832 19024 14884
rect 19340 14832 19392 14884
rect 21456 14832 21508 14884
rect 22284 14875 22336 14884
rect 18052 14764 18104 14816
rect 20536 14764 20588 14816
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 22284 14841 22293 14875
rect 22293 14841 22327 14875
rect 22327 14841 22336 14875
rect 22284 14832 22336 14841
rect 29920 14875 29972 14884
rect 29920 14841 29929 14875
rect 29929 14841 29963 14875
rect 29963 14841 29972 14875
rect 29920 14832 29972 14841
rect 30104 14900 30156 14952
rect 31760 14900 31812 14952
rect 36820 14832 36872 14884
rect 25228 14764 25280 14816
rect 25412 14764 25464 14816
rect 25780 14764 25832 14816
rect 27344 14764 27396 14816
rect 29184 14764 29236 14816
rect 34796 14764 34848 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 14464 14560 14516 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 16212 14560 16264 14612
rect 18052 14560 18104 14612
rect 23664 14560 23716 14612
rect 31760 14603 31812 14612
rect 31760 14569 31769 14603
rect 31769 14569 31803 14603
rect 31803 14569 31812 14603
rect 34060 14603 34112 14612
rect 31760 14560 31812 14569
rect 34060 14569 34069 14603
rect 34069 14569 34103 14603
rect 34103 14569 34112 14603
rect 34060 14560 34112 14569
rect 34704 14560 34756 14612
rect 38108 14603 38160 14612
rect 38108 14569 38117 14603
rect 38117 14569 38151 14603
rect 38151 14569 38160 14603
rect 38108 14560 38160 14569
rect 13912 14492 13964 14544
rect 14556 14492 14608 14544
rect 15660 14492 15712 14544
rect 18696 14492 18748 14544
rect 34428 14492 34480 14544
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 12992 14356 13044 14408
rect 14648 14356 14700 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 15476 14356 15528 14408
rect 25596 14424 25648 14476
rect 25964 14424 26016 14476
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 17868 14356 17920 14408
rect 30288 14356 30340 14408
rect 35992 14399 36044 14408
rect 35992 14365 36001 14399
rect 36001 14365 36035 14399
rect 36035 14365 36044 14399
rect 35992 14356 36044 14365
rect 37004 14399 37056 14408
rect 37004 14365 37008 14399
rect 37008 14365 37042 14399
rect 37042 14365 37056 14399
rect 37004 14356 37056 14365
rect 37188 14399 37240 14408
rect 37188 14365 37197 14399
rect 37197 14365 37231 14399
rect 37231 14365 37240 14399
rect 37188 14356 37240 14365
rect 37372 14399 37424 14408
rect 37372 14365 37380 14399
rect 37380 14365 37414 14399
rect 37414 14365 37424 14399
rect 37372 14356 37424 14365
rect 37464 14399 37516 14408
rect 37464 14365 37473 14399
rect 37473 14365 37507 14399
rect 37507 14365 37516 14399
rect 37464 14356 37516 14365
rect 1400 14288 1452 14340
rect 12348 14288 12400 14340
rect 12624 14288 12676 14340
rect 13084 14288 13136 14340
rect 14924 14288 14976 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2320 14220 2372 14272
rect 9864 14220 9916 14272
rect 12900 14220 12952 14272
rect 13360 14220 13412 14272
rect 16120 14220 16172 14272
rect 17040 14263 17092 14272
rect 17040 14229 17049 14263
rect 17049 14229 17083 14263
rect 17083 14229 17092 14263
rect 17040 14220 17092 14229
rect 17224 14220 17276 14272
rect 17408 14331 17460 14340
rect 17408 14297 17417 14331
rect 17417 14297 17451 14331
rect 17451 14297 17460 14331
rect 17408 14288 17460 14297
rect 17592 14288 17644 14340
rect 17776 14288 17828 14340
rect 21824 14288 21876 14340
rect 29368 14288 29420 14340
rect 34244 14288 34296 14340
rect 37096 14331 37148 14340
rect 37096 14297 37105 14331
rect 37105 14297 37139 14331
rect 37139 14297 37148 14331
rect 37096 14288 37148 14297
rect 37280 14288 37332 14340
rect 17868 14220 17920 14272
rect 29092 14220 29144 14272
rect 30196 14220 30248 14272
rect 36176 14263 36228 14272
rect 36176 14229 36185 14263
rect 36185 14229 36219 14263
rect 36219 14229 36228 14263
rect 36176 14220 36228 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 8300 14016 8352 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 13728 14016 13780 14068
rect 2504 13991 2556 14000
rect 2504 13957 2513 13991
rect 2513 13957 2547 13991
rect 2547 13957 2556 13991
rect 2504 13948 2556 13957
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 8116 13948 8168 14000
rect 12440 13991 12492 14000
rect 12440 13957 12449 13991
rect 12449 13957 12483 13991
rect 12483 13957 12492 13991
rect 12440 13948 12492 13957
rect 13268 13948 13320 14000
rect 13636 13948 13688 14000
rect 14464 13948 14516 14000
rect 14832 13948 14884 14000
rect 2780 13880 2832 13889
rect 9588 13923 9640 13932
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 11796 13880 11848 13932
rect 12532 13880 12584 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 13544 13880 13596 13932
rect 14188 13880 14240 13932
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 17684 14016 17736 14068
rect 17776 14016 17828 14068
rect 29092 14016 29144 14068
rect 29368 14059 29420 14068
rect 29368 14025 29377 14059
rect 29377 14025 29411 14059
rect 29411 14025 29420 14059
rect 29368 14016 29420 14025
rect 29920 14016 29972 14068
rect 30196 14059 30248 14068
rect 30196 14025 30205 14059
rect 30205 14025 30239 14059
rect 30239 14025 30248 14059
rect 30196 14016 30248 14025
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 16028 13923 16080 13932
rect 16028 13889 16037 13923
rect 16037 13889 16071 13923
rect 16071 13889 16080 13923
rect 16028 13880 16080 13889
rect 16120 13880 16172 13932
rect 17224 13948 17276 14000
rect 19340 13948 19392 14000
rect 22008 13948 22060 14000
rect 31760 14016 31812 14068
rect 34428 14059 34480 14068
rect 17132 13880 17184 13932
rect 17684 13880 17736 13932
rect 17960 13880 18012 13932
rect 19432 13880 19484 13932
rect 25964 13880 26016 13932
rect 26056 13923 26108 13932
rect 26056 13889 26065 13923
rect 26065 13889 26099 13923
rect 26099 13889 26108 13923
rect 29184 13923 29236 13932
rect 26056 13880 26108 13889
rect 29184 13889 29193 13923
rect 29193 13889 29227 13923
rect 29227 13889 29236 13923
rect 29184 13880 29236 13889
rect 30196 13880 30248 13932
rect 34428 14025 34437 14059
rect 34437 14025 34471 14059
rect 34471 14025 34480 14059
rect 34428 14016 34480 14025
rect 36084 14016 36136 14068
rect 37096 14016 37148 14068
rect 34796 13948 34848 14000
rect 30564 13880 30616 13932
rect 34152 13880 34204 13932
rect 35900 13880 35952 13932
rect 13268 13812 13320 13864
rect 15384 13812 15436 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 20720 13812 20772 13864
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 4068 13676 4120 13728
rect 10692 13676 10744 13728
rect 15568 13744 15620 13796
rect 15844 13787 15896 13796
rect 15384 13676 15436 13728
rect 15844 13753 15853 13787
rect 15853 13753 15887 13787
rect 15887 13753 15896 13787
rect 15844 13744 15896 13753
rect 16028 13744 16080 13796
rect 17500 13744 17552 13796
rect 20260 13744 20312 13796
rect 21364 13744 21416 13796
rect 30380 13744 30432 13796
rect 34336 13744 34388 13796
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 30932 13676 30984 13728
rect 38016 13719 38068 13728
rect 38016 13685 38025 13719
rect 38025 13685 38059 13719
rect 38059 13685 38068 13719
rect 38016 13676 38068 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2780 13472 2832 13524
rect 9588 13515 9640 13524
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 10692 13404 10744 13456
rect 3700 13336 3752 13388
rect 9496 13336 9548 13388
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 9404 13268 9456 13277
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 7932 13200 7984 13252
rect 8116 13200 8168 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 12256 13472 12308 13524
rect 13820 13472 13872 13524
rect 19984 13472 20036 13524
rect 24676 13515 24728 13524
rect 24676 13481 24685 13515
rect 24685 13481 24719 13515
rect 24719 13481 24728 13515
rect 24676 13472 24728 13481
rect 28540 13515 28592 13524
rect 28540 13481 28549 13515
rect 28549 13481 28583 13515
rect 28583 13481 28592 13515
rect 28540 13472 28592 13481
rect 30564 13472 30616 13524
rect 32036 13515 32088 13524
rect 32036 13481 32045 13515
rect 32045 13481 32079 13515
rect 32079 13481 32088 13515
rect 32036 13472 32088 13481
rect 35900 13472 35952 13524
rect 17132 13404 17184 13456
rect 30012 13447 30064 13456
rect 30012 13413 30021 13447
rect 30021 13413 30055 13447
rect 30055 13413 30064 13447
rect 30012 13404 30064 13413
rect 14740 13336 14792 13388
rect 15752 13336 15804 13388
rect 15936 13336 15988 13388
rect 17224 13336 17276 13388
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 12992 13268 13044 13320
rect 13084 13311 13136 13320
rect 13084 13277 13093 13311
rect 13093 13277 13127 13311
rect 13127 13277 13136 13311
rect 13084 13268 13136 13277
rect 13360 13268 13412 13320
rect 20720 13336 20772 13388
rect 24676 13336 24728 13388
rect 30104 13336 30156 13388
rect 34152 13336 34204 13388
rect 34336 13336 34388 13388
rect 37280 13336 37332 13388
rect 18420 13268 18472 13320
rect 18972 13268 19024 13320
rect 19340 13311 19392 13320
rect 19340 13277 19349 13311
rect 19349 13277 19383 13311
rect 19383 13277 19392 13311
rect 20812 13311 20864 13320
rect 19340 13268 19392 13277
rect 20812 13277 20821 13311
rect 20821 13277 20855 13311
rect 20855 13277 20864 13311
rect 20812 13268 20864 13277
rect 20996 13311 21048 13320
rect 20996 13277 21005 13311
rect 21005 13277 21039 13311
rect 21039 13277 21048 13311
rect 20996 13268 21048 13277
rect 15108 13200 15160 13252
rect 16672 13200 16724 13252
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 12532 13132 12584 13184
rect 14280 13132 14332 13184
rect 16856 13132 16908 13184
rect 19432 13200 19484 13252
rect 17316 13132 17368 13184
rect 17500 13175 17552 13184
rect 17500 13141 17509 13175
rect 17509 13141 17543 13175
rect 17543 13141 17552 13175
rect 17500 13132 17552 13141
rect 18880 13132 18932 13184
rect 21364 13268 21416 13320
rect 21824 13311 21876 13320
rect 21824 13277 21833 13311
rect 21833 13277 21867 13311
rect 21867 13277 21876 13311
rect 21824 13268 21876 13277
rect 24768 13268 24820 13320
rect 25596 13268 25648 13320
rect 26516 13268 26568 13320
rect 29552 13268 29604 13320
rect 30288 13268 30340 13320
rect 30932 13311 30984 13320
rect 30932 13277 30966 13311
rect 30966 13277 30984 13311
rect 30932 13268 30984 13277
rect 31208 13268 31260 13320
rect 37004 13311 37056 13320
rect 37004 13277 37008 13311
rect 37008 13277 37042 13311
rect 37042 13277 37056 13311
rect 37004 13268 37056 13277
rect 37188 13311 37240 13320
rect 37188 13277 37197 13311
rect 37197 13277 37231 13311
rect 37231 13277 37240 13311
rect 37188 13268 37240 13277
rect 38108 13311 38160 13320
rect 26056 13200 26108 13252
rect 29644 13200 29696 13252
rect 34244 13200 34296 13252
rect 35992 13200 36044 13252
rect 38108 13277 38117 13311
rect 38117 13277 38151 13311
rect 38151 13277 38160 13311
rect 38108 13268 38160 13277
rect 19984 13132 20036 13184
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20628 13132 20680 13141
rect 22100 13132 22152 13184
rect 22560 13175 22612 13184
rect 22560 13141 22569 13175
rect 22569 13141 22603 13175
rect 22603 13141 22612 13175
rect 22560 13132 22612 13141
rect 24032 13132 24084 13184
rect 34980 13132 35032 13184
rect 36820 13175 36872 13184
rect 36820 13141 36829 13175
rect 36829 13141 36863 13175
rect 36863 13141 36872 13175
rect 36820 13132 36872 13141
rect 36912 13132 36964 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 6552 12928 6604 12980
rect 8024 12928 8076 12980
rect 11152 12928 11204 12980
rect 11704 12928 11756 12980
rect 6920 12860 6972 12912
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 3700 12835 3752 12844
rect 3700 12801 3706 12835
rect 3706 12801 3752 12835
rect 3700 12792 3752 12801
rect 7012 12792 7064 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 9864 12792 9916 12844
rect 13084 12860 13136 12912
rect 13820 12928 13872 12980
rect 14004 12928 14056 12980
rect 14280 12860 14332 12912
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 13636 12792 13688 12844
rect 15384 12792 15436 12844
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16948 12835 17000 12844
rect 3424 12724 3476 12776
rect 3792 12724 3844 12776
rect 9680 12724 9732 12776
rect 12624 12724 12676 12776
rect 16028 12724 16080 12776
rect 4068 12656 4120 12708
rect 13360 12656 13412 12708
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19800 12792 19852 12844
rect 20260 12860 20312 12912
rect 20628 12792 20680 12844
rect 22560 12860 22612 12912
rect 24768 12860 24820 12912
rect 22100 12835 22152 12844
rect 22100 12801 22134 12835
rect 22134 12801 22152 12835
rect 22100 12792 22152 12801
rect 24308 12835 24360 12844
rect 24308 12801 24342 12835
rect 24342 12801 24360 12835
rect 24308 12792 24360 12801
rect 26148 12792 26200 12844
rect 27160 12928 27212 12980
rect 30012 12971 30064 12980
rect 30012 12937 30021 12971
rect 30021 12937 30055 12971
rect 30055 12937 30064 12971
rect 30012 12928 30064 12937
rect 30472 12928 30524 12980
rect 31208 12928 31260 12980
rect 29460 12860 29512 12912
rect 28540 12792 28592 12844
rect 29092 12792 29144 12844
rect 29644 12792 29696 12844
rect 32036 12928 32088 12980
rect 38108 12928 38160 12980
rect 33508 12792 33560 12844
rect 34980 12792 35032 12844
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 18604 12724 18656 12776
rect 24032 12767 24084 12776
rect 24032 12733 24041 12767
rect 24041 12733 24075 12767
rect 24075 12733 24084 12767
rect 24032 12724 24084 12733
rect 28172 12724 28224 12776
rect 30380 12724 30432 12776
rect 34152 12767 34204 12776
rect 34152 12733 34161 12767
rect 34161 12733 34195 12767
rect 34195 12733 34204 12767
rect 34152 12724 34204 12733
rect 37188 12724 37240 12776
rect 8944 12588 8996 12640
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 17040 12656 17092 12708
rect 18880 12699 18932 12708
rect 18880 12665 18889 12699
rect 18889 12665 18923 12699
rect 18923 12665 18932 12699
rect 18880 12656 18932 12665
rect 17408 12588 17460 12640
rect 19340 12588 19392 12640
rect 20904 12588 20956 12640
rect 22468 12588 22520 12640
rect 25044 12588 25096 12640
rect 25688 12588 25740 12640
rect 29644 12588 29696 12640
rect 31392 12631 31444 12640
rect 31392 12597 31401 12631
rect 31401 12597 31435 12631
rect 31435 12597 31444 12631
rect 31392 12588 31444 12597
rect 34796 12631 34848 12640
rect 34796 12597 34805 12631
rect 34805 12597 34839 12631
rect 34839 12597 34848 12631
rect 34796 12588 34848 12597
rect 35716 12631 35768 12640
rect 35716 12597 35725 12631
rect 35725 12597 35759 12631
rect 35759 12597 35768 12631
rect 35716 12588 35768 12597
rect 38016 12631 38068 12640
rect 38016 12597 38025 12631
rect 38025 12597 38059 12631
rect 38059 12597 38068 12631
rect 38016 12588 38068 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2504 12384 2556 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 7288 12384 7340 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 9772 12384 9824 12436
rect 16488 12427 16540 12436
rect 16488 12393 16497 12427
rect 16497 12393 16531 12427
rect 16531 12393 16540 12427
rect 16488 12384 16540 12393
rect 16764 12384 16816 12436
rect 19800 12427 19852 12436
rect 19800 12393 19809 12427
rect 19809 12393 19843 12427
rect 19843 12393 19852 12427
rect 19800 12384 19852 12393
rect 20260 12384 20312 12436
rect 20720 12384 20772 12436
rect 20812 12384 20864 12436
rect 24308 12384 24360 12436
rect 24676 12384 24728 12436
rect 36912 12384 36964 12436
rect 3700 12316 3752 12368
rect 9864 12316 9916 12368
rect 7472 12248 7524 12300
rect 17500 12316 17552 12368
rect 24768 12359 24820 12368
rect 24768 12325 24777 12359
rect 24777 12325 24811 12359
rect 24811 12325 24820 12359
rect 24768 12316 24820 12325
rect 34796 12359 34848 12368
rect 34796 12325 34805 12359
rect 34805 12325 34839 12359
rect 34839 12325 34848 12359
rect 34796 12316 34848 12325
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3424 12180 3476 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 8944 12223 8996 12232
rect 3516 12112 3568 12164
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9220 12180 9272 12232
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 12992 12180 13044 12232
rect 13544 12248 13596 12300
rect 20996 12248 21048 12300
rect 16764 12180 16816 12232
rect 17776 12180 17828 12232
rect 19984 12180 20036 12232
rect 20904 12180 20956 12232
rect 22008 12180 22060 12232
rect 22284 12180 22336 12232
rect 24032 12248 24084 12300
rect 25412 12291 25464 12300
rect 25412 12257 25421 12291
rect 25421 12257 25455 12291
rect 25455 12257 25464 12291
rect 25412 12248 25464 12257
rect 24400 12180 24452 12232
rect 15108 12112 15160 12164
rect 25320 12180 25372 12232
rect 25688 12223 25740 12232
rect 25688 12189 25722 12223
rect 25722 12189 25740 12223
rect 25688 12180 25740 12189
rect 29552 12223 29604 12232
rect 29552 12189 29561 12223
rect 29561 12189 29595 12223
rect 29595 12189 29604 12223
rect 29552 12180 29604 12189
rect 29644 12180 29696 12232
rect 34060 12180 34112 12232
rect 34428 12180 34480 12232
rect 36268 12180 36320 12232
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 7564 12044 7616 12096
rect 12716 12044 12768 12096
rect 26516 12112 26568 12164
rect 34244 12112 34296 12164
rect 35808 12112 35860 12164
rect 18420 12044 18472 12096
rect 18604 12087 18656 12096
rect 18604 12053 18613 12087
rect 18613 12053 18647 12087
rect 18647 12053 18656 12087
rect 18604 12044 18656 12053
rect 25320 12044 25372 12096
rect 26608 12044 26660 12096
rect 30932 12087 30984 12096
rect 30932 12053 30941 12087
rect 30941 12053 30975 12087
rect 30975 12053 30984 12087
rect 30932 12044 30984 12053
rect 34152 12087 34204 12096
rect 34152 12053 34161 12087
rect 34161 12053 34195 12087
rect 34195 12053 34204 12087
rect 34152 12044 34204 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 11336 11840 11388 11892
rect 13452 11840 13504 11892
rect 2596 11772 2648 11824
rect 7472 11704 7524 11756
rect 8944 11772 8996 11824
rect 11612 11772 11664 11824
rect 19248 11840 19300 11892
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 24400 11883 24452 11892
rect 24400 11849 24409 11883
rect 24409 11849 24443 11883
rect 24443 11849 24452 11883
rect 24400 11840 24452 11849
rect 26148 11883 26200 11892
rect 26148 11849 26157 11883
rect 26157 11849 26191 11883
rect 26191 11849 26200 11883
rect 26148 11840 26200 11849
rect 26884 11840 26936 11892
rect 28540 11883 28592 11892
rect 28540 11849 28549 11883
rect 28549 11849 28583 11883
rect 28583 11849 28592 11883
rect 28540 11840 28592 11849
rect 29092 11883 29144 11892
rect 29092 11849 29101 11883
rect 29101 11849 29135 11883
rect 29135 11849 29144 11883
rect 29092 11840 29144 11849
rect 16396 11772 16448 11824
rect 34152 11772 34204 11824
rect 9864 11704 9916 11756
rect 12624 11704 12676 11756
rect 20536 11704 20588 11756
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 22836 11704 22888 11756
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 24584 11704 24636 11713
rect 25044 11747 25096 11756
rect 17408 11636 17460 11688
rect 19340 11636 19392 11688
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 25320 11704 25372 11756
rect 25964 11747 26016 11756
rect 25136 11636 25188 11688
rect 25964 11713 25973 11747
rect 25973 11713 26007 11747
rect 26007 11713 26016 11747
rect 25964 11704 26016 11713
rect 29276 11747 29328 11756
rect 29276 11713 29285 11747
rect 29285 11713 29319 11747
rect 29319 11713 29328 11747
rect 29276 11704 29328 11713
rect 28540 11636 28592 11688
rect 1492 11611 1544 11620
rect 1492 11577 1501 11611
rect 1501 11577 1535 11611
rect 1535 11577 1544 11611
rect 1492 11568 1544 11577
rect 2872 11568 2924 11620
rect 9864 11611 9916 11620
rect 9864 11577 9873 11611
rect 9873 11577 9907 11611
rect 9907 11577 9916 11611
rect 9864 11568 9916 11577
rect 10140 11568 10192 11620
rect 18144 11568 18196 11620
rect 24768 11568 24820 11620
rect 25044 11568 25096 11620
rect 25320 11568 25372 11620
rect 2780 11500 2832 11552
rect 9220 11500 9272 11552
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 28908 11568 28960 11620
rect 30932 11704 30984 11756
rect 31024 11704 31076 11756
rect 31392 11704 31444 11756
rect 34428 11704 34480 11756
rect 32496 11568 32548 11620
rect 30472 11500 30524 11552
rect 37004 11840 37056 11892
rect 37096 11772 37148 11824
rect 37280 11747 37332 11756
rect 37280 11713 37289 11747
rect 37289 11713 37323 11747
rect 37323 11713 37332 11747
rect 37280 11704 37332 11713
rect 37372 11747 37424 11756
rect 37372 11713 37382 11747
rect 37382 11713 37416 11747
rect 37416 11713 37424 11747
rect 37372 11704 37424 11713
rect 37188 11636 37240 11688
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7380 11296 7432 11348
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2780 11092 2832 11144
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 10968 11296 11020 11348
rect 12716 11339 12768 11348
rect 9680 11024 9732 11076
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 15384 11296 15436 11348
rect 13176 11228 13228 11280
rect 15660 11228 15712 11280
rect 15844 11296 15896 11348
rect 16396 11296 16448 11348
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 17132 11296 17184 11348
rect 25412 11296 25464 11348
rect 29276 11296 29328 11348
rect 31760 11296 31812 11348
rect 33048 11296 33100 11348
rect 37372 11296 37424 11348
rect 38016 11339 38068 11348
rect 38016 11305 38025 11339
rect 38025 11305 38059 11339
rect 38059 11305 38068 11339
rect 38016 11296 38068 11305
rect 25596 11271 25648 11280
rect 11612 11092 11664 11144
rect 12440 11024 12492 11076
rect 14188 11092 14240 11144
rect 15200 11160 15252 11212
rect 17408 11160 17460 11212
rect 25320 11160 25372 11212
rect 25596 11237 25605 11271
rect 25605 11237 25639 11271
rect 25639 11237 25648 11271
rect 25596 11228 25648 11237
rect 32496 11228 32548 11280
rect 36084 11228 36136 11280
rect 37188 11228 37240 11280
rect 15936 11092 15988 11144
rect 24676 11092 24728 11144
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 2688 10999 2740 11008
rect 2688 10965 2697 10999
rect 2697 10965 2731 10999
rect 2731 10965 2740 10999
rect 2688 10956 2740 10965
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 15108 10999 15160 11008
rect 15108 10965 15117 10999
rect 15117 10965 15151 10999
rect 15151 10965 15160 10999
rect 15108 10956 15160 10965
rect 15292 10956 15344 11008
rect 19064 11024 19116 11076
rect 19432 11024 19484 11076
rect 24584 11024 24636 11076
rect 25964 11092 26016 11144
rect 30380 11160 30432 11212
rect 33508 11092 33560 11144
rect 36452 11135 36504 11144
rect 36452 11101 36461 11135
rect 36461 11101 36495 11135
rect 36495 11101 36504 11135
rect 36452 11092 36504 11101
rect 37648 11092 37700 11144
rect 30564 11067 30616 11076
rect 30564 11033 30573 11067
rect 30573 11033 30607 11067
rect 30607 11033 30616 11067
rect 30564 11024 30616 11033
rect 32680 11024 32732 11076
rect 19156 10956 19208 11008
rect 30288 10956 30340 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 9588 10752 9640 10804
rect 11520 10684 11572 10736
rect 12256 10684 12308 10736
rect 12532 10684 12584 10736
rect 2596 10616 2648 10668
rect 8208 10616 8260 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 15292 10684 15344 10736
rect 16948 10752 17000 10804
rect 21180 10752 21232 10804
rect 22376 10752 22428 10804
rect 25504 10752 25556 10804
rect 37280 10752 37332 10804
rect 38292 10752 38344 10804
rect 15844 10727 15896 10736
rect 15844 10693 15853 10727
rect 15853 10693 15887 10727
rect 15887 10693 15896 10727
rect 15844 10684 15896 10693
rect 12992 10616 13044 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 15108 10616 15160 10668
rect 15568 10616 15620 10668
rect 27620 10684 27672 10736
rect 31024 10684 31076 10736
rect 17500 10616 17552 10668
rect 17960 10616 18012 10668
rect 19340 10616 19392 10668
rect 19432 10616 19484 10668
rect 19984 10616 20036 10668
rect 25412 10616 25464 10668
rect 25780 10616 25832 10668
rect 32312 10616 32364 10668
rect 12440 10548 12492 10600
rect 12624 10548 12676 10600
rect 16764 10548 16816 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 18144 10548 18196 10600
rect 22560 10548 22612 10600
rect 6920 10480 6972 10532
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 2044 10412 2096 10464
rect 2964 10412 3016 10464
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 8392 10412 8444 10464
rect 10968 10412 11020 10464
rect 12716 10412 12768 10464
rect 18512 10480 18564 10532
rect 29736 10548 29788 10600
rect 29552 10480 29604 10532
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 16856 10412 16908 10464
rect 18972 10412 19024 10464
rect 22100 10412 22152 10464
rect 22376 10412 22428 10464
rect 28172 10412 28224 10464
rect 38016 10455 38068 10464
rect 38016 10421 38025 10455
rect 38025 10421 38059 10455
rect 38059 10421 38068 10455
rect 38016 10412 38068 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2320 10208 2372 10260
rect 10784 10208 10836 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 12900 10208 12952 10260
rect 13544 10208 13596 10260
rect 13912 10208 13964 10260
rect 17500 10208 17552 10260
rect 22560 10251 22612 10260
rect 22560 10217 22569 10251
rect 22569 10217 22603 10251
rect 22603 10217 22612 10251
rect 23756 10251 23808 10260
rect 22560 10208 22612 10217
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 27620 10251 27672 10260
rect 27620 10217 27629 10251
rect 27629 10217 27663 10251
rect 27663 10217 27672 10251
rect 27620 10208 27672 10217
rect 32680 10208 32732 10260
rect 35808 10251 35860 10260
rect 35808 10217 35817 10251
rect 35817 10217 35851 10251
rect 35851 10217 35860 10251
rect 35808 10208 35860 10217
rect 36268 10251 36320 10260
rect 36268 10217 36277 10251
rect 36277 10217 36311 10251
rect 36311 10217 36320 10251
rect 36268 10208 36320 10217
rect 2596 10140 2648 10192
rect 16120 10140 16172 10192
rect 16764 10140 16816 10192
rect 19156 10140 19208 10192
rect 30288 10183 30340 10192
rect 30288 10149 30297 10183
rect 30297 10149 30331 10183
rect 30331 10149 30340 10183
rect 30288 10140 30340 10149
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 3240 10004 3292 10056
rect 8300 10072 8352 10124
rect 9404 10072 9456 10124
rect 10600 10115 10652 10124
rect 10600 10081 10609 10115
rect 10609 10081 10643 10115
rect 10643 10081 10652 10115
rect 10600 10072 10652 10081
rect 12440 10072 12492 10124
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 9772 10004 9824 10056
rect 11060 10004 11112 10056
rect 9220 9936 9272 9988
rect 11520 9936 11572 9988
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 7288 9868 7340 9920
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 11704 9868 11756 9920
rect 15200 10072 15252 10124
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 16488 10004 16540 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 17960 10072 18012 10124
rect 18512 10115 18564 10124
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 25504 10115 25556 10124
rect 25504 10081 25513 10115
rect 25513 10081 25547 10115
rect 25547 10081 25556 10115
rect 25504 10072 25556 10081
rect 18236 10047 18288 10056
rect 13912 9936 13964 9988
rect 17316 9936 17368 9988
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 20076 10004 20128 10056
rect 20536 10004 20588 10056
rect 23756 10004 23808 10056
rect 25780 10047 25832 10056
rect 25504 9936 25556 9988
rect 25780 10013 25789 10047
rect 25789 10013 25823 10047
rect 25823 10013 25832 10047
rect 25780 10004 25832 10013
rect 30564 10072 30616 10124
rect 36636 10072 36688 10124
rect 29552 10004 29604 10056
rect 37740 10004 37792 10056
rect 26976 9936 27028 9988
rect 27712 9936 27764 9988
rect 30012 9979 30064 9988
rect 30012 9945 30021 9979
rect 30021 9945 30055 9979
rect 30055 9945 30064 9979
rect 30012 9936 30064 9945
rect 30840 9936 30892 9988
rect 17868 9868 17920 9920
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 22100 9911 22152 9920
rect 22100 9877 22109 9911
rect 22109 9877 22143 9911
rect 22143 9877 22152 9911
rect 22100 9868 22152 9877
rect 22376 9868 22428 9920
rect 22928 9868 22980 9920
rect 24584 9911 24636 9920
rect 24584 9877 24593 9911
rect 24593 9877 24627 9911
rect 24627 9877 24636 9911
rect 24584 9868 24636 9877
rect 26148 9868 26200 9920
rect 30656 9868 30708 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3884 9664 3936 9716
rect 8024 9664 8076 9716
rect 2780 9596 2832 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2872 9528 2924 9580
rect 4988 9528 5040 9580
rect 8300 9596 8352 9648
rect 11520 9664 11572 9716
rect 11796 9664 11848 9716
rect 17408 9664 17460 9716
rect 17868 9664 17920 9716
rect 18880 9664 18932 9716
rect 22376 9707 22428 9716
rect 22376 9673 22385 9707
rect 22385 9673 22419 9707
rect 22419 9673 22428 9707
rect 22376 9664 22428 9673
rect 23756 9664 23808 9716
rect 26976 9707 27028 9716
rect 26976 9673 26985 9707
rect 26985 9673 27019 9707
rect 27019 9673 27028 9707
rect 26976 9664 27028 9673
rect 30840 9707 30892 9716
rect 30840 9673 30849 9707
rect 30849 9673 30883 9707
rect 30883 9673 30892 9707
rect 30840 9664 30892 9673
rect 10876 9596 10928 9648
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 7012 9528 7064 9580
rect 8024 9528 8076 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 9404 9528 9456 9580
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2504 9324 2556 9376
rect 5264 9392 5316 9444
rect 9772 9528 9824 9580
rect 9864 9528 9916 9580
rect 11980 9528 12032 9580
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13544 9596 13596 9648
rect 18052 9596 18104 9648
rect 19340 9596 19392 9648
rect 13176 9528 13228 9537
rect 19248 9528 19300 9580
rect 19524 9528 19576 9580
rect 20076 9528 20128 9580
rect 20628 9596 20680 9648
rect 12256 9460 12308 9469
rect 13636 9460 13688 9512
rect 17132 9460 17184 9512
rect 19156 9460 19208 9512
rect 12164 9435 12216 9444
rect 12164 9401 12173 9435
rect 12173 9401 12207 9435
rect 12207 9401 12216 9435
rect 12164 9392 12216 9401
rect 3792 9324 3844 9376
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 5448 9324 5500 9376
rect 7380 9324 7432 9376
rect 8300 9324 8352 9376
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 12072 9324 12124 9376
rect 12256 9324 12308 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13360 9392 13412 9444
rect 20444 9392 20496 9444
rect 22560 9596 22612 9648
rect 23020 9596 23072 9648
rect 23296 9596 23348 9648
rect 22744 9528 22796 9580
rect 23388 9571 23440 9580
rect 23388 9537 23397 9571
rect 23397 9537 23431 9571
rect 23431 9537 23440 9571
rect 23388 9528 23440 9537
rect 24492 9528 24544 9580
rect 25412 9528 25464 9580
rect 25596 9528 25648 9580
rect 27252 9596 27304 9648
rect 31300 9596 31352 9648
rect 32588 9596 32640 9648
rect 28632 9528 28684 9580
rect 30656 9571 30708 9580
rect 30656 9537 30665 9571
rect 30665 9537 30699 9571
rect 30699 9537 30708 9571
rect 30656 9528 30708 9537
rect 31760 9528 31812 9580
rect 34612 9528 34664 9580
rect 35808 9528 35860 9580
rect 37280 9571 37332 9580
rect 37280 9537 37289 9571
rect 37289 9537 37323 9571
rect 37323 9537 37332 9571
rect 37280 9528 37332 9537
rect 22284 9460 22336 9512
rect 37556 9503 37608 9512
rect 37556 9469 37565 9503
rect 37565 9469 37599 9503
rect 37599 9469 37608 9503
rect 37556 9460 37608 9469
rect 37372 9392 37424 9444
rect 15200 9324 15252 9376
rect 17776 9324 17828 9376
rect 19064 9324 19116 9376
rect 19340 9324 19392 9376
rect 22008 9324 22060 9376
rect 22100 9324 22152 9376
rect 25504 9324 25556 9376
rect 26056 9324 26108 9376
rect 30288 9324 30340 9376
rect 34520 9324 34572 9376
rect 35440 9324 35492 9376
rect 38016 9324 38068 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2320 9120 2372 9172
rect 3700 9120 3752 9172
rect 1584 9052 1636 9104
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 7012 9120 7064 9172
rect 7380 9120 7432 9172
rect 22376 9120 22428 9172
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 25596 9120 25648 9172
rect 12072 9052 12124 9104
rect 12164 9095 12216 9104
rect 12164 9061 12173 9095
rect 12173 9061 12207 9095
rect 12207 9061 12216 9095
rect 12164 9052 12216 9061
rect 12532 9052 12584 9104
rect 13268 9052 13320 9104
rect 18236 9052 18288 9104
rect 19248 9095 19300 9104
rect 19248 9061 19257 9095
rect 19257 9061 19291 9095
rect 19291 9061 19300 9095
rect 19248 9052 19300 9061
rect 20444 9095 20496 9104
rect 20444 9061 20453 9095
rect 20453 9061 20487 9095
rect 20487 9061 20496 9095
rect 20444 9052 20496 9061
rect 22008 9052 22060 9104
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 12256 9027 12308 9036
rect 12256 8993 12265 9027
rect 12265 8993 12299 9027
rect 12299 8993 12308 9027
rect 12256 8984 12308 8993
rect 14740 8984 14792 9036
rect 3792 8916 3844 8925
rect 2780 8780 2832 8832
rect 4068 8891 4120 8900
rect 4068 8857 4102 8891
rect 4102 8857 4120 8891
rect 9588 8916 9640 8968
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 11980 8916 12032 8968
rect 4068 8848 4120 8857
rect 7104 8848 7156 8900
rect 4804 8780 4856 8832
rect 9864 8848 9916 8900
rect 11336 8848 11388 8900
rect 11704 8848 11756 8900
rect 13360 8916 13412 8968
rect 16856 8959 16908 8968
rect 16856 8925 16874 8959
rect 16874 8925 16908 8959
rect 17132 8959 17184 8968
rect 16856 8916 16908 8925
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 17868 8916 17920 8968
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 19524 8916 19576 8968
rect 22468 8984 22520 9036
rect 20076 8916 20128 8968
rect 21916 8916 21968 8968
rect 22100 8916 22152 8968
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 25136 9052 25188 9104
rect 32128 9120 32180 9172
rect 37464 9120 37516 9172
rect 34704 9052 34756 9104
rect 24584 8984 24636 9036
rect 7748 8780 7800 8832
rect 8208 8780 8260 8832
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 11796 8780 11848 8832
rect 11980 8780 12032 8832
rect 16396 8780 16448 8832
rect 16948 8780 17000 8832
rect 17224 8848 17276 8900
rect 23480 8916 23532 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 31760 8984 31812 9036
rect 25596 8916 25648 8968
rect 25964 8959 26016 8968
rect 25964 8925 25973 8959
rect 25973 8925 26007 8959
rect 26007 8925 26016 8959
rect 25964 8916 26016 8925
rect 30656 8959 30708 8968
rect 20628 8780 20680 8832
rect 21824 8823 21876 8832
rect 21824 8789 21833 8823
rect 21833 8789 21867 8823
rect 21867 8789 21876 8823
rect 21824 8780 21876 8789
rect 25228 8848 25280 8900
rect 26148 8848 26200 8900
rect 30656 8925 30665 8959
rect 30665 8925 30699 8959
rect 30699 8925 30708 8959
rect 30656 8916 30708 8925
rect 28632 8848 28684 8900
rect 32128 8916 32180 8968
rect 34336 8916 34388 8968
rect 36176 8916 36228 8968
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 36360 8891 36412 8900
rect 36360 8857 36394 8891
rect 36394 8857 36412 8891
rect 36360 8848 36412 8857
rect 27252 8780 27304 8832
rect 27988 8823 28040 8832
rect 27988 8789 27997 8823
rect 27997 8789 28031 8823
rect 28031 8789 28040 8823
rect 27988 8780 28040 8789
rect 29736 8823 29788 8832
rect 29736 8789 29745 8823
rect 29745 8789 29779 8823
rect 29779 8789 29788 8823
rect 29736 8780 29788 8789
rect 31024 8780 31076 8832
rect 31760 8780 31812 8832
rect 35808 8780 35860 8832
rect 37648 8780 37700 8832
rect 37924 8823 37976 8832
rect 37924 8789 37933 8823
rect 37933 8789 37967 8823
rect 37967 8789 37976 8823
rect 37924 8780 37976 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1492 8619 1544 8628
rect 1492 8585 1501 8619
rect 1501 8585 1535 8619
rect 1535 8585 1544 8619
rect 1492 8576 1544 8585
rect 5356 8576 5408 8628
rect 5448 8576 5500 8628
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8484 8576 8536 8628
rect 25780 8619 25832 8628
rect 2596 8440 2648 8492
rect 3792 8508 3844 8560
rect 3332 8440 3384 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 5356 8440 5408 8492
rect 5264 8372 5316 8424
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8300 8440 8352 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 10232 8508 10284 8560
rect 11980 8508 12032 8560
rect 12256 8551 12308 8560
rect 12256 8517 12265 8551
rect 12265 8517 12299 8551
rect 12299 8517 12308 8551
rect 12256 8508 12308 8517
rect 12440 8508 12492 8560
rect 17132 8508 17184 8560
rect 8392 8440 8444 8449
rect 11060 8440 11112 8492
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12900 8440 12952 8492
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 21548 8508 21600 8560
rect 21916 8551 21968 8560
rect 21916 8517 21925 8551
rect 21925 8517 21959 8551
rect 21959 8517 21968 8551
rect 21916 8508 21968 8517
rect 22008 8508 22060 8560
rect 19064 8483 19116 8492
rect 19064 8449 19098 8483
rect 19098 8449 19116 8483
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 13268 8415 13320 8424
rect 8484 8372 8536 8381
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 1584 8304 1636 8356
rect 7012 8304 7064 8356
rect 10232 8304 10284 8356
rect 3608 8236 3660 8288
rect 11060 8236 11112 8288
rect 12808 8304 12860 8356
rect 12992 8304 13044 8356
rect 13544 8347 13596 8356
rect 13544 8313 13553 8347
rect 13553 8313 13587 8347
rect 13587 8313 13596 8347
rect 13544 8304 13596 8313
rect 19064 8440 19116 8449
rect 23388 8508 23440 8560
rect 25780 8585 25789 8619
rect 25789 8585 25823 8619
rect 25823 8585 25832 8619
rect 25780 8576 25832 8585
rect 27252 8576 27304 8628
rect 29736 8576 29788 8628
rect 34060 8576 34112 8628
rect 36728 8619 36780 8628
rect 36728 8585 36737 8619
rect 36737 8585 36771 8619
rect 36771 8585 36780 8619
rect 36728 8576 36780 8585
rect 37372 8619 37424 8628
rect 37372 8585 37381 8619
rect 37381 8585 37415 8619
rect 37415 8585 37424 8619
rect 37372 8576 37424 8585
rect 32312 8508 32364 8560
rect 36176 8508 36228 8560
rect 37740 8551 37792 8560
rect 37740 8517 37749 8551
rect 37749 8517 37783 8551
rect 37783 8517 37792 8551
rect 37740 8508 37792 8517
rect 20076 8304 20128 8356
rect 22100 8304 22152 8356
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 25228 8440 25280 8492
rect 25596 8483 25648 8492
rect 25596 8449 25605 8483
rect 25605 8449 25639 8483
rect 25639 8449 25648 8483
rect 25596 8440 25648 8449
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 35348 8483 35400 8492
rect 22560 8372 22612 8424
rect 22928 8304 22980 8356
rect 21548 8236 21600 8288
rect 24860 8372 24912 8424
rect 27436 8372 27488 8424
rect 27988 8372 28040 8424
rect 30012 8372 30064 8424
rect 30288 8372 30340 8424
rect 34428 8372 34480 8424
rect 23388 8236 23440 8288
rect 25964 8304 26016 8356
rect 29552 8304 29604 8356
rect 33600 8347 33652 8356
rect 33600 8313 33609 8347
rect 33609 8313 33643 8347
rect 33643 8313 33652 8347
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35440 8440 35492 8492
rect 37556 8483 37608 8492
rect 37556 8449 37560 8483
rect 37560 8449 37594 8483
rect 37594 8449 37608 8483
rect 37556 8440 37608 8449
rect 37648 8483 37700 8492
rect 37648 8449 37657 8483
rect 37657 8449 37691 8483
rect 37691 8449 37700 8483
rect 37924 8483 37976 8492
rect 37648 8440 37700 8449
rect 37924 8449 37932 8483
rect 37932 8449 37966 8483
rect 37966 8449 37976 8483
rect 37924 8440 37976 8449
rect 38016 8483 38068 8492
rect 38016 8449 38025 8483
rect 38025 8449 38059 8483
rect 38059 8449 38068 8483
rect 38016 8440 38068 8449
rect 33600 8304 33652 8313
rect 30104 8236 30156 8288
rect 34796 8236 34848 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2872 8032 2924 8084
rect 11060 8032 11112 8084
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 13084 8075 13136 8084
rect 13084 8041 13093 8075
rect 13093 8041 13127 8075
rect 13127 8041 13136 8075
rect 13084 8032 13136 8041
rect 17408 8032 17460 8084
rect 4620 7964 4672 8016
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 4988 7896 5040 7948
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 1768 7692 1820 7744
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5264 7828 5316 7880
rect 5448 7964 5500 8016
rect 5448 7828 5500 7880
rect 11520 7828 11572 7880
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 21456 7896 21508 7948
rect 27988 8007 28040 8016
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 25964 7939 26016 7948
rect 25964 7905 25973 7939
rect 25973 7905 26007 7939
rect 26007 7905 26016 7939
rect 25964 7896 26016 7905
rect 26056 7828 26108 7880
rect 27988 7973 27997 8007
rect 27997 7973 28031 8007
rect 28031 7973 28040 8007
rect 27988 7964 28040 7973
rect 28632 8007 28684 8016
rect 28632 7973 28641 8007
rect 28641 7973 28675 8007
rect 28675 7973 28684 8007
rect 28632 7964 28684 7973
rect 30104 8007 30156 8016
rect 30104 7973 30113 8007
rect 30113 7973 30147 8007
rect 30147 7973 30156 8007
rect 30104 7964 30156 7973
rect 30656 7964 30708 8016
rect 32312 8007 32364 8016
rect 32312 7973 32321 8007
rect 32321 7973 32355 8007
rect 32355 7973 32364 8007
rect 32312 7964 32364 7973
rect 32772 8032 32824 8084
rect 35348 8032 35400 8084
rect 36360 8032 36412 8084
rect 38016 8075 38068 8084
rect 38016 8041 38025 8075
rect 38025 8041 38059 8075
rect 38059 8041 38068 8075
rect 38016 8032 38068 8041
rect 38936 7964 38988 8016
rect 7840 7760 7892 7812
rect 18972 7760 19024 7812
rect 21824 7803 21876 7812
rect 21824 7769 21858 7803
rect 21858 7769 21876 7803
rect 21824 7760 21876 7769
rect 30012 7896 30064 7948
rect 34060 7939 34112 7948
rect 34060 7905 34069 7939
rect 34069 7905 34103 7939
rect 34103 7905 34112 7939
rect 34060 7896 34112 7905
rect 30840 7828 30892 7880
rect 31024 7828 31076 7880
rect 4436 7692 4488 7744
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 8484 7692 8536 7744
rect 19984 7692 20036 7744
rect 34520 7760 34572 7812
rect 38108 7896 38160 7948
rect 35808 7828 35860 7880
rect 36728 7828 36780 7880
rect 37188 7828 37240 7880
rect 22560 7692 22612 7744
rect 27436 7692 27488 7744
rect 34704 7735 34756 7744
rect 34704 7701 34713 7735
rect 34713 7701 34747 7735
rect 34747 7701 34756 7735
rect 34704 7692 34756 7701
rect 37648 7692 37700 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3332 7531 3384 7540
rect 3332 7497 3341 7531
rect 3341 7497 3375 7531
rect 3375 7497 3384 7531
rect 3332 7488 3384 7497
rect 4068 7488 4120 7540
rect 4528 7488 4580 7540
rect 7932 7488 7984 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 3608 7352 3660 7404
rect 4068 7352 4120 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 7472 7352 7524 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 19340 7488 19392 7540
rect 22928 7488 22980 7540
rect 33600 7488 33652 7540
rect 34612 7488 34664 7540
rect 35348 7531 35400 7540
rect 35348 7497 35357 7531
rect 35357 7497 35391 7531
rect 35391 7497 35400 7531
rect 35348 7488 35400 7497
rect 35808 7488 35860 7540
rect 36084 7488 36136 7540
rect 4804 7284 4856 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8392 7284 8444 7336
rect 4528 7216 4580 7268
rect 7564 7216 7616 7268
rect 30288 7420 30340 7472
rect 34336 7420 34388 7472
rect 37188 7420 37240 7472
rect 37740 7463 37792 7472
rect 37740 7429 37749 7463
rect 37749 7429 37783 7463
rect 37783 7429 37792 7463
rect 37740 7420 37792 7429
rect 15384 7352 15436 7404
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 17408 7352 17460 7404
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 19248 7327 19300 7336
rect 19248 7293 19257 7327
rect 19257 7293 19291 7327
rect 19291 7293 19300 7327
rect 19248 7284 19300 7293
rect 27804 7352 27856 7404
rect 30288 7327 30340 7336
rect 30288 7293 30297 7327
rect 30297 7293 30331 7327
rect 30331 7293 30340 7327
rect 30288 7284 30340 7293
rect 30472 7352 30524 7404
rect 37556 7395 37608 7404
rect 37556 7361 37560 7395
rect 37560 7361 37594 7395
rect 37594 7361 37608 7395
rect 37556 7352 37608 7361
rect 36636 7284 36688 7336
rect 38016 7395 38068 7404
rect 38016 7361 38025 7395
rect 38025 7361 38059 7395
rect 38059 7361 38068 7395
rect 38016 7352 38068 7361
rect 16764 7216 16816 7268
rect 34796 7259 34848 7268
rect 34796 7225 34805 7259
rect 34805 7225 34839 7259
rect 34839 7225 34848 7259
rect 34796 7216 34848 7225
rect 37372 7259 37424 7268
rect 37372 7225 37381 7259
rect 37381 7225 37415 7259
rect 37415 7225 37424 7259
rect 37372 7216 37424 7225
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 3148 7148 3200 7200
rect 4620 7148 4672 7200
rect 4896 7148 4948 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 7288 7148 7340 7200
rect 12900 7148 12952 7200
rect 13636 7148 13688 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 16488 7148 16540 7200
rect 27528 7191 27580 7200
rect 27528 7157 27537 7191
rect 27537 7157 27571 7191
rect 27571 7157 27580 7191
rect 27528 7148 27580 7157
rect 30104 7148 30156 7200
rect 31116 7148 31168 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3884 6944 3936 6996
rect 4896 6944 4948 6996
rect 11704 6944 11756 6996
rect 15844 6944 15896 6996
rect 16856 6944 16908 6996
rect 30840 6944 30892 6996
rect 32772 6987 32824 6996
rect 32772 6953 32781 6987
rect 32781 6953 32815 6987
rect 32815 6953 32824 6987
rect 32772 6944 32824 6953
rect 36636 6987 36688 6996
rect 36636 6953 36645 6987
rect 36645 6953 36679 6987
rect 36679 6953 36688 6987
rect 36636 6944 36688 6953
rect 38016 6987 38068 6996
rect 38016 6953 38025 6987
rect 38025 6953 38059 6987
rect 38059 6953 38068 6987
rect 38016 6944 38068 6953
rect 3976 6808 4028 6860
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 11428 6808 11480 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2044 6740 2096 6792
rect 7288 6783 7340 6792
rect 7288 6749 7322 6783
rect 7322 6749 7340 6783
rect 7288 6740 7340 6749
rect 11980 6808 12032 6860
rect 27528 6876 27580 6928
rect 30104 6919 30156 6928
rect 30104 6885 30113 6919
rect 30113 6885 30147 6919
rect 30147 6885 30156 6919
rect 30104 6876 30156 6885
rect 12808 6851 12860 6860
rect 2872 6672 2924 6724
rect 5540 6672 5592 6724
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2412 6604 2464 6656
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4712 6604 4764 6656
rect 8576 6604 8628 6656
rect 11244 6672 11296 6724
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 12532 6740 12584 6792
rect 16304 6740 16356 6792
rect 19248 6808 19300 6860
rect 23296 6851 23348 6860
rect 17500 6783 17552 6792
rect 15752 6672 15804 6724
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 14464 6604 14516 6656
rect 16856 6604 16908 6656
rect 18420 6740 18472 6792
rect 21824 6740 21876 6792
rect 17776 6672 17828 6724
rect 23296 6817 23305 6851
rect 23305 6817 23339 6851
rect 23339 6817 23348 6851
rect 23296 6808 23348 6817
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 25320 6808 25372 6860
rect 26056 6808 26108 6860
rect 29092 6808 29144 6860
rect 30012 6808 30064 6860
rect 30472 6808 30524 6860
rect 30840 6851 30892 6860
rect 30840 6817 30849 6851
rect 30849 6817 30883 6851
rect 30883 6817 30892 6851
rect 30840 6808 30892 6817
rect 31116 6783 31168 6792
rect 31116 6749 31150 6783
rect 31150 6749 31168 6783
rect 31116 6740 31168 6749
rect 36452 6783 36504 6792
rect 36452 6749 36461 6783
rect 36461 6749 36495 6783
rect 36495 6749 36504 6783
rect 36452 6740 36504 6749
rect 37096 6783 37148 6792
rect 37096 6749 37105 6783
rect 37105 6749 37139 6783
rect 37139 6749 37148 6783
rect 37096 6740 37148 6749
rect 30288 6672 30340 6724
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 37280 6647 37332 6656
rect 37280 6613 37289 6647
rect 37289 6613 37323 6647
rect 37323 6613 37332 6647
rect 37280 6604 37332 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 7564 6400 7616 6452
rect 7656 6400 7708 6452
rect 12164 6400 12216 6452
rect 36820 6400 36872 6452
rect 1860 6375 1912 6384
rect 1860 6341 1869 6375
rect 1869 6341 1903 6375
rect 1903 6341 1912 6375
rect 1860 6332 1912 6341
rect 5724 6332 5776 6384
rect 7104 6332 7156 6384
rect 2872 6307 2924 6316
rect 2872 6273 2881 6307
rect 2881 6273 2915 6307
rect 2915 6273 2924 6307
rect 2872 6264 2924 6273
rect 4160 6264 4212 6316
rect 4804 6264 4856 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 9588 6264 9640 6316
rect 10784 6264 10836 6316
rect 12716 6264 12768 6316
rect 15660 6332 15712 6384
rect 19340 6332 19392 6384
rect 20536 6332 20588 6384
rect 23112 6375 23164 6384
rect 23112 6341 23121 6375
rect 23121 6341 23155 6375
rect 23155 6341 23164 6375
rect 23112 6332 23164 6341
rect 1676 6196 1728 6248
rect 11704 6196 11756 6248
rect 16580 6264 16632 6316
rect 17132 6264 17184 6316
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 3700 6128 3752 6180
rect 11152 6128 11204 6180
rect 15108 6128 15160 6180
rect 22468 6196 22520 6248
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 24584 6332 24636 6384
rect 23388 6264 23440 6273
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 34796 6264 34848 6316
rect 34704 6196 34756 6248
rect 29000 6128 29052 6180
rect 34520 6171 34572 6180
rect 34520 6137 34529 6171
rect 34529 6137 34563 6171
rect 34563 6137 34572 6171
rect 34520 6128 34572 6137
rect 37188 6128 37240 6180
rect 38108 6128 38160 6180
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3240 6060 3292 6112
rect 4068 6060 4120 6112
rect 4620 6060 4672 6112
rect 4804 6060 4856 6112
rect 7564 6060 7616 6112
rect 8116 6060 8168 6112
rect 12532 6060 12584 6112
rect 12716 6060 12768 6112
rect 13360 6060 13412 6112
rect 15752 6060 15804 6112
rect 20352 6103 20404 6112
rect 20352 6069 20361 6103
rect 20361 6069 20395 6103
rect 20395 6069 20404 6103
rect 20352 6060 20404 6069
rect 22560 6060 22612 6112
rect 25964 6060 26016 6112
rect 26056 6060 26108 6112
rect 35624 6060 35676 6112
rect 35716 6060 35768 6112
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 7104 5856 7156 5908
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 7840 5856 7892 5908
rect 12440 5856 12492 5908
rect 2504 5788 2556 5840
rect 3424 5720 3476 5772
rect 6368 5788 6420 5840
rect 12992 5788 13044 5840
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 7472 5720 7524 5729
rect 9588 5720 9640 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 3332 5652 3384 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 10324 5652 10376 5704
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 11888 5720 11940 5772
rect 18328 5856 18380 5908
rect 20536 5856 20588 5908
rect 22192 5856 22244 5908
rect 23204 5856 23256 5908
rect 20628 5788 20680 5840
rect 16580 5763 16632 5772
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 23664 5856 23716 5908
rect 24124 5856 24176 5908
rect 25872 5856 25924 5908
rect 29000 5856 29052 5908
rect 33416 5899 33468 5908
rect 33416 5865 33425 5899
rect 33425 5865 33459 5899
rect 33459 5865 33468 5899
rect 33416 5856 33468 5865
rect 36820 5899 36872 5908
rect 36820 5865 36829 5899
rect 36829 5865 36863 5899
rect 36863 5865 36872 5899
rect 36820 5856 36872 5865
rect 23572 5788 23624 5840
rect 25136 5788 25188 5840
rect 10876 5652 10928 5661
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 12072 5695 12124 5704
rect 11152 5652 11204 5661
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 14188 5652 14240 5704
rect 16488 5652 16540 5704
rect 18236 5652 18288 5704
rect 19340 5695 19392 5704
rect 19340 5661 19349 5695
rect 19349 5661 19383 5695
rect 19383 5661 19392 5695
rect 19340 5652 19392 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2780 5516 2832 5568
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 7104 5516 7156 5568
rect 11520 5584 11572 5636
rect 12164 5627 12216 5636
rect 12164 5593 12173 5627
rect 12173 5593 12207 5627
rect 12207 5593 12216 5627
rect 19984 5652 20036 5704
rect 12164 5584 12216 5593
rect 20076 5584 20128 5636
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 20352 5516 20404 5568
rect 20628 5516 20680 5568
rect 21732 5516 21784 5568
rect 22468 5695 22520 5704
rect 22468 5661 22477 5695
rect 22477 5661 22511 5695
rect 22511 5661 22520 5695
rect 22468 5652 22520 5661
rect 22560 5695 22612 5704
rect 22560 5661 22569 5695
rect 22569 5661 22603 5695
rect 22603 5661 22612 5695
rect 22744 5695 22796 5704
rect 22560 5652 22612 5661
rect 22744 5661 22753 5695
rect 22753 5661 22787 5695
rect 22787 5661 22796 5695
rect 22744 5652 22796 5661
rect 23572 5695 23624 5704
rect 23572 5661 23581 5695
rect 23581 5661 23615 5695
rect 23615 5661 23624 5695
rect 23756 5695 23808 5704
rect 23572 5652 23624 5661
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 24860 5695 24912 5704
rect 24124 5584 24176 5636
rect 24860 5661 24869 5695
rect 24869 5661 24903 5695
rect 24903 5661 24912 5695
rect 24860 5652 24912 5661
rect 25964 5788 26016 5840
rect 32864 5788 32916 5840
rect 26424 5720 26476 5772
rect 27712 5720 27764 5772
rect 34612 5720 34664 5772
rect 26056 5652 26108 5704
rect 34520 5652 34572 5704
rect 35716 5652 35768 5704
rect 37096 5695 37148 5704
rect 37096 5661 37130 5695
rect 37130 5661 37148 5695
rect 27528 5584 27580 5636
rect 36912 5584 36964 5636
rect 34428 5516 34480 5568
rect 35440 5559 35492 5568
rect 35440 5525 35449 5559
rect 35449 5525 35483 5559
rect 35483 5525 35492 5559
rect 35440 5516 35492 5525
rect 37096 5652 37148 5661
rect 37924 5652 37976 5704
rect 38108 5695 38160 5704
rect 38108 5661 38117 5695
rect 38117 5661 38151 5695
rect 38151 5661 38160 5695
rect 38108 5652 38160 5661
rect 37740 5584 37792 5636
rect 37556 5516 37608 5568
rect 37924 5559 37976 5568
rect 37924 5525 37933 5559
rect 37933 5525 37967 5559
rect 37967 5525 37976 5559
rect 37924 5516 37976 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3792 5355 3844 5364
rect 3792 5321 3801 5355
rect 3801 5321 3835 5355
rect 3835 5321 3844 5355
rect 3792 5312 3844 5321
rect 7196 5312 7248 5364
rect 11244 5312 11296 5364
rect 2412 5244 2464 5296
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2688 5176 2740 5228
rect 3424 5219 3476 5228
rect 2596 5108 2648 5160
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5540 5176 5592 5228
rect 5632 5108 5684 5160
rect 3056 5040 3108 5092
rect 6920 5244 6972 5296
rect 7196 5176 7248 5228
rect 7380 5176 7432 5228
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 8116 5244 8168 5296
rect 12072 5287 12124 5296
rect 10324 5219 10376 5228
rect 7288 5108 7340 5160
rect 7472 5108 7524 5160
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 12072 5253 12081 5287
rect 12081 5253 12115 5287
rect 12115 5253 12124 5287
rect 12072 5244 12124 5253
rect 12716 5312 12768 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 14004 5355 14056 5364
rect 14004 5321 14013 5355
rect 14013 5321 14047 5355
rect 14047 5321 14056 5355
rect 14004 5312 14056 5321
rect 14464 5312 14516 5364
rect 19432 5312 19484 5364
rect 20628 5312 20680 5364
rect 23388 5312 23440 5364
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 26148 5312 26200 5364
rect 13268 5287 13320 5296
rect 13268 5253 13277 5287
rect 13277 5253 13311 5287
rect 13311 5253 13320 5287
rect 13268 5244 13320 5253
rect 13544 5244 13596 5296
rect 14740 5244 14792 5296
rect 15292 5287 15344 5296
rect 10416 5176 10468 5185
rect 8392 5108 8444 5160
rect 11060 5176 11112 5228
rect 11796 5151 11848 5160
rect 11796 5117 11805 5151
rect 11805 5117 11839 5151
rect 11839 5117 11848 5151
rect 11796 5108 11848 5117
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 15292 5253 15301 5287
rect 15301 5253 15335 5287
rect 15335 5253 15344 5287
rect 15292 5244 15344 5253
rect 21732 5244 21784 5296
rect 17316 5176 17368 5228
rect 18236 5219 18288 5228
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 18604 5176 18656 5228
rect 19064 5176 19116 5228
rect 19984 5176 20036 5228
rect 20628 5176 20680 5228
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20996 5219 21048 5228
rect 20812 5176 20864 5185
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 24308 5244 24360 5296
rect 24124 5219 24176 5228
rect 21088 5176 21140 5185
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 24400 5219 24452 5228
rect 20536 5108 20588 5160
rect 22376 5108 22428 5160
rect 23940 5108 23992 5160
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 24400 5176 24452 5185
rect 27712 5244 27764 5296
rect 29000 5312 29052 5364
rect 32220 5355 32272 5364
rect 32220 5321 32229 5355
rect 32229 5321 32263 5355
rect 32263 5321 32272 5355
rect 32220 5312 32272 5321
rect 32864 5355 32916 5364
rect 32864 5321 32873 5355
rect 32873 5321 32907 5355
rect 32907 5321 32916 5355
rect 32864 5312 32916 5321
rect 34336 5312 34388 5364
rect 37832 5312 37884 5364
rect 37740 5287 37792 5296
rect 37740 5253 37749 5287
rect 37749 5253 37783 5287
rect 37783 5253 37792 5287
rect 37740 5244 37792 5253
rect 24676 5108 24728 5160
rect 29092 5108 29144 5160
rect 29460 5151 29512 5160
rect 29460 5117 29469 5151
rect 29469 5117 29503 5151
rect 29503 5117 29512 5151
rect 29460 5108 29512 5117
rect 5080 4972 5132 5024
rect 6276 4972 6328 5024
rect 10968 5040 11020 5092
rect 12992 5040 13044 5092
rect 24216 5040 24268 5092
rect 27804 5040 27856 5092
rect 29184 5040 29236 5092
rect 30196 5108 30248 5160
rect 35532 5176 35584 5228
rect 34612 5151 34664 5160
rect 34612 5117 34621 5151
rect 34621 5117 34655 5151
rect 34655 5117 34664 5151
rect 34612 5108 34664 5117
rect 37556 5219 37608 5228
rect 37556 5185 37560 5219
rect 37560 5185 37594 5219
rect 37594 5185 37608 5219
rect 37556 5176 37608 5185
rect 37924 5219 37976 5228
rect 37924 5185 37932 5219
rect 37932 5185 37966 5219
rect 37966 5185 37976 5219
rect 37924 5176 37976 5185
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 23112 4972 23164 5024
rect 25688 4972 25740 5024
rect 25780 5015 25832 5024
rect 25780 4981 25789 5015
rect 25789 4981 25823 5015
rect 25823 4981 25832 5015
rect 25780 4972 25832 4981
rect 28632 4972 28684 5024
rect 35440 5083 35492 5092
rect 35440 5049 35449 5083
rect 35449 5049 35483 5083
rect 35483 5049 35492 5083
rect 35440 5040 35492 5049
rect 37372 5083 37424 5092
rect 37372 5049 37381 5083
rect 37381 5049 37415 5083
rect 37415 5049 37424 5083
rect 37372 5040 37424 5049
rect 30196 5015 30248 5024
rect 30196 4981 30205 5015
rect 30205 4981 30239 5015
rect 30239 4981 30248 5015
rect 30196 4972 30248 4981
rect 33600 4972 33652 5024
rect 36268 5015 36320 5024
rect 36268 4981 36277 5015
rect 36277 4981 36311 5015
rect 36311 4981 36320 5015
rect 36268 4972 36320 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1952 4768 2004 4820
rect 2596 4768 2648 4820
rect 3516 4768 3568 4820
rect 5632 4768 5684 4820
rect 4896 4700 4948 4752
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 3240 4564 3292 4616
rect 3608 4564 3660 4616
rect 4160 4607 4212 4616
rect 1860 4539 1912 4548
rect 1860 4505 1869 4539
rect 1869 4505 1903 4539
rect 1903 4505 1912 4539
rect 1860 4496 1912 4505
rect 3884 4496 3936 4548
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 6000 4632 6052 4684
rect 7012 4768 7064 4820
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 11060 4811 11112 4820
rect 11060 4777 11069 4811
rect 11069 4777 11103 4811
rect 11103 4777 11112 4811
rect 11060 4768 11112 4777
rect 13636 4768 13688 4820
rect 15568 4811 15620 4820
rect 13268 4700 13320 4752
rect 14280 4700 14332 4752
rect 15568 4777 15577 4811
rect 15577 4777 15611 4811
rect 15611 4777 15620 4811
rect 15568 4768 15620 4777
rect 17040 4768 17092 4820
rect 17592 4811 17644 4820
rect 17592 4777 17601 4811
rect 17601 4777 17635 4811
rect 17635 4777 17644 4811
rect 17592 4768 17644 4777
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 22652 4768 22704 4820
rect 23756 4768 23808 4820
rect 24952 4811 25004 4820
rect 24952 4777 24961 4811
rect 24961 4777 24995 4811
rect 24995 4777 25004 4811
rect 24952 4768 25004 4777
rect 26792 4811 26844 4820
rect 26792 4777 26801 4811
rect 26801 4777 26835 4811
rect 26835 4777 26844 4811
rect 26792 4768 26844 4777
rect 27436 4811 27488 4820
rect 27436 4777 27445 4811
rect 27445 4777 27479 4811
rect 27479 4777 27488 4811
rect 27436 4768 27488 4777
rect 29460 4768 29512 4820
rect 34796 4768 34848 4820
rect 37096 4768 37148 4820
rect 12624 4632 12676 4684
rect 20352 4700 20404 4752
rect 20628 4700 20680 4752
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 5448 4564 5500 4616
rect 7012 4607 7064 4616
rect 7012 4573 7046 4607
rect 7046 4573 7064 4607
rect 7012 4564 7064 4573
rect 10324 4564 10376 4616
rect 10784 4607 10836 4616
rect 7472 4496 7524 4548
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 10968 4564 11020 4616
rect 11704 4564 11756 4616
rect 10692 4496 10744 4548
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 3976 4428 4028 4480
rect 13636 4428 13688 4480
rect 13820 4428 13872 4480
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14740 4564 14792 4616
rect 15108 4564 15160 4616
rect 17224 4632 17276 4684
rect 17960 4632 18012 4684
rect 21088 4632 21140 4684
rect 23112 4700 23164 4752
rect 24584 4700 24636 4752
rect 25688 4743 25740 4752
rect 25688 4709 25697 4743
rect 25697 4709 25731 4743
rect 25731 4709 25740 4743
rect 25688 4700 25740 4709
rect 25780 4743 25832 4752
rect 25780 4709 25789 4743
rect 25789 4709 25823 4743
rect 25823 4709 25832 4743
rect 31668 4743 31720 4752
rect 25780 4700 25832 4709
rect 31668 4709 31677 4743
rect 31677 4709 31711 4743
rect 31711 4709 31720 4743
rect 31668 4700 31720 4709
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16764 4607 16816 4616
rect 14372 4496 14424 4548
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 17040 4607 17092 4616
rect 16856 4564 16908 4573
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 18052 4607 18104 4616
rect 17868 4564 17920 4573
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 17224 4496 17276 4548
rect 18236 4564 18288 4616
rect 18788 4564 18840 4616
rect 21548 4564 21600 4616
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 24032 4632 24084 4684
rect 22100 4564 22152 4573
rect 23388 4564 23440 4616
rect 23664 4607 23716 4616
rect 22836 4496 22888 4548
rect 23664 4573 23673 4607
rect 23673 4573 23707 4607
rect 23707 4573 23716 4607
rect 23664 4564 23716 4573
rect 24216 4564 24268 4616
rect 24308 4564 24360 4616
rect 24492 4607 24544 4616
rect 24492 4573 24501 4607
rect 24501 4573 24535 4607
rect 24535 4573 24544 4607
rect 24676 4607 24728 4616
rect 24492 4564 24544 4573
rect 24676 4573 24685 4607
rect 24685 4573 24719 4607
rect 24719 4573 24728 4607
rect 24676 4564 24728 4573
rect 18788 4428 18840 4480
rect 23664 4428 23716 4480
rect 29184 4632 29236 4684
rect 31300 4632 31352 4684
rect 33876 4632 33928 4684
rect 34336 4632 34388 4684
rect 34612 4632 34664 4684
rect 35900 4632 35952 4684
rect 36360 4675 36412 4684
rect 36360 4641 36369 4675
rect 36369 4641 36403 4675
rect 36403 4641 36412 4675
rect 36360 4632 36412 4641
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 26424 4607 26476 4616
rect 25872 4564 25924 4573
rect 26424 4573 26433 4607
rect 26433 4573 26467 4607
rect 26467 4573 26476 4607
rect 26424 4564 26476 4573
rect 27712 4564 27764 4616
rect 28540 4564 28592 4616
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 29552 4607 29604 4616
rect 28632 4564 28684 4573
rect 29552 4573 29561 4607
rect 29561 4573 29595 4607
rect 29595 4573 29604 4607
rect 29552 4564 29604 4573
rect 30196 4564 30248 4616
rect 33416 4564 33468 4616
rect 36268 4564 36320 4616
rect 30288 4496 30340 4548
rect 28540 4471 28592 4480
rect 28540 4437 28549 4471
rect 28549 4437 28583 4471
rect 28583 4437 28592 4471
rect 29000 4471 29052 4480
rect 28540 4428 28592 4437
rect 29000 4437 29009 4471
rect 29009 4437 29043 4471
rect 29043 4437 29052 4471
rect 29000 4428 29052 4437
rect 32128 4428 32180 4480
rect 34612 4496 34664 4548
rect 33968 4428 34020 4480
rect 34428 4428 34480 4480
rect 36084 4428 36136 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 6644 4224 6696 4276
rect 10784 4224 10836 4276
rect 10968 4224 11020 4276
rect 13544 4224 13596 4276
rect 13636 4224 13688 4276
rect 23112 4224 23164 4276
rect 24308 4224 24360 4276
rect 26424 4224 26476 4276
rect 27896 4224 27948 4276
rect 28632 4224 28684 4276
rect 31668 4224 31720 4276
rect 35532 4224 35584 4276
rect 3792 4156 3844 4208
rect 4160 4156 4212 4208
rect 2320 4088 2372 4140
rect 2504 4088 2556 4140
rect 5080 4131 5132 4140
rect 2136 4063 2188 4072
rect 2136 4029 2145 4063
rect 2145 4029 2179 4063
rect 2179 4029 2188 4063
rect 2136 4020 2188 4029
rect 1768 3952 1820 4004
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 7104 4156 7156 4208
rect 6920 4088 6972 4140
rect 7564 4156 7616 4208
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 5448 3952 5500 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2964 3884 3016 3936
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5724 3884 5776 3936
rect 7380 4020 7432 4072
rect 7840 4088 7892 4140
rect 10324 4088 10376 4140
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 11428 4088 11480 4140
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8300 3884 8352 3936
rect 8760 3884 8812 3936
rect 13820 4131 13872 4140
rect 12348 4063 12400 4072
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 15292 4088 15344 4140
rect 16672 4131 16724 4140
rect 14188 4020 14240 4072
rect 14832 4020 14884 4072
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 16764 4088 16816 4140
rect 17132 4131 17184 4140
rect 16396 4020 16448 4072
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 18972 4063 19024 4072
rect 18972 4029 18981 4063
rect 18981 4029 19015 4063
rect 19015 4029 19024 4063
rect 18972 4020 19024 4029
rect 19064 4020 19116 4072
rect 20628 4088 20680 4140
rect 22744 4088 22796 4140
rect 23388 4156 23440 4208
rect 23112 4131 23164 4140
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 23848 4131 23900 4140
rect 19984 4063 20036 4072
rect 19984 4029 19993 4063
rect 19993 4029 20027 4063
rect 20027 4029 20036 4063
rect 19984 4020 20036 4029
rect 14464 3952 14516 4004
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 21548 3952 21600 4004
rect 22560 3952 22612 4004
rect 14832 3884 14884 3936
rect 16672 3884 16724 3936
rect 16948 3884 17000 3936
rect 17684 3884 17736 3936
rect 17776 3884 17828 3936
rect 23204 3884 23256 3936
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 24032 4131 24084 4140
rect 24032 4097 24041 4131
rect 24041 4097 24075 4131
rect 24075 4097 24084 4131
rect 24032 4088 24084 4097
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 29092 4156 29144 4208
rect 29828 4156 29880 4208
rect 34428 4156 34480 4208
rect 24124 4088 24176 4097
rect 24860 4131 24912 4140
rect 24860 4097 24869 4131
rect 24869 4097 24903 4131
rect 24903 4097 24912 4131
rect 24860 4088 24912 4097
rect 25044 4131 25096 4140
rect 25044 4097 25053 4131
rect 25053 4097 25087 4131
rect 25087 4097 25096 4131
rect 25044 4088 25096 4097
rect 28908 4088 28960 4140
rect 25412 4020 25464 4072
rect 30288 4088 30340 4140
rect 32128 4131 32180 4140
rect 32128 4097 32137 4131
rect 32137 4097 32171 4131
rect 32171 4097 32180 4131
rect 32128 4088 32180 4097
rect 32772 4088 32824 4140
rect 34612 4131 34664 4140
rect 34612 4097 34646 4131
rect 34646 4097 34664 4131
rect 34612 4088 34664 4097
rect 37832 4224 37884 4276
rect 37740 4199 37792 4208
rect 37740 4165 37749 4199
rect 37749 4165 37783 4199
rect 37783 4165 37792 4199
rect 37740 4156 37792 4165
rect 37556 4131 37608 4140
rect 37556 4097 37560 4131
rect 37560 4097 37594 4131
rect 37594 4097 37608 4131
rect 37556 4088 37608 4097
rect 30104 4020 30156 4072
rect 33416 4063 33468 4072
rect 33416 4029 33425 4063
rect 33425 4029 33459 4063
rect 33459 4029 33468 4063
rect 33416 4020 33468 4029
rect 33876 4063 33928 4072
rect 33876 4029 33885 4063
rect 33885 4029 33919 4063
rect 33919 4029 33928 4063
rect 33876 4020 33928 4029
rect 36084 4020 36136 4072
rect 37832 4131 37884 4140
rect 37832 4097 37877 4131
rect 37877 4097 37884 4131
rect 37832 4088 37884 4097
rect 25136 3995 25188 4004
rect 25136 3961 25145 3995
rect 25145 3961 25179 3995
rect 25179 3961 25188 3995
rect 25136 3952 25188 3961
rect 25228 3995 25280 4004
rect 25228 3961 25237 3995
rect 25237 3961 25271 3995
rect 25271 3961 25280 3995
rect 25228 3952 25280 3961
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 29000 3952 29052 4004
rect 31208 3952 31260 4004
rect 33600 3995 33652 4004
rect 33600 3961 33609 3995
rect 33609 3961 33643 3995
rect 33643 3961 33652 3995
rect 33600 3952 33652 3961
rect 37372 3995 37424 4004
rect 37372 3961 37381 3995
rect 37381 3961 37415 3995
rect 37415 3961 37424 3995
rect 37372 3952 37424 3961
rect 29460 3927 29512 3936
rect 29460 3893 29469 3927
rect 29469 3893 29503 3927
rect 29503 3893 29512 3927
rect 29460 3884 29512 3893
rect 32312 3927 32364 3936
rect 32312 3893 32321 3927
rect 32321 3893 32355 3927
rect 32355 3893 32364 3927
rect 32312 3884 32364 3893
rect 32864 3884 32916 3936
rect 35716 3884 35768 3936
rect 36636 3927 36688 3936
rect 36636 3893 36645 3927
rect 36645 3893 36679 3927
rect 36679 3893 36688 3927
rect 36636 3884 36688 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 3424 3680 3476 3732
rect 5540 3680 5592 3732
rect 6644 3680 6696 3732
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 10416 3680 10468 3732
rect 10692 3680 10744 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 15476 3680 15528 3732
rect 16672 3723 16724 3732
rect 16672 3689 16681 3723
rect 16681 3689 16715 3723
rect 16715 3689 16724 3723
rect 16672 3680 16724 3689
rect 17040 3680 17092 3732
rect 18052 3680 18104 3732
rect 22100 3680 22152 3732
rect 23112 3680 23164 3732
rect 23664 3680 23716 3732
rect 24492 3680 24544 3732
rect 25412 3723 25464 3732
rect 25412 3689 25421 3723
rect 25421 3689 25455 3723
rect 25455 3689 25464 3723
rect 25412 3680 25464 3689
rect 29368 3680 29420 3732
rect 29828 3680 29880 3732
rect 30288 3680 30340 3732
rect 8208 3612 8260 3664
rect 10324 3612 10376 3664
rect 22560 3655 22612 3664
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 7012 3544 7064 3596
rect 2504 3476 2556 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 3056 3476 3108 3528
rect 6276 3519 6328 3528
rect 6276 3485 6310 3519
rect 6310 3485 6328 3519
rect 6276 3476 6328 3485
rect 7840 3519 7892 3528
rect 1400 3408 1452 3460
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 3884 3408 3936 3460
rect 4896 3408 4948 3460
rect 6368 3408 6420 3460
rect 4712 3340 4764 3392
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 22560 3621 22569 3655
rect 22569 3621 22603 3655
rect 22603 3621 22612 3655
rect 22560 3612 22612 3621
rect 25228 3612 25280 3664
rect 25780 3612 25832 3664
rect 9680 3476 9732 3485
rect 10324 3408 10376 3460
rect 10968 3544 11020 3596
rect 12900 3544 12952 3596
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 10784 3476 10836 3528
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 25136 3544 25188 3596
rect 12440 3408 12492 3460
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 17684 3408 17736 3460
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 18788 3476 18840 3528
rect 22376 3519 22428 3528
rect 22376 3485 22385 3519
rect 22385 3485 22419 3519
rect 22419 3485 22428 3519
rect 22376 3476 22428 3485
rect 22744 3476 22796 3528
rect 24216 3476 24268 3528
rect 10692 3340 10744 3392
rect 13176 3340 13228 3392
rect 17408 3340 17460 3392
rect 18972 3408 19024 3460
rect 25044 3476 25096 3528
rect 25228 3408 25280 3460
rect 26976 3476 27028 3528
rect 28724 3476 28776 3528
rect 18512 3340 18564 3392
rect 20628 3340 20680 3392
rect 23204 3340 23256 3392
rect 27896 3408 27948 3460
rect 26240 3340 26292 3392
rect 28816 3383 28868 3392
rect 28816 3349 28825 3383
rect 28825 3349 28859 3383
rect 28859 3349 28868 3383
rect 28816 3340 28868 3349
rect 32772 3680 32824 3732
rect 36084 3723 36136 3732
rect 36084 3689 36093 3723
rect 36093 3689 36127 3723
rect 36127 3689 36136 3723
rect 36084 3680 36136 3689
rect 36360 3680 36412 3732
rect 34152 3655 34204 3664
rect 34152 3621 34161 3655
rect 34161 3621 34195 3655
rect 34195 3621 34204 3655
rect 34152 3612 34204 3621
rect 32312 3476 32364 3528
rect 33968 3519 34020 3528
rect 33968 3485 33977 3519
rect 33977 3485 34011 3519
rect 34011 3485 34020 3519
rect 33968 3476 34020 3485
rect 31116 3408 31168 3460
rect 34152 3408 34204 3460
rect 37280 3383 37332 3392
rect 37280 3349 37289 3383
rect 37289 3349 37323 3383
rect 37323 3349 37332 3383
rect 37280 3340 37332 3349
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3148 3136 3200 3188
rect 4620 3136 4672 3188
rect 4712 3136 4764 3188
rect 1584 3068 1636 3120
rect 7012 3068 7064 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 2780 2932 2832 2984
rect 3148 2932 3200 2984
rect 1584 2864 1636 2916
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 5172 3000 5224 3052
rect 5264 3000 5316 3052
rect 5448 3000 5500 3052
rect 6644 3043 6696 3052
rect 3516 2932 3568 2941
rect 5540 2932 5592 2984
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 10508 3136 10560 3188
rect 13268 3136 13320 3188
rect 8300 3000 8352 3052
rect 8392 3000 8444 3052
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 10784 3000 10836 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 12348 3000 12400 3052
rect 17132 3136 17184 3188
rect 19340 3136 19392 3188
rect 20720 3136 20772 3188
rect 22744 3179 22796 3188
rect 22744 3145 22753 3179
rect 22753 3145 22787 3179
rect 22787 3145 22796 3179
rect 22744 3136 22796 3145
rect 24216 3179 24268 3188
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 24400 3136 24452 3188
rect 24952 3136 25004 3188
rect 13176 3043 13228 3052
rect 3608 2864 3660 2916
rect 940 2796 992 2848
rect 4988 2796 5040 2848
rect 5632 2864 5684 2916
rect 6644 2796 6696 2848
rect 8760 2864 8812 2916
rect 10692 2864 10744 2916
rect 11704 2907 11756 2916
rect 11704 2873 11713 2907
rect 11713 2873 11747 2907
rect 11747 2873 11756 2907
rect 11704 2864 11756 2873
rect 9588 2796 9640 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 10416 2796 10468 2848
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 14464 3000 14516 3052
rect 16396 3000 16448 3052
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 18972 3000 19024 3052
rect 19432 3000 19484 3052
rect 17316 2932 17368 2984
rect 19708 3000 19760 3052
rect 20996 3068 21048 3120
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 22652 3000 22704 3052
rect 25136 3136 25188 3188
rect 26976 3179 27028 3188
rect 26976 3145 26985 3179
rect 26985 3145 27019 3179
rect 27019 3145 27028 3179
rect 26976 3136 27028 3145
rect 28540 3136 28592 3188
rect 31116 3136 31168 3188
rect 31208 3136 31260 3188
rect 28816 3068 28868 3120
rect 29460 3068 29512 3120
rect 17224 2864 17276 2916
rect 18420 2864 18472 2916
rect 20536 2932 20588 2984
rect 26700 3000 26752 3052
rect 29552 3043 29604 3052
rect 29552 3009 29561 3043
rect 29561 3009 29595 3043
rect 29595 3009 29604 3043
rect 29552 3000 29604 3009
rect 32772 3000 32824 3052
rect 34796 3068 34848 3120
rect 38200 3136 38252 3188
rect 37832 3068 37884 3120
rect 24676 2932 24728 2984
rect 34704 3000 34756 3052
rect 35716 3043 35768 3052
rect 35716 3009 35725 3043
rect 35725 3009 35759 3043
rect 35759 3009 35768 3043
rect 35716 3000 35768 3009
rect 36176 3000 36228 3052
rect 15844 2796 15896 2848
rect 18512 2796 18564 2848
rect 19984 2864 20036 2916
rect 20720 2864 20772 2916
rect 24124 2864 24176 2916
rect 25228 2864 25280 2916
rect 26608 2864 26660 2916
rect 26976 2864 27028 2916
rect 26240 2839 26292 2848
rect 26240 2805 26249 2839
rect 26249 2805 26283 2839
rect 26283 2805 26292 2839
rect 26240 2796 26292 2805
rect 27804 2796 27856 2848
rect 35072 2932 35124 2984
rect 35256 2932 35308 2984
rect 37372 2975 37424 2984
rect 37372 2941 37381 2975
rect 37381 2941 37415 2975
rect 37415 2941 37424 2975
rect 37372 2932 37424 2941
rect 30748 2796 30800 2848
rect 36176 2796 36228 2848
rect 37464 2864 37516 2916
rect 39580 3000 39632 3052
rect 37648 2864 37700 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4068 2592 4120 2644
rect 5540 2592 5592 2644
rect 10876 2592 10928 2644
rect 2872 2524 2924 2576
rect 4804 2524 4856 2576
rect 296 2388 348 2440
rect 2412 2388 2464 2440
rect 2872 2388 2924 2440
rect 3884 2388 3936 2440
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7748 2388 7800 2440
rect 8024 2388 8076 2440
rect 9680 2456 9732 2508
rect 10324 2524 10376 2576
rect 14740 2592 14792 2644
rect 18604 2592 18656 2644
rect 20444 2592 20496 2644
rect 25780 2592 25832 2644
rect 26056 2592 26108 2644
rect 20536 2524 20588 2576
rect 24124 2524 24176 2576
rect 9588 2388 9640 2440
rect 10692 2388 10744 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11612 2388 11664 2440
rect 15752 2456 15804 2508
rect 16304 2456 16356 2508
rect 13636 2388 13688 2440
rect 15200 2388 15252 2440
rect 15384 2388 15436 2440
rect 16488 2388 16540 2440
rect 16948 2388 17000 2440
rect 17868 2388 17920 2440
rect 18696 2388 18748 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20720 2388 20772 2440
rect 26240 2456 26292 2508
rect 23664 2431 23716 2440
rect 3976 2320 4028 2372
rect 8392 2320 8444 2372
rect 20812 2320 20864 2372
rect 23664 2397 23673 2431
rect 23673 2397 23707 2431
rect 23707 2397 23716 2431
rect 23664 2388 23716 2397
rect 22836 2320 22888 2372
rect 25780 2388 25832 2440
rect 27712 2431 27764 2440
rect 24768 2320 24820 2372
rect 27712 2397 27721 2431
rect 27721 2397 27755 2431
rect 27755 2397 27764 2431
rect 27712 2388 27764 2397
rect 26976 2320 27028 2372
rect 29368 2388 29420 2440
rect 32128 2524 32180 2576
rect 30748 2388 30800 2440
rect 32220 2388 32272 2440
rect 32864 2431 32916 2440
rect 32864 2397 32873 2431
rect 32873 2397 32907 2431
rect 32907 2397 32916 2431
rect 32864 2388 32916 2397
rect 33508 2388 33560 2440
rect 36912 2456 36964 2508
rect 37188 2456 37240 2508
rect 35624 2431 35676 2440
rect 35624 2397 35633 2431
rect 35633 2397 35667 2431
rect 35667 2397 35676 2431
rect 35624 2388 35676 2397
rect 36084 2388 36136 2440
rect 37556 2431 37608 2440
rect 37556 2397 37565 2431
rect 37565 2397 37599 2431
rect 37599 2397 37608 2431
rect 37556 2388 37608 2397
rect 28908 2320 28960 2372
rect 2964 2252 3016 2304
rect 7012 2252 7064 2304
rect 7748 2252 7800 2304
rect 9036 2252 9088 2304
rect 11060 2252 11112 2304
rect 11796 2252 11848 2304
rect 13176 2252 13228 2304
rect 13820 2252 13872 2304
rect 15200 2252 15252 2304
rect 17224 2252 17276 2304
rect 17868 2252 17920 2304
rect 19248 2252 19300 2304
rect 19984 2252 20036 2304
rect 21272 2252 21324 2304
rect 22008 2252 22060 2304
rect 23296 2252 23348 2304
rect 24032 2252 24084 2304
rect 25320 2252 25372 2304
rect 26056 2252 26108 2304
rect 27344 2252 27396 2304
rect 28080 2252 28132 2304
rect 29460 2252 29512 2304
rect 30104 2252 30156 2304
rect 31484 2252 31536 2304
rect 33508 2252 33560 2304
rect 34152 2252 34204 2304
rect 35532 2252 35584 2304
rect 36636 2295 36688 2304
rect 36636 2261 36645 2295
rect 36645 2261 36679 2295
rect 36679 2261 36688 2295
rect 36636 2252 36688 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 20260 2048 20312 2100
rect 23664 2048 23716 2100
rect 25872 2048 25924 2100
rect 37556 2048 37608 2100
rect 20168 1980 20220 2032
rect 27712 1980 27764 2032
rect 23664 1912 23716 1964
rect 26148 1912 26200 1964
rect 27528 1912 27580 1964
rect 32864 1912 32916 1964
rect 3976 212 4028 264
rect 5724 212 5776 264
<< metal2 >>
rect 2870 39672 2926 39681
rect 2870 39607 2926 39616
rect 2778 38856 2834 38865
rect 2778 38791 2834 38800
rect 1490 37904 1546 37913
rect 1490 37839 1546 37848
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1412 37097 1440 37198
rect 1398 37088 1454 37097
rect 1398 37023 1454 37032
rect 1504 36786 1532 37839
rect 2792 37466 2820 38791
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 2884 37398 2912 39607
rect 19982 39200 20038 40000
rect 35714 39536 35770 39545
rect 35714 39471 35770 39480
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 2872 37392 2924 37398
rect 2872 37334 2924 37340
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 1492 36780 1544 36786
rect 1492 36722 1544 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 19444 36378 19472 37198
rect 19996 37126 20024 39200
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35728 37194 35756 39471
rect 38198 38856 38254 38865
rect 38198 38791 38254 38800
rect 35806 38176 35862 38185
rect 35806 38111 35862 38120
rect 35820 37262 35848 38111
rect 38106 37496 38162 37505
rect 38106 37431 38162 37440
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 35716 37188 35768 37194
rect 35716 37130 35768 37136
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 35820 36922 35848 37198
rect 35992 37120 36044 37126
rect 35992 37062 36044 37068
rect 35808 36916 35860 36922
rect 35808 36858 35860 36864
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 1400 36168 1452 36174
rect 1398 36136 1400 36145
rect 18972 36168 19024 36174
rect 1452 36136 1454 36145
rect 18972 36110 19024 36116
rect 1398 36071 1454 36080
rect 18984 35894 19012 36110
rect 32128 36100 32180 36106
rect 32128 36042 32180 36048
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 18984 35866 19196 35894
rect 1400 35488 1452 35494
rect 1400 35430 1452 35436
rect 1412 35329 1440 35430
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 1398 35320 1454 35329
rect 4214 35312 4522 35332
rect 1398 35255 1454 35264
rect 1398 34504 1454 34513
rect 1398 34439 1400 34448
rect 1452 34439 1454 34448
rect 1400 34410 1452 34416
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1412 33561 1440 33934
rect 1398 33552 1454 33561
rect 1398 33487 1454 33496
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1412 32745 1440 32846
rect 1398 32736 1454 32745
rect 1398 32671 1454 32680
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1490 31784 1546 31793
rect 1412 31385 1440 31758
rect 1490 31719 1546 31728
rect 1398 31376 1454 31385
rect 1504 31346 1532 31719
rect 1398 31311 1454 31320
rect 1492 31340 1544 31346
rect 1492 31282 1544 31288
rect 2596 31136 2648 31142
rect 2596 31078 2648 31084
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30433 1440 30670
rect 2504 30592 2556 30598
rect 2504 30534 2556 30540
rect 1398 30424 1454 30433
rect 1398 30359 1454 30368
rect 1400 30048 1452 30054
rect 1398 30016 1400 30025
rect 1452 30016 1454 30025
rect 1398 29951 1454 29960
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29209 1440 29582
rect 1584 29504 1636 29510
rect 1584 29446 1636 29452
rect 1596 29238 1624 29446
rect 1584 29232 1636 29238
rect 1398 29200 1454 29209
rect 1584 29174 1636 29180
rect 2516 29170 2544 30534
rect 1398 29135 1454 29144
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2608 29102 2636 31078
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 2596 29096 2648 29102
rect 2596 29038 2648 29044
rect 1400 29028 1452 29034
rect 1400 28970 1452 28976
rect 3516 29028 3568 29034
rect 3516 28970 3568 28976
rect 1412 28801 1440 28970
rect 1584 28960 1636 28966
rect 1584 28902 1636 28908
rect 1398 28792 1454 28801
rect 1398 28727 1454 28736
rect 1596 28218 1624 28902
rect 1584 28212 1636 28218
rect 1584 28154 1636 28160
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27849 1440 28018
rect 1398 27840 1454 27849
rect 1398 27775 1454 27784
rect 1400 27464 1452 27470
rect 1398 27432 1400 27441
rect 1452 27432 1454 27441
rect 1398 27367 1454 27376
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1412 26489 1440 26930
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 1398 26480 1454 26489
rect 1398 26415 1454 26424
rect 2228 26308 2280 26314
rect 2228 26250 2280 26256
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 26081 1532 26182
rect 1490 26072 1546 26081
rect 1490 26007 1546 26016
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 25673 1440 25842
rect 1398 25664 1454 25673
rect 1398 25599 1454 25608
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1860 24812 1912 24818
rect 1860 24754 1912 24760
rect 1490 24712 1546 24721
rect 1490 24647 1546 24656
rect 1504 24410 1532 24647
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 1872 24313 1900 24754
rect 2240 24342 2268 26250
rect 2780 25424 2832 25430
rect 2780 25366 2832 25372
rect 2688 25152 2740 25158
rect 2688 25094 2740 25100
rect 2228 24336 2280 24342
rect 1858 24304 1914 24313
rect 2228 24278 2280 24284
rect 2700 24274 2728 25094
rect 1858 24239 1914 24248
rect 2688 24268 2740 24274
rect 2688 24210 2740 24216
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2148 23905 2176 24142
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 2134 23896 2190 23905
rect 2134 23831 2190 23840
rect 2424 23730 2452 24006
rect 2412 23724 2464 23730
rect 2412 23666 2464 23672
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 1492 23520 1544 23526
rect 1490 23488 1492 23497
rect 1544 23488 1546 23497
rect 1490 23423 1546 23432
rect 1858 23080 1914 23089
rect 1858 23015 1860 23024
rect 1912 23015 1914 23024
rect 1860 22986 1912 22992
rect 2516 22778 2544 23666
rect 2792 23526 2820 25366
rect 2884 23730 2912 26726
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 2148 22545 2176 22578
rect 2134 22536 2190 22545
rect 2134 22471 2190 22480
rect 1492 22432 1544 22438
rect 1492 22374 1544 22380
rect 1504 22137 1532 22374
rect 1490 22128 1546 22137
rect 1490 22063 1546 22072
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1872 21729 1900 21898
rect 1858 21720 1914 21729
rect 1858 21655 1914 21664
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21321 1440 21490
rect 3056 21344 3108 21350
rect 1398 21312 1454 21321
rect 3056 21286 3108 21292
rect 1398 21247 1454 21256
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 1492 20800 1544 20806
rect 1490 20768 1492 20777
rect 1860 20800 1912 20806
rect 1544 20768 1546 20777
rect 1860 20742 1912 20748
rect 1490 20703 1546 20712
rect 1872 20466 1900 20742
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1872 20369 1900 20402
rect 1858 20360 1914 20369
rect 1858 20295 1914 20304
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19553 1532 19654
rect 1490 19544 1546 19553
rect 1490 19479 1546 19488
rect 1872 19378 1900 19722
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1872 19009 1900 19314
rect 1858 19000 1914 19009
rect 1858 18935 1914 18944
rect 1964 18850 1992 19654
rect 1872 18822 1992 18850
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 18601 1440 18702
rect 1398 18592 1454 18601
rect 1398 18527 1454 18536
rect 1412 18426 1440 18527
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1872 18290 1900 18822
rect 2240 18358 2268 21082
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2792 19961 2820 20402
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2778 19952 2834 19961
rect 2778 19887 2834 19896
rect 2884 19378 2912 20198
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2884 18902 2912 19314
rect 3068 19310 3096 21286
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2872 18896 2924 18902
rect 2872 18838 2924 18844
rect 2976 18698 3004 19246
rect 3068 19174 3096 19246
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18970 3096 19110
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3344 18834 3372 23462
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 3436 21894 3464 22374
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3528 18970 3556 28970
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 3620 23050 3648 23462
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 3608 23044 3660 23050
rect 3608 22986 3660 22992
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 13832 21146 13860 21558
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 13556 19854 13584 20538
rect 14292 20534 14320 21286
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1490 18184 1546 18193
rect 1490 18119 1546 18128
rect 1504 17882 1532 18119
rect 1492 17876 1544 17882
rect 1492 17818 1544 17824
rect 1872 17785 1900 18226
rect 3068 17882 3096 18702
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18290 3280 18566
rect 3344 18290 3372 18770
rect 3528 18290 3556 18906
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 1858 17776 1914 17785
rect 1858 17711 1914 17720
rect 3068 17678 3096 17818
rect 3344 17814 3372 18226
rect 3528 17882 3556 18226
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 3712 17678 3740 19450
rect 3896 19446 3924 19654
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3804 18766 3832 19110
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 2148 17377 2176 17614
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 2134 17368 2190 17377
rect 3344 17338 3372 17546
rect 3988 17338 4016 18770
rect 2134 17303 2136 17312
rect 2188 17303 2190 17312
rect 3332 17332 3384 17338
rect 2136 17274 2188 17280
rect 3332 17274 3384 17280
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4080 17202 4108 18838
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 5460 17678 5488 18566
rect 6368 17808 6420 17814
rect 6274 17776 6330 17785
rect 6368 17750 6420 17756
rect 6274 17711 6330 17720
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 1490 16824 1546 16833
rect 4214 16816 4522 16836
rect 6288 16794 6316 17711
rect 6380 17542 6408 17750
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 1490 16759 1546 16768
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 1872 16425 1900 16458
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1674 16144 1730 16153
rect 6288 16114 6316 16458
rect 1674 16079 1676 16088
rect 1728 16079 1730 16088
rect 2136 16108 2188 16114
rect 1676 16050 1728 16056
rect 2136 16050 2188 16056
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 2148 16017 2176 16050
rect 2134 16008 2190 16017
rect 2134 15943 2190 15952
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 1504 15609 1532 15846
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1872 15065 1900 15370
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 1858 15056 1914 15065
rect 1400 15020 1452 15026
rect 1858 14991 1914 15000
rect 1400 14962 1452 14968
rect 1412 14657 1440 14962
rect 1398 14648 1454 14657
rect 1398 14583 1454 14592
rect 1674 14512 1730 14521
rect 1674 14447 1730 14456
rect 1688 14414 1716 14447
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1412 13938 1440 14282
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13841 1440 13874
rect 1398 13832 1454 13841
rect 1398 13767 1454 13776
rect 1674 13424 1730 13433
rect 1674 13359 1730 13368
rect 1688 13326 1716 13359
rect 1676 13320 1728 13326
rect 2136 13320 2188 13326
rect 1676 13262 1728 13268
rect 2134 13288 2136 13297
rect 2188 13288 2190 13297
rect 2134 13223 2190 13232
rect 1492 13184 1544 13190
rect 2240 13138 2268 15098
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 1492 13126 1544 13132
rect 1504 12889 1532 13126
rect 2148 13110 2268 13138
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1872 12481 1900 12786
rect 1858 12472 1914 12481
rect 1858 12407 1914 12416
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 12073 1440 12174
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1490 11656 1546 11665
rect 1490 11591 1492 11600
rect 1544 11591 1546 11600
rect 1492 11562 1544 11568
rect 1860 11144 1912 11150
rect 1858 11112 1860 11121
rect 1912 11112 1914 11121
rect 1858 11047 1914 11056
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1504 10305 1532 10406
rect 1490 10296 1546 10305
rect 1490 10231 1546 10240
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9897 1900 9998
rect 1858 9888 1914 9897
rect 1858 9823 1914 9832
rect 2056 9586 2084 10406
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1412 8129 1440 9522
rect 1584 9376 1636 9382
rect 2056 9353 2084 9522
rect 1584 9318 1636 9324
rect 2042 9344 2098 9353
rect 1596 9110 1624 9318
rect 2042 9279 2098 9288
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1504 8634 1532 8871
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 7585 1532 7686
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 7177 1440 7346
rect 1398 7168 1454 7177
rect 1398 7103 1454 7112
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6361 1532 6598
rect 1490 6352 1546 6361
rect 1490 6287 1546 6296
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 3460 1452 3466
rect 1400 3402 1452 3408
rect 1412 3233 1440 3402
rect 1398 3224 1454 3233
rect 1398 3159 1454 3168
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 296 2440 348 2446
rect 296 2382 348 2388
rect 308 800 336 2382
rect 952 800 980 2790
rect 1504 2417 1532 5510
rect 1596 5234 1624 8298
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6254 1716 6734
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1676 5704 1728 5710
rect 1674 5672 1676 5681
rect 1728 5672 1730 5681
rect 1674 5607 1730 5616
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4185 1624 5170
rect 1582 4176 1638 4185
rect 1582 4111 1638 4120
rect 1780 4010 1808 7686
rect 2044 6792 2096 6798
rect 2042 6760 2044 6769
rect 2096 6760 2098 6769
rect 2042 6695 2098 6704
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 1872 5953 1900 6326
rect 1858 5944 1914 5953
rect 1858 5879 1914 5888
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1858 4584 1914 4593
rect 1858 4519 1860 4528
rect 1912 4519 1914 4528
rect 1860 4490 1912 4496
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3126 1624 3878
rect 1780 3738 1808 3946
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1964 3058 1992 4762
rect 2148 4078 2176 13110
rect 2332 10266 2360 14214
rect 2516 14006 2544 14758
rect 2504 14000 2556 14006
rect 2504 13942 2556 13948
rect 2608 13870 2636 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 6288 15162 6316 16050
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 12442 2544 13670
rect 2792 13530 2820 13874
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3712 12850 3740 13330
rect 4080 13326 4108 13670
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 3436 12238 3464 12718
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2608 10674 2636 11766
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 11150 2820 11494
rect 2884 11150 2912 11562
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 4128 2268 7142
rect 2332 6662 2360 9114
rect 2516 8974 2544 9318
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2608 8498 2636 10134
rect 2700 9042 2728 10950
rect 2884 10713 2912 11086
rect 2870 10704 2926 10713
rect 2870 10639 2926 10648
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9654 2820 9862
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2792 8838 2820 8871
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8537 2820 8774
rect 2778 8528 2834 8537
rect 2596 8492 2648 8498
rect 2778 8463 2834 8472
rect 2596 8434 2648 8440
rect 2884 8090 2912 9522
rect 2976 8945 3004 10406
rect 2962 8936 3018 8945
rect 2962 8871 3018 8880
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 5794 2452 6598
rect 2884 6322 2912 6666
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2332 5766 2452 5794
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2332 4298 2360 5766
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 5302 2452 5646
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2332 4270 2452 4298
rect 2320 4140 2372 4146
rect 2240 4100 2320 4128
rect 2320 4082 2372 4088
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1584 2916 1636 2922
rect 1584 2858 1636 2864
rect 1490 2408 1546 2417
rect 1490 2343 1546 2352
rect 1596 800 1624 2858
rect 2332 800 2360 4082
rect 2424 2446 2452 4270
rect 2516 4146 2544 5782
rect 2700 5234 2728 6054
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2608 4826 2636 5102
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2700 4622 2728 5170
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3534 2544 4082
rect 2792 3641 2820 5510
rect 2884 5409 2912 6258
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2870 5400 2926 5409
rect 2870 5335 2926 5344
rect 2976 5001 3004 5510
rect 3068 5098 3096 12174
rect 3528 12170 3556 12786
rect 3712 12374 3740 12786
rect 3804 12782 3832 13262
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 4080 12714 4108 13262
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4080 12442 4108 12650
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10062 3280 10406
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7206 3188 7822
rect 3344 7546 3372 8434
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3056 5092 3108 5098
rect 3056 5034 3108 5040
rect 2962 4992 3018 5001
rect 2962 4927 3018 4936
rect 3252 4729 3280 6054
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2778 3632 2834 3641
rect 2778 3567 2834 3576
rect 2976 3534 3004 3878
rect 3068 3534 3096 4014
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3160 2990 3188 3130
rect 3252 3058 3280 4558
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2792 1465 2820 2926
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2884 2446 2912 2518
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2884 1873 2912 2382
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2870 1864 2926 1873
rect 2870 1799 2926 1808
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 2976 800 3004 2246
rect 3344 1057 3372 5646
rect 3436 5234 3464 5714
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3436 3738 3464 5170
rect 3528 4826 3556 12106
rect 3712 9178 3740 12310
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3804 8974 3832 9318
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8566 3832 8910
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3896 8378 3924 9658
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3804 8350 3924 8378
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3620 7410 3648 8230
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3620 4622 3648 5170
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3712 3890 3740 6122
rect 3804 5370 3832 8350
rect 4080 7546 4108 8842
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4632 8022 4660 9318
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4816 7886 4844 8774
rect 5000 8498 5028 9522
rect 5276 9450 5304 9522
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5000 7954 5028 8434
rect 5276 8430 5304 9386
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8634 5488 9318
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5368 8498 5396 8570
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 7970 5304 8366
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5092 7942 5304 7970
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4448 7410 4476 7686
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3896 4554 3924 6938
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 5710 4016 6802
rect 4080 6118 4108 7346
rect 4540 7274 4568 7482
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4632 7206 4660 7346
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4172 6322 4200 6598
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 4250 4720 4306 4729
rect 4250 4655 4252 4664
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3804 4214 3832 4422
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3528 3862 3740 3890
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3528 2990 3556 3862
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3528 2825 3556 2926
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3514 2816 3570 2825
rect 3514 2751 3570 2760
rect 3330 1048 3386 1057
rect 3330 983 3386 992
rect 3620 800 3648 2858
rect 3896 2446 3924 3402
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3988 2378 4016 4422
rect 4080 2650 4108 4655
rect 4304 4655 4306 4664
rect 4252 4626 4304 4632
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4172 4214 4200 4558
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3194 4660 6054
rect 4724 3398 4752 6598
rect 4816 6322 4844 7278
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 7002 4936 7142
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6316 4856 6322
rect 4856 6276 4936 6304
rect 4804 6258 4856 6264
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2318 0 2374 800
rect 2962 0 3018 800
rect 3606 0 3662 800
rect 3988 649 4016 2314
rect 4356 870 4476 898
rect 4356 800 4384 870
rect 3974 640 4030 649
rect 3974 575 4030 584
rect 3976 264 4028 270
rect 3974 232 3976 241
rect 4028 232 4030 241
rect 3974 167 4030 176
rect 4342 0 4398 800
rect 4448 762 4476 870
rect 4724 762 4752 3130
rect 4816 2582 4844 6054
rect 4908 4758 4936 6276
rect 5092 5114 5120 7942
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5368 7868 5396 8434
rect 5460 8022 5488 8570
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5448 7880 5500 7886
rect 5368 7840 5448 7868
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5000 5086 5120 5114
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3466 4936 3878
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 5000 2938 5028 5086
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4146 5120 4966
rect 5184 4622 5212 5170
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5276 3058 5304 7822
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5184 2938 5212 2994
rect 5368 2938 5396 7840
rect 5448 7822 5500 7828
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 5914 5580 6666
rect 5736 6390 5764 7142
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5552 5352 5580 5850
rect 6380 5846 6408 17478
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6564 16726 6592 17274
rect 6840 17134 6868 17614
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6840 16794 6868 17070
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 6564 12986 6592 16662
rect 6932 16250 6960 17138
rect 7300 16998 7328 17614
rect 7392 17134 7420 17682
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7010 16552 7066 16561
rect 7010 16487 7012 16496
rect 7064 16487 7066 16496
rect 7012 16458 7064 16464
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6932 12918 6960 15982
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6932 10538 6960 12854
rect 7024 12850 7052 13262
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7024 9586 7052 12786
rect 7300 12442 7328 16934
rect 7392 16658 7420 17070
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7484 15706 7512 18634
rect 9324 18358 9352 19178
rect 10336 18426 10364 19790
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 7562 17640 7618 17649
rect 7562 17575 7564 17584
rect 7616 17575 7618 17584
rect 7564 17546 7616 17552
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 7748 17128 7800 17134
rect 7746 17096 7748 17105
rect 8116 17128 8168 17134
rect 7800 17096 7802 17105
rect 8116 17070 8168 17076
rect 7746 17031 7802 17040
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7944 16046 7972 16526
rect 8128 16182 8156 17070
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 8128 14006 8156 16118
rect 8312 16114 8340 16390
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8956 15706 8984 17138
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9140 15502 9168 18022
rect 9508 16590 9536 18226
rect 10060 18086 10088 18226
rect 10048 18080 10100 18086
rect 10232 18080 10284 18086
rect 10048 18022 10100 18028
rect 10152 18028 10232 18034
rect 10152 18022 10284 18028
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 14074 8340 15302
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8956 13326 8984 14010
rect 9508 13394 9536 16526
rect 9600 14090 9628 17818
rect 10060 17066 10088 18022
rect 10152 18006 10272 18022
rect 10152 17746 10180 18006
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 15910 9996 16526
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9600 14062 9720 14090
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9600 13530 9628 13874
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9692 13410 9720 14062
rect 9784 13938 9812 15642
rect 9968 15162 9996 15846
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13938 9904 14214
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9600 13382 9720 13410
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 7944 12442 7972 13194
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7288 12436 7340 12442
rect 7932 12436 7984 12442
rect 7340 12406 7604 12434
rect 7288 12378 7340 12384
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11354 7420 12038
rect 7484 11762 7512 12242
rect 7576 12102 7604 12406
rect 7932 12378 7984 12384
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 9178 7052 9522
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7024 8362 7052 9114
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7116 8634 7144 8842
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7300 8498 7328 9862
rect 8036 9722 8064 12922
rect 8128 12238 8156 13194
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12238 8984 12582
rect 9140 12238 9168 13262
rect 9416 12238 9444 13262
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8956 11830 8984 12174
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 9232 11558 9260 12174
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8220 10062 8248 10610
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9178 7420 9318
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7024 6866 7052 8298
rect 7484 7410 7512 8434
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7576 7274 7604 8366
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 5552 5324 5672 5352
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4010 5488 4558
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3058 5488 3946
rect 5552 3738 5580 5170
rect 5644 5166 5672 5324
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4826 5672 5102
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5000 2910 5120 2938
rect 5184 2910 5396 2938
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 5000 800 5028 2790
rect 5092 2774 5120 2910
rect 5092 2746 5396 2774
rect 5368 2446 5396 2746
rect 5552 2650 5580 2926
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5644 800 5672 2858
rect 4448 734 4752 762
rect 4986 0 5042 800
rect 5630 0 5686 800
rect 5736 270 5764 3878
rect 6012 3602 6040 4626
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6288 3534 6316 4966
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6656 3738 6684 4218
rect 6932 4146 6960 5238
rect 7024 4826 7052 6802
rect 7300 6798 7328 7142
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7576 6474 7604 7210
rect 7484 6458 7604 6474
rect 7668 6458 7696 7346
rect 7484 6452 7616 6458
rect 7484 6446 7564 6452
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7116 5914 7144 6326
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7116 5794 7144 5850
rect 7116 5766 7328 5794
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7012 4616 7064 4622
rect 7116 4604 7144 5510
rect 7208 5370 7236 5646
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7064 4576 7144 4604
rect 7012 4558 7064 4564
rect 7208 4298 7236 5170
rect 7300 5166 7328 5766
rect 7392 5234 7420 5850
rect 7484 5778 7512 6446
rect 7564 6394 7616 6400
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7576 5234 7604 6054
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4554 7512 5102
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7116 4270 7236 4298
rect 7116 4214 7144 4270
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7484 4146 7512 4490
rect 7576 4214 7604 5170
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7392 3738 7420 4014
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 800 6408 3402
rect 6656 3058 6684 3674
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7024 3126 7052 3538
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 7392 3058 7420 3674
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2446 6684 2790
rect 7760 2446 7788 8774
rect 8036 8634 8064 9522
rect 8220 8838 8248 9998
rect 8312 9654 8340 10066
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8312 8498 8340 9318
rect 8404 8498 8432 10406
rect 9232 9994 9260 11494
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10130 9444 10950
rect 9600 10810 9628 13382
rect 9784 12968 9812 13874
rect 9784 12940 9904 12968
rect 9876 12850 9904 12940
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 11082 9720 12718
rect 9784 12442 9812 12786
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9876 12374 9904 12786
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11626 9904 11698
rect 10152 11626 10180 17682
rect 10336 17678 10364 18362
rect 11808 18086 11836 18566
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10336 16522 10364 17614
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10704 16454 10732 17070
rect 10796 16590 10824 17478
rect 10980 17202 11008 17614
rect 11072 17202 11100 17750
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11164 17513 11192 17614
rect 11808 17542 11836 18022
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11796 17536 11848 17542
rect 11150 17504 11206 17513
rect 11796 17478 11848 17484
rect 11150 17439 11206 17448
rect 11808 17202 11836 17478
rect 12084 17338 12112 17818
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 15706 10732 16390
rect 10796 16114 10824 16526
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10888 15502 10916 15846
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 13462 10732 13670
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10704 13326 10732 13398
rect 10692 13320 10744 13326
rect 10690 13288 10692 13297
rect 10744 13288 10746 13297
rect 10690 13223 10746 13232
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10980 11354 11008 15846
rect 11072 15094 11100 17138
rect 12268 16658 12296 18022
rect 12360 17270 12388 18226
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17882 12664 18158
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12452 16726 12480 17818
rect 13188 17610 13216 18226
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12268 16114 12296 16594
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12452 16046 12480 16662
rect 12544 16590 12572 17138
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11900 15706 11928 15914
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11164 13190 11192 15302
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12986 11192 13126
rect 11716 12986 11744 13262
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9692 10690 9720 11018
rect 9600 10662 9720 10690
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 9586 9260 9930
rect 9416 9586 9444 10066
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9600 8974 9628 10662
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9586 9812 9998
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8496 8430 8524 8570
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7852 7410 7880 7754
rect 8496 7750 8524 8366
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 7944 7546 7972 7686
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 5914 7880 7346
rect 7944 7342 7972 7482
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8404 6322 8432 7278
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6322 8616 6598
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 8128 6118 8156 6258
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8128 4826 8156 5238
rect 8404 5166 8432 6258
rect 9600 5778 9628 6258
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7852 3534 7880 4082
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8128 2774 8156 4762
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8220 3670 8248 3878
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8312 3058 8340 3878
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8036 2746 8156 2774
rect 8036 2446 8064 2746
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8404 2378 8432 2994
rect 8772 2922 8800 3878
rect 9600 3058 9628 5714
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9692 3369 9720 3470
rect 9678 3360 9734 3369
rect 9678 3295 9734 3304
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9784 2938 9812 9522
rect 9876 8906 9904 9522
rect 10612 9518 10640 10066
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10796 9382 10824 10202
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9654 10916 9862
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10980 8974 11008 10406
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8566 10272 8774
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10244 8362 10272 8502
rect 11072 8498 11100 9998
rect 11348 8906 11376 11834
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11624 11150 11652 11766
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11532 9994 11560 10678
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11532 9722 11560 9930
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 8090 11100 8230
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11440 6866 11468 8774
rect 11532 7886 11560 9658
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10796 5710 10824 6258
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11164 5710 11192 6122
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10336 5234 10364 5646
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10336 4622 10364 5170
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4146 10364 4558
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10322 3904 10378 3913
rect 10322 3839 10378 3848
rect 10336 3670 10364 3839
rect 10428 3738 10456 5170
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10322 3496 10378 3505
rect 10322 3431 10324 3440
rect 10376 3431 10378 3440
rect 10324 3402 10376 3408
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 9692 2910 9812 2938
rect 10336 3040 10364 3402
rect 10520 3194 10548 4082
rect 10704 3738 10732 4490
rect 10796 4282 10824 4558
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10692 3392 10744 3398
rect 10796 3369 10824 3470
rect 10692 3334 10744 3340
rect 10782 3360 10838 3369
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10600 3052 10652 3058
rect 10336 3012 10600 3040
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9600 2446 9628 2790
rect 9692 2514 9720 2910
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7024 800 7052 2246
rect 7760 800 7788 2246
rect 8404 800 8432 2314
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 800 9076 2246
rect 9784 800 9812 2790
rect 10336 2582 10364 3012
rect 10600 2994 10652 3000
rect 10704 2922 10732 3334
rect 10782 3295 10838 3304
rect 10796 3058 10824 3295
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10428 800 10456 2790
rect 10704 2446 10732 2858
rect 10796 2446 10824 2994
rect 10888 2650 10916 5646
rect 11256 5370 11284 6666
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 4622 11008 5034
rect 11072 4826 11100 5170
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10980 4282 11008 4558
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11428 4140 11480 4146
rect 11532 4128 11560 5578
rect 11480 4100 11560 4128
rect 11428 4082 11480 4088
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10980 3505 11008 3538
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11624 2446 11652 11086
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 8906 11744 9862
rect 11808 9722 11836 13874
rect 12268 13530 12296 15370
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12268 10742 12296 11494
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11716 6254 11744 6938
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11808 5166 11836 8774
rect 11900 5778 11928 9318
rect 11992 8974 12020 9522
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9110 12112 9318
rect 12176 9110 12204 9386
rect 12268 9382 12296 9454
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12268 9042 12296 9318
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 11980 8968 12032 8974
rect 11978 8936 11980 8945
rect 12032 8936 12034 8945
rect 11978 8871 12034 8880
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 12070 8800 12126 8809
rect 11992 8566 12020 8774
rect 12070 8735 12126 8744
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 12084 8498 12112 8735
rect 12256 8560 12308 8566
rect 12176 8520 12256 8548
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11980 6860 12032 6866
rect 12176 6848 12204 8520
rect 12360 8548 12388 14282
rect 12452 14006 12480 15982
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12636 14346 12664 15914
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 13190 12572 13874
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12728 12850 12756 17138
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 15609 12848 16390
rect 12806 15600 12862 15609
rect 12806 15535 12808 15544
rect 12860 15535 12862 15544
rect 12808 15506 12860 15512
rect 12912 15434 12940 16934
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13004 15570 13032 16526
rect 13096 15706 13124 16730
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13188 15638 13216 17546
rect 13280 16658 13308 18090
rect 13372 17513 13400 18634
rect 13464 18426 13492 19790
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13740 19281 13768 19382
rect 13924 19378 13952 20334
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 13726 19272 13782 19281
rect 13726 19207 13782 19216
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13464 17610 13492 17818
rect 13556 17746 13584 18090
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13358 17504 13414 17513
rect 13358 17439 13414 17448
rect 13372 17338 13400 17439
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13464 17218 13492 17546
rect 13372 17190 13492 17218
rect 13372 16726 13400 17190
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 14822 12940 15370
rect 13004 14890 13032 15506
rect 13188 15314 13216 15574
rect 13280 15502 13308 16594
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13096 15286 13216 15314
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 13004 14414 13032 14826
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12636 11762 12664 12718
rect 12728 12102 12756 12786
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10606 12480 11018
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10130 12480 10542
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12544 9110 12572 10678
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 10146 12664 10542
rect 12728 10470 12756 11290
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10266 12756 10406
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12636 10118 12756 10146
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12308 8520 12388 8548
rect 12440 8560 12492 8566
rect 12256 8502 12308 8508
rect 12440 8502 12492 8508
rect 12032 6820 12204 6848
rect 11980 6802 12032 6808
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 12084 5710 12112 6820
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 5302 12112 5646
rect 12176 5642 12204 6394
rect 12452 5914 12480 8502
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12544 6118 12572 6734
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12254 5808 12310 5817
rect 12254 5743 12310 5752
rect 12268 5710 12296 5743
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12254 5264 12310 5273
rect 12254 5199 12256 5208
rect 12308 5199 12310 5208
rect 12256 5170 12308 5176
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 12636 4690 12664 8026
rect 12728 6322 12756 10118
rect 12820 8362 12848 10610
rect 12912 10266 12940 14214
rect 13004 13326 13032 14350
rect 13096 14346 13124 15286
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 13326 13124 14282
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13096 12918 13124 13262
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13188 12434 13216 14826
rect 13280 14006 13308 15438
rect 13372 14278 13400 16662
rect 13556 16114 13584 16934
rect 13924 16250 13952 19314
rect 14200 18426 14228 19314
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14384 18290 14412 20742
rect 14476 20058 14504 21490
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 14568 21078 14596 21286
rect 14556 21072 14608 21078
rect 14556 21014 14608 21020
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 18766 14504 19654
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14568 18698 14596 21014
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14936 20058 14964 20878
rect 15028 20618 15056 20946
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20806 15700 20878
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15028 20590 15240 20618
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14936 18766 14964 19994
rect 15212 19786 15240 20590
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15212 18766 15240 19722
rect 15672 19514 15700 20742
rect 16500 20330 16528 21286
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15948 18970 15976 19790
rect 16500 19718 16528 20266
rect 16684 20262 16712 21014
rect 16960 20398 16988 23530
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21690 17264 22034
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17144 20806 17172 20878
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16684 20058 16712 20198
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16500 19174 16528 19654
rect 16684 19446 16712 19790
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16684 19174 16712 19382
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 14568 18290 14596 18634
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14200 17882 14228 18158
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14200 17785 14228 17818
rect 14186 17776 14242 17785
rect 14186 17711 14242 17720
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14384 16182 14412 17138
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15638 14320 15846
rect 14384 15706 14412 16118
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13358 13968 13414 13977
rect 13358 13903 13360 13912
rect 13412 13903 13414 13912
rect 13360 13874 13412 13880
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13096 12406 13216 12434
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 10674 13032 12174
rect 13096 10674 13124 12406
rect 13280 11370 13308 13806
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12714 13400 13262
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13464 11898 13492 15370
rect 14384 15094 14412 15642
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14476 15026 14504 15846
rect 14568 15502 14596 17274
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 12306 13584 13874
rect 13648 12850 13676 13942
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13188 11342 13308 11370
rect 13188 11286 13216 11342
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13188 9586 13216 11222
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13556 10062 13584 10202
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9654 13584 9998
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 8498 12940 9318
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7426 12848 7822
rect 12820 7398 12940 7426
rect 12806 7304 12862 7313
rect 12806 7239 12862 7248
rect 12820 6866 12848 7239
rect 12912 7206 12940 7398
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5370 12756 6054
rect 13004 5846 13032 8298
rect 13096 8090 13124 8434
rect 13280 8430 13308 9046
rect 13372 8974 13400 9386
rect 13360 8968 13412 8974
rect 13358 8936 13360 8945
rect 13412 8936 13414 8945
rect 13358 8871 13414 8880
rect 13372 8498 13400 8871
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12898 5672 12954 5681
rect 12898 5607 12954 5616
rect 12912 5370 12940 5607
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12728 5137 12756 5306
rect 12714 5128 12770 5137
rect 13004 5098 13032 5782
rect 13268 5296 13320 5302
rect 13372 5250 13400 6054
rect 13556 5302 13584 8298
rect 13648 7206 13676 9454
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13320 5244 13400 5250
rect 13268 5238 13400 5244
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13176 5228 13228 5234
rect 13280 5222 13400 5238
rect 13176 5170 13228 5176
rect 12714 5063 12770 5072
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 13188 5001 13216 5170
rect 13174 4992 13230 5001
rect 13174 4927 13230 4936
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11716 2922 11744 4558
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 11796 3528 11848 3534
rect 11794 3496 11796 3505
rect 11848 3496 11850 3505
rect 11794 3431 11850 3440
rect 11808 3058 11836 3431
rect 12360 3058 12388 4014
rect 12898 3768 12954 3777
rect 12898 3703 12900 3712
rect 12952 3703 12954 3712
rect 12900 3674 12952 3680
rect 12912 3602 12940 3674
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11072 800 11100 2246
rect 11808 800 11836 2246
rect 12452 800 12480 3402
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 3058 13216 3334
rect 13280 3194 13308 4694
rect 13372 4049 13400 5222
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 4282 13584 5102
rect 13648 4826 13676 7142
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13648 4486 13676 4762
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13648 4282 13676 4422
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13358 4040 13414 4049
rect 13358 3975 13414 3984
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13740 2774 13768 14010
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13832 12986 13860 13466
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13924 10266 13952 14486
rect 14476 14006 14504 14554
rect 14568 14550 14596 15438
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14660 13938 14688 14350
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13924 9994 13952 10202
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 14016 5370 14044 12922
rect 14200 12646 14228 13874
rect 14752 13394 14780 14826
rect 14830 14376 14886 14385
rect 14936 14346 14964 17070
rect 15948 16726 15976 17614
rect 16316 17542 16344 18634
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 15948 16114 15976 16662
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15212 15502 15240 16050
rect 16040 15910 16068 16594
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16040 15570 16068 15846
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15026 15700 15370
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15304 14414 15332 14962
rect 16040 14958 16068 15506
rect 16132 15502 16160 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 15706 16252 16730
rect 16316 16522 16344 17478
rect 16408 16590 16436 17546
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15396 14482 15424 14894
rect 16224 14890 16252 15642
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14830 14311 14886 14320
rect 14924 14340 14976 14346
rect 14844 14006 14872 14311
rect 14924 14282 14976 14288
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12918 14320 13126
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 11150 14228 12582
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14752 9042 14780 13330
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14464 6656 14516 6662
rect 14462 6624 14464 6633
rect 14516 6624 14518 6633
rect 14462 6559 14518 6568
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4146 13860 4422
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14200 4078 14228 5646
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14280 4752 14332 4758
rect 14332 4700 14412 4706
rect 14280 4694 14412 4700
rect 14292 4678 14412 4694
rect 14384 4554 14412 4678
rect 14476 4622 14504 5306
rect 14752 5302 14780 8978
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14476 4010 14504 4558
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 13648 2746 13768 2774
rect 13648 2446 13676 2746
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13188 800 13216 2246
rect 13832 800 13860 2246
rect 14476 800 14504 2994
rect 14752 2650 14780 4558
rect 14844 4078 14872 13942
rect 15396 13870 15424 14418
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15120 12170 15148 13194
rect 15396 12850 15424 13670
rect 15488 13297 15516 14350
rect 15580 13802 15608 14554
rect 15672 14550 15700 14758
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 16040 13938 16068 14758
rect 16224 14618 16252 14826
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13938 16160 14214
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15764 13394 15792 13874
rect 16316 13818 16344 16458
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16132 13790 16344 13818
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15474 13288 15530 13297
rect 15474 13223 15530 13232
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10674 15148 10950
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15212 10130 15240 11154
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 10742 15332 10950
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 9382 15240 10066
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15396 7410 15424 11290
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15120 4622 15148 6122
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15108 4616 15160 4622
rect 15212 4593 15240 5510
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15108 4558 15160 4564
rect 15198 4584 15254 4593
rect 15198 4519 15254 4528
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14844 3942 14872 4014
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 15212 2446 15240 4519
rect 15304 4146 15332 5238
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15488 3738 15516 13223
rect 15856 12850 15884 13738
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15948 12850 15976 13330
rect 15844 12844 15896 12850
rect 15764 12804 15844 12832
rect 15764 12434 15792 12804
rect 15844 12786 15896 12792
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15672 12406 15792 12434
rect 15672 11286 15700 12406
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15856 10742 15884 11290
rect 15948 11150 15976 12786
rect 16040 12782 16068 13738
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16132 12434 16160 13790
rect 16040 12406 16160 12434
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 4826 15608 10610
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 6390 15700 7142
rect 15856 7002 15884 7346
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15764 6118 15792 6666
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15764 4604 15792 6054
rect 15844 4616 15896 4622
rect 15764 4576 15844 4604
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15488 2774 15516 3674
rect 15396 2746 15516 2774
rect 15396 2446 15424 2746
rect 15764 2514 15792 4576
rect 15844 4558 15896 4564
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 800 15240 2246
rect 15856 800 15884 2790
rect 16040 2774 16068 12406
rect 16408 11914 16436 15438
rect 16500 15366 16528 19110
rect 16684 18630 16712 19110
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16960 18426 16988 20334
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17144 18358 17172 20742
rect 17420 20602 17448 21490
rect 18788 21344 18840 21350
rect 18708 21292 18788 21298
rect 18708 21286 18840 21292
rect 18708 21270 18828 21286
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18064 20602 18092 20878
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18248 20534 18276 20742
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 17236 20058 17264 20402
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 18616 19786 18644 20402
rect 18708 19854 18736 21270
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17338 16620 17478
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 17512 17066 17540 18566
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16684 16590 16712 16730
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16776 16046 16804 16186
rect 16960 16046 16988 16594
rect 17512 16590 17540 17002
rect 18248 16658 18276 18702
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17604 16114 17632 16526
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 16114 18184 16390
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16224 11886 16436 11914
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 10198 16160 10406
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16224 4865 16252 11886
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16408 11354 16436 11766
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16500 10062 16528 12378
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 6792 16356 6798
rect 16302 6760 16304 6769
rect 16356 6760 16358 6769
rect 16302 6695 16358 6704
rect 16210 4856 16266 4865
rect 16210 4791 16266 4800
rect 16408 4078 16436 8774
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 5710 16528 7142
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16592 5778 16620 6258
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16684 4146 16712 13194
rect 16776 12442 16804 15982
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16868 15026 16896 15574
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16856 14884 16908 14890
rect 16960 14872 16988 15982
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17052 14958 17080 15574
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17328 15065 17356 15098
rect 17314 15056 17370 15065
rect 17132 15020 17184 15026
rect 17314 14991 17370 15000
rect 17132 14962 17184 14968
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16908 14844 16988 14872
rect 16856 14826 16908 14832
rect 16868 13870 16896 14826
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 17052 13433 17080 14214
rect 17144 13938 17172 14962
rect 17406 14784 17462 14793
rect 17406 14719 17462 14728
rect 17420 14346 17448 14719
rect 17408 14340 17460 14346
rect 17328 14300 17408 14328
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17236 14006 17264 14214
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17132 13456 17184 13462
rect 17038 13424 17094 13433
rect 17132 13398 17184 13404
rect 17038 13359 17094 13368
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12832 16896 13126
rect 17144 12850 17172 13398
rect 17236 13394 17264 13670
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17328 13190 17356 14300
rect 17408 14282 17460 14288
rect 17512 13802 17540 15302
rect 17684 15088 17736 15094
rect 17960 15088 18012 15094
rect 17736 15048 17908 15076
rect 17684 15030 17736 15036
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17788 14521 17816 14758
rect 17774 14512 17830 14521
rect 17774 14447 17830 14456
rect 17880 14414 17908 15048
rect 18012 15036 18092 15042
rect 17960 15030 18092 15036
rect 17972 15014 18092 15030
rect 18064 14929 18092 15014
rect 18050 14920 18106 14929
rect 17960 14884 18012 14890
rect 18050 14855 18106 14864
rect 17960 14826 18012 14832
rect 17972 14793 18000 14826
rect 18052 14816 18104 14822
rect 17958 14784 18014 14793
rect 18052 14758 18104 14764
rect 17958 14719 18014 14728
rect 18064 14618 18092 14758
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17684 14408 17736 14414
rect 17868 14408 17920 14414
rect 17684 14350 17736 14356
rect 17774 14376 17830 14385
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 16948 12844 17000 12850
rect 16868 12804 16948 12832
rect 16948 12786 17000 12792
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11354 16804 12174
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16960 10810 16988 12786
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16776 10198 16804 10542
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16776 7274 16804 10134
rect 16868 8974 16896 10406
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16960 8838 16988 9998
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16868 7002 16896 7346
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 4622 16896 6598
rect 17052 4826 17080 12650
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 11694 17448 12582
rect 17512 12374 17540 13126
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17144 10606 17172 11290
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17144 8974 17172 9454
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8566 17172 8910
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17236 8809 17264 8842
rect 17222 8800 17278 8809
rect 17222 8735 17278 8744
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 6322 17172 8502
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17328 5234 17356 9930
rect 17420 9722 17448 11154
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17420 8090 17448 9658
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17420 7410 17448 8026
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17500 6792 17552 6798
rect 17498 6760 17500 6769
rect 17552 6760 17554 6769
rect 17498 6695 17554 6704
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17236 4690 17264 4966
rect 17604 4826 17632 14282
rect 17696 14074 17724 14350
rect 17920 14356 18000 14362
rect 17868 14350 18000 14356
rect 17880 14334 18000 14350
rect 17774 14311 17776 14320
rect 17828 14311 17830 14320
rect 17776 14282 17828 14288
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 16764 4616 16816 4622
rect 16856 4616 16908 4622
rect 16764 4558 16816 4564
rect 16854 4584 16856 4593
rect 17040 4616 17092 4622
rect 16908 4584 16910 4593
rect 16776 4146 16804 4558
rect 17040 4558 17092 4564
rect 16854 4519 16910 4528
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3058 16436 4014
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16684 3738 16712 3878
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16040 2746 16344 2774
rect 16316 2514 16344 2746
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 16960 2446 16988 3878
rect 17052 3738 17080 4558
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17236 4146 17264 4490
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17144 3194 17172 4082
rect 17696 3942 17724 13874
rect 17788 12238 17816 14010
rect 17880 13870 17908 14214
rect 17972 13938 18000 14334
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17868 13864 17920 13870
rect 17866 13832 17868 13841
rect 17920 13832 17922 13841
rect 17866 13767 17922 13776
rect 17868 12776 17920 12782
rect 17866 12744 17868 12753
rect 17920 12744 17922 12753
rect 17866 12679 17922 12688
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 18156 11626 18184 16050
rect 18248 15638 18276 16594
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 18340 15348 18368 17206
rect 18432 15502 18460 17274
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18524 16153 18552 17206
rect 18616 17082 18644 19722
rect 18708 19242 18736 19790
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 17270 18828 17614
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18616 17054 18828 17082
rect 18800 16454 18828 17054
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18510 16144 18566 16153
rect 18510 16079 18566 16088
rect 18800 16046 18828 16390
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18340 15320 18460 15348
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17972 10130 18000 10610
rect 18156 10606 18184 11562
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9722 17908 9862
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9376 17828 9382
rect 17828 9336 17908 9364
rect 17776 9318 17828 9324
rect 17880 8974 17908 9336
rect 17972 8974 18000 10066
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18064 9654 18092 9862
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18248 9110 18276 9998
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17788 6633 17816 6666
rect 17774 6624 17830 6633
rect 17774 6559 17830 6568
rect 17880 4622 17908 8910
rect 17972 6769 18000 8910
rect 17958 6760 18014 6769
rect 17958 6695 18014 6704
rect 18340 5914 18368 15030
rect 18432 13326 18460 15320
rect 18524 13977 18552 15370
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18602 15056 18658 15065
rect 18602 14991 18658 15000
rect 18616 14958 18644 14991
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18708 14550 18736 15098
rect 18786 14920 18842 14929
rect 18786 14855 18788 14864
rect 18840 14855 18842 14864
rect 18788 14826 18840 14832
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18510 13968 18566 13977
rect 18510 13903 18566 13912
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18892 13190 18920 19382
rect 19062 17232 19118 17241
rect 19062 17167 19064 17176
rect 19116 17167 19118 17176
rect 19064 17128 19116 17134
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18984 16250 19012 17002
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18984 14793 19012 14826
rect 18970 14784 19026 14793
rect 18970 14719 19026 14728
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18984 12850 19012 13262
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18616 12102 18644 12718
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18892 12434 18920 12650
rect 18800 12406 18920 12434
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18432 6798 18460 12038
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18524 10130 18552 10474
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5234 18276 5646
rect 18616 5234 18644 12038
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17972 4690 18000 5102
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 18248 4622 18276 5170
rect 18602 4856 18658 4865
rect 18602 4791 18604 4800
rect 18656 4791 18658 4800
rect 18604 4762 18656 4768
rect 18616 4706 18644 4762
rect 18616 4678 18736 4706
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 17684 3936 17736 3942
rect 17776 3936 17828 3942
rect 17684 3878 17736 3884
rect 17774 3904 17776 3913
rect 17828 3904 17830 3913
rect 17774 3839 17830 3848
rect 17408 3596 17460 3602
rect 17236 3556 17408 3584
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17236 2922 17264 3556
rect 17408 3538 17460 3544
rect 17592 3528 17644 3534
rect 17328 3476 17592 3482
rect 17328 3470 17644 3476
rect 17328 3454 17632 3470
rect 17684 3460 17736 3466
rect 17328 2990 17356 3454
rect 17684 3402 17736 3408
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 3058 17448 3334
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17592 3052 17644 3058
rect 17696 3040 17724 3402
rect 17644 3012 17724 3040
rect 17592 2994 17644 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17880 2446 17908 4558
rect 18064 3738 18092 4558
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18432 2922 18460 3470
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18420 2916 18472 2922
rect 18420 2858 18472 2864
rect 18524 2854 18552 3334
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 16500 800 16528 2382
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17236 800 17264 2246
rect 17880 800 17908 2246
rect 18524 898 18552 2790
rect 18616 2650 18644 3470
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18708 2446 18736 4678
rect 18800 4622 18828 12406
rect 19076 11082 19104 15438
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 19168 11014 19196 35866
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 25780 34944 25832 34950
rect 25780 34886 25832 34892
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 25792 27606 25820 34886
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 25780 27600 25832 27606
rect 25780 27542 25832 27548
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 22296 26042 22324 26930
rect 22388 26586 22416 27338
rect 22940 26994 22968 27406
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 23664 27328 23716 27334
rect 23664 27270 23716 27276
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23492 26586 23520 26930
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21192 25702 21220 25842
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19260 18714 19288 19450
rect 19352 18902 19380 19722
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19444 18834 19472 19994
rect 19996 19718 20024 20198
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19310 20024 19654
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19996 18873 20024 19246
rect 19982 18864 20038 18873
rect 19432 18828 19484 18834
rect 19982 18799 20038 18808
rect 19432 18770 19484 18776
rect 19706 18728 19762 18737
rect 19260 18686 19380 18714
rect 19352 18086 19380 18686
rect 19706 18663 19708 18672
rect 19760 18663 19762 18672
rect 19708 18634 19760 18640
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18080 19392 18086
rect 19338 18048 19340 18057
rect 19392 18048 19394 18057
rect 19338 17983 19394 17992
rect 19444 17338 19472 18294
rect 19800 18284 19852 18290
rect 19720 18244 19800 18272
rect 19616 18216 19668 18222
rect 19614 18184 19616 18193
rect 19668 18184 19670 18193
rect 19614 18119 19670 18128
rect 19720 17610 19748 18244
rect 19800 18226 19852 18232
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19812 17882 19840 18022
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19904 17746 19932 18158
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19708 17604 19760 17610
rect 19708 17546 19760 17552
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19248 17264 19300 17270
rect 19246 17232 19248 17241
rect 19300 17232 19302 17241
rect 19246 17167 19302 17176
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16794 19288 17070
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19720 16726 19748 17002
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19260 11898 19288 15982
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 14890 19380 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19352 13326 19380 13942
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19444 13258 19472 13874
rect 19996 13530 20024 18362
rect 20088 17678 20116 20946
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20272 19922 20300 20402
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20180 18970 20208 19314
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20166 18864 20222 18873
rect 20166 18799 20222 18808
rect 20180 18766 20208 18799
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19352 11694 19380 12582
rect 19812 12442 19840 12786
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19996 12238 20024 13126
rect 20180 12594 20208 18702
rect 20272 17270 20300 19450
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20350 18728 20406 18737
rect 20350 18663 20406 18672
rect 20364 17678 20392 18663
rect 20456 18222 20484 18770
rect 20548 18358 20576 20470
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20640 18698 20668 19246
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20824 18986 20852 19178
rect 20824 18958 20944 18986
rect 20916 18902 20944 18958
rect 20720 18896 20772 18902
rect 20904 18896 20956 18902
rect 20772 18856 20852 18884
rect 20720 18838 20772 18844
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 17746 20484 18158
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20456 17338 20484 17478
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20364 17218 20392 17274
rect 20548 17218 20576 18294
rect 20640 18154 20668 18634
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20626 18048 20682 18057
rect 20626 17983 20682 17992
rect 20640 17678 20668 17983
rect 20732 17882 20760 18702
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20824 17746 20852 18856
rect 20904 18838 20956 18844
rect 20916 18290 20944 18838
rect 21100 18630 21128 19314
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20916 17814 20944 18226
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20272 16658 20300 17206
rect 20364 17190 20576 17218
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20272 12918 20300 13738
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20171 12566 20208 12594
rect 20171 12356 20199 12566
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20171 12328 20208 12356
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19352 10674 19380 11630
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19444 10792 19472 11018
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19444 10764 19564 10792
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18892 7698 18920 9658
rect 18984 7818 19012 10406
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19168 9518 19196 10134
rect 19352 9654 19380 10610
rect 19444 10062 19472 10610
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19536 9908 19564 10764
rect 19996 10674 20024 12174
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19444 9880 19564 9908
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 8498 19104 9318
rect 19260 9110 19288 9522
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18892 7670 19196 7698
rect 19168 7426 19196 7670
rect 19352 7546 19380 9318
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19168 7398 19380 7426
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19260 6866 19288 7278
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19352 6390 19380 7398
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18800 4486 18828 4558
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 3534 18828 4422
rect 19076 4078 19104 5170
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18984 3466 19012 4014
rect 19076 3777 19104 4014
rect 19062 3768 19118 3777
rect 19062 3703 19118 3712
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18984 3058 19012 3402
rect 19352 3194 19380 5646
rect 19444 5370 19472 9880
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19536 8974 19564 9522
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19996 7750 20024 10066
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20088 9586 20116 9998
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20088 8362 20116 8910
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19996 7410 20024 7686
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19996 5234 20024 5646
rect 20088 5642 20116 8298
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19432 3052 19484 3058
rect 19708 3052 19760 3058
rect 19484 3012 19708 3040
rect 19432 2994 19484 3000
rect 19708 2994 19760 3000
rect 19996 2922 20024 4014
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 20088 2446 20116 5578
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 18524 870 18644 898
rect 18616 800 18644 870
rect 19260 800 19288 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 1170 20024 2246
rect 20180 2038 20208 12328
rect 20272 2106 20300 12378
rect 20364 7562 20392 17190
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20456 9450 20484 17002
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20548 14822 20576 15030
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 12434 20576 14758
rect 20640 13274 20668 17614
rect 20916 17202 20944 17750
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 21008 17066 21036 18294
rect 21100 18290 21128 18566
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 21100 16998 21128 17682
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20732 15570 20760 16594
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20824 15570 20852 15914
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20732 13394 20760 13806
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20812 13320 20864 13326
rect 20640 13246 20760 13274
rect 20812 13262 20864 13268
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20640 12850 20668 13126
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20732 12442 20760 13246
rect 20824 12442 20852 13262
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20720 12436 20772 12442
rect 20548 12406 20668 12434
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20548 10062 20576 11698
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20640 9738 20668 12406
rect 20720 12378 20772 12384
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20916 12238 20944 12582
rect 21008 12306 21036 13262
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20640 9710 20760 9738
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20444 9444 20496 9450
rect 20444 9386 20496 9392
rect 20456 9110 20484 9386
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20640 8838 20668 9590
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20732 8650 20760 9710
rect 20640 8622 20760 8650
rect 20364 7534 20484 7562
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20364 5574 20392 6054
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 4758 20392 5510
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20456 2650 20484 7534
rect 20640 6662 20668 8622
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20548 5914 20576 6326
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20548 5166 20576 5850
rect 20640 5846 20668 6598
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20640 5370 20668 5510
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20812 5228 20864 5234
rect 20916 5216 20944 12174
rect 21192 10810 21220 25638
rect 22480 25226 22508 25774
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22572 25430 22600 25638
rect 22664 25498 22692 26318
rect 22928 26308 22980 26314
rect 22928 26250 22980 26256
rect 22940 25838 22968 26250
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 23020 25764 23072 25770
rect 23020 25706 23072 25712
rect 23032 25498 23060 25706
rect 23400 25498 23428 26454
rect 22652 25492 22704 25498
rect 22652 25434 22704 25440
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 23584 25362 23612 26726
rect 23676 26234 23704 27270
rect 24872 27130 24900 27338
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24688 26246 24716 26454
rect 23756 26240 23808 26246
rect 23676 26206 23756 26234
rect 23676 25838 23704 26206
rect 23756 26182 23808 26188
rect 24676 26240 24728 26246
rect 24676 26182 24728 26188
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21652 24682 21680 25094
rect 21640 24676 21692 24682
rect 21640 24618 21692 24624
rect 22480 24614 22508 25162
rect 23020 24676 23072 24682
rect 23020 24618 23072 24624
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 18426 21312 19654
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21376 18193 21404 21014
rect 21454 18728 21510 18737
rect 21454 18663 21510 18672
rect 21468 18290 21496 18663
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21362 18184 21418 18193
rect 21362 18119 21418 18128
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21284 17270 21312 17614
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 21376 13802 21404 18119
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21468 17202 21496 17546
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21652 16250 21680 23598
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21744 18426 21772 18702
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21744 16998 21772 18022
rect 21836 17338 21864 24074
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22112 22438 22140 23666
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22020 18970 22048 19722
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 21916 18760 21968 18766
rect 21968 18720 22048 18748
rect 21916 18702 21968 18708
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21928 17814 21956 18158
rect 21916 17808 21968 17814
rect 21916 17750 21968 17756
rect 22020 17746 22048 18720
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 14890 21496 16050
rect 21560 15502 21588 16118
rect 21744 15638 21772 16526
rect 21836 16522 21864 17138
rect 21916 17060 21968 17066
rect 22020 17048 22048 17682
rect 22112 17218 22140 22374
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 18970 22232 20402
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22388 19514 22416 19654
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22296 18850 22324 19110
rect 22204 18822 22324 18850
rect 22204 18290 22232 18822
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22204 18086 22232 18226
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22112 17190 22232 17218
rect 21968 17020 22048 17048
rect 21916 17002 21968 17008
rect 21928 16590 21956 17002
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21836 16114 21864 16458
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21836 15910 21864 16050
rect 21928 15978 21956 16526
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21560 15026 21588 15438
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21376 13326 21404 13738
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21468 7954 21496 14826
rect 21836 14822 21864 15642
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22020 15026 22048 15506
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14346 21864 14758
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 22020 14006 22048 14962
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21836 11898 21864 13262
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 12850 22140 13126
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 22020 11762 22048 12174
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 9926 22140 10406
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9382 22140 9862
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22020 9110 22048 9318
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21548 8560 21600 8566
rect 21548 8502 21600 8508
rect 21560 8294 21588 8502
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21560 7886 21588 8230
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21836 7818 21864 8774
rect 21928 8566 21956 8910
rect 22020 8566 22048 9046
rect 22112 8974 22140 9318
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 22112 8362 22140 8910
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21836 6322 21864 6734
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 22204 5914 22232 17190
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22296 14890 22324 17138
rect 22388 17066 22416 17478
rect 22480 17066 22508 24550
rect 22848 24274 22876 24550
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22572 23746 22600 24006
rect 22664 23866 22692 24210
rect 23032 24138 23060 24618
rect 23584 24342 23612 25298
rect 23676 24750 23704 25774
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24412 25158 24440 25638
rect 25792 25498 25820 27542
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 26988 26994 27016 27406
rect 27528 27056 27580 27062
rect 27528 26998 27580 27004
rect 26976 26988 27028 26994
rect 26976 26930 27028 26936
rect 27068 26988 27120 26994
rect 27068 26930 27120 26936
rect 27080 26586 27108 26930
rect 27068 26580 27120 26586
rect 27068 26522 27120 26528
rect 27540 26382 27568 26998
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 26252 26042 26280 26318
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 27436 25832 27488 25838
rect 27436 25774 27488 25780
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25792 25294 25820 25434
rect 26252 25362 26280 25774
rect 27068 25764 27120 25770
rect 27068 25706 27120 25712
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 24400 25152 24452 25158
rect 24400 25094 24452 25100
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23860 24614 23888 24754
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22572 23718 22692 23746
rect 22664 23662 22692 23718
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 23050 22692 23598
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22664 22098 22692 22986
rect 22652 22092 22704 22098
rect 22940 22094 22968 23054
rect 22652 22034 22704 22040
rect 22848 22066 22968 22094
rect 23032 22094 23060 24074
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23186 23520 24006
rect 23584 23730 23612 24278
rect 23860 24138 23888 24550
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23860 23730 23888 24074
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 24412 23254 24440 25094
rect 24504 24410 24532 25230
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24504 24070 24532 24346
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24400 23248 24452 23254
rect 24400 23190 24452 23196
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 23204 23044 23256 23050
rect 23204 22986 23256 22992
rect 23032 22066 23152 22094
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22572 17882 22600 21966
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22756 21690 22784 21898
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22664 21418 22692 21626
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22652 20324 22704 20330
rect 22652 20266 22704 20272
rect 22664 19990 22692 20266
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22388 16726 22416 17002
rect 22376 16720 22428 16726
rect 22376 16662 22428 16668
rect 22388 16454 22416 16662
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22388 15978 22416 16390
rect 22664 16182 22692 17138
rect 22652 16176 22704 16182
rect 22466 16144 22522 16153
rect 22652 16118 22704 16124
rect 22466 16079 22468 16088
rect 22520 16079 22522 16088
rect 22468 16050 22520 16056
rect 22376 15972 22428 15978
rect 22376 15914 22428 15920
rect 22388 15094 22416 15914
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15570 22508 15846
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22572 12918 22600 13126
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22296 11762 22324 12174
rect 22480 11762 22508 12582
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22388 10470 22416 10746
rect 22664 10690 22692 15030
rect 22480 10662 22692 10690
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22388 10010 22416 10406
rect 22296 9982 22416 10010
rect 22296 9518 22324 9982
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22388 9722 22416 9862
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22388 9178 22416 9658
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22480 9042 22508 10662
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22572 10266 22600 10542
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22572 9654 22600 10202
rect 22756 9738 22784 19790
rect 22848 16794 22876 22066
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22940 20534 22968 20810
rect 22928 20528 22980 20534
rect 22928 20470 22980 20476
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 22940 19446 22968 19926
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 22926 19272 22982 19281
rect 22926 19207 22928 19216
rect 22980 19207 22982 19216
rect 22928 19178 22980 19184
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23032 17202 23060 17750
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23020 17060 23072 17066
rect 23020 17002 23072 17008
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22848 16153 22876 16186
rect 22834 16144 22890 16153
rect 22834 16079 22890 16088
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22940 15910 22968 15982
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22664 9710 22784 9738
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22572 7750 22600 8366
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22480 5710 22508 6190
rect 22572 6118 22600 7686
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5710 22600 6054
rect 22468 5704 22520 5710
rect 22468 5646 22520 5652
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21744 5302 21772 5510
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 20864 5188 20944 5216
rect 20996 5228 21048 5234
rect 20812 5170 20864 5176
rect 20996 5170 21048 5176
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20640 4758 20668 5170
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3602 20668 4082
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20640 3482 20668 3538
rect 20640 3454 20760 3482
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20640 3058 20668 3334
rect 20732 3194 20760 3454
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20548 2582 20576 2926
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 20732 2446 20760 2858
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20260 2100 20312 2106
rect 20260 2042 20312 2048
rect 20168 2032 20220 2038
rect 20168 1974 20220 1980
rect 20732 1714 20760 2382
rect 20824 2378 20852 5170
rect 21008 3126 21036 5170
rect 21100 4690 21128 5170
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 21560 4010 21588 4558
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 22112 3738 22140 4558
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22388 3534 22416 5102
rect 22664 4826 22692 9710
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22756 9178 22784 9522
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22756 4146 22784 5646
rect 22848 4554 22876 11698
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 8974 22968 9862
rect 23032 9654 23060 17002
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22940 8362 22968 8910
rect 22928 8356 22980 8362
rect 22928 8298 22980 8304
rect 22940 7546 22968 8298
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23124 6390 23152 22066
rect 23112 6384 23164 6390
rect 23112 6326 23164 6332
rect 23216 5914 23244 22986
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23308 16658 23336 22034
rect 24044 22030 24072 22374
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23584 21146 23612 21422
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23400 19174 23428 20334
rect 23492 19666 23520 20538
rect 23584 19922 23612 20742
rect 23676 20602 23704 21082
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23768 20466 23796 21830
rect 24124 21684 24176 21690
rect 24124 21626 24176 21632
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 19922 23796 20198
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23572 19712 23624 19718
rect 23492 19660 23572 19666
rect 23492 19654 23624 19660
rect 23492 19638 23612 19654
rect 23584 19514 23612 19638
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23296 16652 23348 16658
rect 23296 16594 23348 16600
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23308 15910 23336 16390
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15706 23336 15846
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23676 14618 23704 17002
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23768 10062 23796 10202
rect 23756 10056 23808 10062
rect 23756 9998 23808 10004
rect 23768 9722 23796 9998
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23308 6866 23336 9590
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23400 8566 23428 9522
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23492 8378 23520 8910
rect 23400 8350 23520 8378
rect 23400 8294 23428 8350
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23400 6322 23428 8230
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 5914 23704 6258
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23572 5840 23624 5846
rect 23572 5782 23624 5788
rect 23584 5710 23612 5782
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 23124 4758 23152 4966
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 22572 3670 22600 3946
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22756 3194 22784 3470
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 20812 2372 20864 2378
rect 20812 2314 20864 2320
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 19904 1142 20024 1170
rect 20640 1686 20760 1714
rect 19904 800 19932 1142
rect 20640 800 20668 1686
rect 21284 800 21312 2246
rect 22020 1170 22048 2246
rect 21928 1142 22048 1170
rect 21928 800 21956 1142
rect 22664 800 22692 2994
rect 22848 2378 22876 4490
rect 23124 4282 23152 4694
rect 23400 4622 23428 5306
rect 23768 4826 23796 5646
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23124 4146 23152 4218
rect 23400 4214 23428 4558
rect 23676 4486 23704 4558
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23388 4208 23440 4214
rect 23388 4150 23440 4156
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23124 3738 23152 4082
rect 23204 4072 23256 4078
rect 23676 4026 23704 4422
rect 23860 4146 23888 19178
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 5370 23980 19110
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12782 24072 13126
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 24044 12306 24072 12718
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24136 5914 24164 21626
rect 24320 21622 24348 22374
rect 24412 22030 24440 22578
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24412 21622 24440 21966
rect 24308 21616 24360 21622
rect 24308 21558 24360 21564
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24228 18154 24256 19790
rect 24320 19378 24348 21286
rect 24412 20942 24440 21558
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24504 21350 24532 21490
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24412 20534 24440 20878
rect 24688 20806 24716 25162
rect 26252 25158 26280 25298
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 26240 25152 26292 25158
rect 26292 25112 26372 25140
rect 26240 25094 26292 25100
rect 25884 24886 25912 25094
rect 25872 24880 25924 24886
rect 25872 24822 25924 24828
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 24872 23322 24900 24686
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24872 22710 24900 23258
rect 24964 22778 24992 23802
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25056 22982 25084 23666
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24964 22030 24992 22714
rect 24952 22024 25004 22030
rect 24766 21992 24822 22001
rect 24952 21966 25004 21972
rect 24766 21927 24822 21936
rect 24780 21418 24808 21927
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24676 20800 24728 20806
rect 24676 20742 24728 20748
rect 24400 20528 24452 20534
rect 24400 20470 24452 20476
rect 24412 20058 24440 20470
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24688 19446 24716 19994
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24872 18698 24900 19790
rect 25056 18698 25084 22918
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 24216 18148 24268 18154
rect 24216 18090 24268 18096
rect 24872 17678 24900 18634
rect 24952 18216 25004 18222
rect 24952 18158 25004 18164
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24780 16590 24808 16934
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24872 16250 24900 17138
rect 24964 16998 24992 18158
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24964 16114 24992 16458
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 25056 15994 25084 18090
rect 25148 17542 25176 20742
rect 25240 20602 25268 22510
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25148 17134 25176 17478
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 24964 15966 25084 15994
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24688 13394 24716 13466
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 12918 24808 13262
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12442 24348 12786
rect 24308 12436 24360 12442
rect 24308 12378 24360 12384
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24412 11898 24440 12174
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24596 11082 24624 11698
rect 24688 11150 24716 12378
rect 24780 12374 24808 12854
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24596 9926 24624 11018
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24504 6866 24532 9522
rect 24596 9042 24624 9862
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24124 5636 24176 5642
rect 24124 5578 24176 5584
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24136 5234 24164 5578
rect 24308 5296 24360 5302
rect 24308 5238 24360 5244
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23256 4020 23704 4026
rect 23204 4014 23704 4020
rect 23216 3998 23704 4014
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23216 3398 23244 3878
rect 23676 3738 23704 3998
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23952 2774 23980 5102
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24032 4684 24084 4690
rect 24032 4626 24084 4632
rect 24044 4146 24072 4626
rect 24228 4622 24256 5034
rect 24320 4622 24348 5238
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24320 4282 24348 4558
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24136 2922 24164 4082
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 3194 24256 3470
rect 24412 3194 24440 5170
rect 24596 4758 24624 6326
rect 24688 5166 24716 11086
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24676 4616 24728 4622
rect 24780 4570 24808 11562
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24872 8430 24900 8910
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24728 4564 24808 4570
rect 24676 4558 24808 4564
rect 24504 3738 24532 4558
rect 24688 4542 24808 4558
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24124 2916 24176 2922
rect 24124 2858 24176 2864
rect 23952 2746 24164 2774
rect 24136 2582 24164 2746
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23308 800 23336 2246
rect 23676 2106 23704 2382
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 23676 1970 23704 2042
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 24044 800 24072 2246
rect 24688 800 24716 2926
rect 24780 2378 24808 4542
rect 24872 4146 24900 5646
rect 24964 4826 24992 15966
rect 25148 15094 25176 17070
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25240 15910 25268 16934
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25240 15706 25268 15846
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25056 11762 25084 12582
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25056 11626 25084 11698
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 25044 11620 25096 11626
rect 25044 11562 25096 11568
rect 25148 11150 25176 11630
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25240 9330 25268 14758
rect 25332 12238 25360 22374
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25608 17202 25636 17478
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25424 16114 25452 16390
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25424 14822 25452 16050
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25332 11762 25360 12038
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25320 11620 25372 11626
rect 25320 11562 25372 11568
rect 25332 11218 25360 11562
rect 25424 11354 25452 12242
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25516 10810 25544 15030
rect 25608 14482 25636 15302
rect 25792 14940 25820 18634
rect 25884 16114 25912 24822
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 26252 23322 26280 24754
rect 26344 24682 26372 25112
rect 27080 24954 27108 25706
rect 27344 25220 27396 25226
rect 27344 25162 27396 25168
rect 27068 24948 27120 24954
rect 27068 24890 27120 24896
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27068 24336 27120 24342
rect 27068 24278 27120 24284
rect 26884 23520 26936 23526
rect 26884 23462 26936 23468
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26896 23254 26924 23462
rect 26884 23248 26936 23254
rect 26884 23190 26936 23196
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26148 22094 26200 22098
rect 26252 22094 26280 23122
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 26804 22574 26832 22918
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 27080 22506 27108 24278
rect 27172 24070 27200 24618
rect 27356 24614 27384 25162
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27448 24274 27476 25774
rect 27540 25226 27568 26318
rect 27632 26314 27660 28358
rect 28368 27130 28396 32846
rect 28448 30592 28500 30598
rect 28448 30534 28500 30540
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 27620 26308 27672 26314
rect 27620 26250 27672 26256
rect 27896 26308 27948 26314
rect 27896 26250 27948 26256
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27436 24268 27488 24274
rect 27436 24210 27488 24216
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 27172 22658 27200 24006
rect 27344 23588 27396 23594
rect 27344 23530 27396 23536
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 27264 22778 27292 22986
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27172 22630 27292 22658
rect 27068 22500 27120 22506
rect 27068 22442 27120 22448
rect 26332 22160 26384 22166
rect 26332 22102 26384 22108
rect 26148 22092 26280 22094
rect 26200 22066 26280 22092
rect 26148 22034 26200 22040
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25976 21554 26004 21830
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25976 17814 26004 18226
rect 25964 17808 26016 17814
rect 25964 17750 26016 17756
rect 25976 17202 26004 17750
rect 26148 17672 26200 17678
rect 26252 17660 26280 21966
rect 26344 21418 26372 22102
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26528 21690 26556 21898
rect 26516 21684 26568 21690
rect 26516 21626 26568 21632
rect 27160 21480 27212 21486
rect 27160 21422 27212 21428
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 27172 20874 27200 21422
rect 27160 20868 27212 20874
rect 27160 20810 27212 20816
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 26200 17632 26280 17660
rect 26148 17614 26200 17620
rect 25964 17196 26016 17202
rect 25964 17138 26016 17144
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 25884 15094 25912 16050
rect 25976 15434 26004 17138
rect 26252 16794 26280 17632
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26252 16114 26280 16390
rect 26436 16250 26464 17546
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26896 16046 26924 16526
rect 26988 16114 27016 17274
rect 27080 16590 27108 17478
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25976 15314 26004 15370
rect 26896 15366 26924 15982
rect 27080 15638 27108 16526
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 27080 15434 27108 15574
rect 27068 15428 27120 15434
rect 27068 15370 27120 15376
rect 26884 15360 26936 15366
rect 25976 15286 26096 15314
rect 26884 15302 26936 15308
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25792 14912 25912 14940
rect 25780 14816 25832 14822
rect 25780 14758 25832 14764
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25608 11286 25636 13262
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 12238 25728 12582
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25596 11280 25648 11286
rect 25596 11222 25648 11228
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25424 9586 25452 10610
rect 25516 10130 25544 10746
rect 25792 10674 25820 14758
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25516 9382 25544 9930
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25504 9376 25556 9382
rect 25240 9302 25360 9330
rect 25504 9318 25556 9324
rect 25136 9104 25188 9110
rect 25136 9046 25188 9052
rect 25148 8498 25176 9046
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25240 8498 25268 8842
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25148 5846 25176 8434
rect 25332 6866 25360 9302
rect 25608 9178 25636 9522
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25608 8498 25636 8910
rect 25792 8634 25820 9998
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25884 5914 25912 14912
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25976 13938 26004 14418
rect 26068 13938 26096 15286
rect 26896 15094 26924 15302
rect 26884 15088 26936 15094
rect 26884 15030 26936 15036
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 26068 13258 26096 13874
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26160 11898 26188 12786
rect 26528 12170 26556 13262
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25976 11150 26004 11698
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25976 8362 26004 8910
rect 25964 8356 26016 8362
rect 25964 8298 26016 8304
rect 25976 7954 26004 8298
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 26068 7886 26096 9318
rect 26160 8906 26188 9862
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26056 6860 26108 6866
rect 26056 6802 26108 6808
rect 26068 6118 26096 6802
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 25976 5846 26004 6054
rect 25136 5840 25188 5846
rect 25136 5782 25188 5788
rect 25964 5840 26016 5846
rect 25964 5782 26016 5788
rect 26146 5808 26202 5817
rect 26146 5743 26202 5752
rect 26424 5772 26476 5778
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 25700 4758 25728 4966
rect 25792 4758 25820 4966
rect 25688 4752 25740 4758
rect 25688 4694 25740 4700
rect 25780 4752 25832 4758
rect 25780 4694 25832 4700
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 25056 3534 25084 4082
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 25136 4004 25188 4010
rect 25136 3946 25188 3952
rect 25228 4004 25280 4010
rect 25228 3946 25280 3952
rect 25148 3602 25176 3946
rect 25240 3670 25268 3946
rect 25424 3738 25452 4014
rect 25412 3732 25464 3738
rect 25412 3674 25464 3680
rect 25228 3664 25280 3670
rect 25228 3606 25280 3612
rect 25780 3664 25832 3670
rect 25780 3606 25832 3612
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25056 3210 25084 3470
rect 24964 3194 25084 3210
rect 25148 3194 25176 3538
rect 25240 3466 25268 3606
rect 25228 3460 25280 3466
rect 25228 3402 25280 3408
rect 24952 3188 25084 3194
rect 25004 3182 25084 3188
rect 25136 3188 25188 3194
rect 24952 3130 25004 3136
rect 25136 3130 25188 3136
rect 25240 2922 25268 3402
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 25792 2650 25820 3606
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25792 2446 25820 2586
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 25332 800 25360 2246
rect 25884 2106 25912 4558
rect 26068 2650 26096 5646
rect 26160 5370 26188 5743
rect 26424 5714 26476 5720
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 26436 4622 26464 5714
rect 26424 4616 26476 4622
rect 26424 4558 26476 4564
rect 26436 4282 26464 4558
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 2938 26280 3334
rect 26160 2910 26280 2938
rect 26620 2922 26648 12038
rect 26896 11898 26924 15030
rect 27172 12986 27200 18158
rect 27264 18086 27292 22630
rect 27356 22574 27384 23530
rect 27448 23186 27476 24210
rect 27540 23202 27568 25162
rect 27632 23594 27660 26250
rect 27908 26042 27936 26250
rect 27896 26036 27948 26042
rect 27896 25978 27948 25984
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 27712 24948 27764 24954
rect 27712 24890 27764 24896
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 27540 23186 27660 23202
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27540 23180 27672 23186
rect 27540 23174 27620 23180
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27448 22098 27476 23122
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27356 21078 27384 21490
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27448 20602 27476 22034
rect 27540 22030 27568 23174
rect 27620 23122 27672 23128
rect 27620 22976 27672 22982
rect 27620 22918 27672 22924
rect 27632 22778 27660 22918
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27540 21622 27568 21966
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27632 21486 27660 22510
rect 27724 21978 27752 24890
rect 28092 24410 28120 25842
rect 28264 24948 28316 24954
rect 28264 24890 28316 24896
rect 28276 24750 28304 24890
rect 28368 24818 28396 27066
rect 28460 25498 28488 30534
rect 32140 28218 32168 36042
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 36004 31822 36032 37062
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 32128 28212 32180 28218
rect 32128 28154 32180 28160
rect 32864 28212 32916 28218
rect 32864 28154 32916 28160
rect 32036 27532 32088 27538
rect 32036 27474 32088 27480
rect 30564 27396 30616 27402
rect 30564 27338 30616 27344
rect 30576 27130 30604 27338
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 30852 26586 30880 26930
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 30288 26512 30340 26518
rect 30288 26454 30340 26460
rect 30932 26512 30984 26518
rect 30932 26454 30984 26460
rect 30300 25498 30328 26454
rect 30944 26042 30972 26454
rect 31312 26314 31340 27066
rect 31392 26852 31444 26858
rect 31392 26794 31444 26800
rect 31300 26308 31352 26314
rect 31300 26250 31352 26256
rect 30932 26036 30984 26042
rect 30932 25978 30984 25984
rect 30380 25900 30432 25906
rect 30380 25842 30432 25848
rect 28448 25492 28500 25498
rect 28448 25434 28500 25440
rect 30288 25492 30340 25498
rect 30288 25434 30340 25440
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 28264 24744 28316 24750
rect 28264 24686 28316 24692
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 28460 24342 28488 25434
rect 30392 24750 30420 25842
rect 31312 25158 31340 26250
rect 31404 26042 31432 26794
rect 31760 26784 31812 26790
rect 31760 26726 31812 26732
rect 31772 26382 31800 26726
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 32048 26314 32076 27474
rect 32220 26988 32272 26994
rect 32220 26930 32272 26936
rect 32232 26586 32260 26930
rect 32220 26580 32272 26586
rect 32220 26522 32272 26528
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32036 26308 32088 26314
rect 32036 26250 32088 26256
rect 32600 26246 32628 26386
rect 32588 26240 32640 26246
rect 32588 26182 32640 26188
rect 31392 26036 31444 26042
rect 31392 25978 31444 25984
rect 32600 25838 32628 26182
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32588 25832 32640 25838
rect 32588 25774 32640 25780
rect 32600 25702 32628 25774
rect 32588 25696 32640 25702
rect 32588 25638 32640 25644
rect 32600 25362 32628 25638
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 30472 25152 30524 25158
rect 30472 25094 30524 25100
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 30484 24818 30512 25094
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 27896 24336 27948 24342
rect 27896 24278 27948 24284
rect 28448 24336 28500 24342
rect 28448 24278 28500 24284
rect 27908 23866 27936 24278
rect 28908 24132 28960 24138
rect 28908 24074 28960 24080
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 28264 22704 28316 22710
rect 28264 22646 28316 22652
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 22166 27844 22374
rect 27804 22160 27856 22166
rect 27804 22102 27856 22108
rect 28276 22098 28304 22646
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 28264 22092 28316 22098
rect 28264 22034 28316 22040
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 27802 21992 27858 22001
rect 27724 21950 27802 21978
rect 27858 21950 28028 21978
rect 28092 21962 28120 22034
rect 27802 21927 27858 21936
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27540 19854 27568 20266
rect 27632 19922 27660 21422
rect 27816 21418 27844 21830
rect 27804 21412 27856 21418
rect 27804 21354 27856 21360
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 27724 20262 27752 20402
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27540 18358 27568 19790
rect 27632 19446 27660 19858
rect 27620 19440 27672 19446
rect 27620 19382 27672 19388
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27632 18630 27660 19110
rect 27724 18766 27752 20198
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27632 18290 27660 18566
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 26976 9988 27028 9994
rect 26976 9930 27028 9936
rect 26988 9722 27016 9930
rect 26976 9716 27028 9722
rect 26976 9658 27028 9664
rect 27264 9654 27292 18022
rect 27632 17882 27660 18226
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27356 14822 27384 17070
rect 27632 16561 27660 17818
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 27618 16552 27674 16561
rect 27436 16516 27488 16522
rect 27618 16487 27674 16496
rect 27436 16458 27488 16464
rect 27448 16114 27476 16458
rect 27724 16250 27752 17138
rect 28000 17134 28028 21950
rect 28080 21956 28132 21962
rect 28080 21898 28132 21904
rect 28460 21706 28488 22034
rect 28644 22030 28672 24006
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28736 22574 28764 23462
rect 28828 22930 28856 23598
rect 28920 23118 28948 24074
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28828 22902 28948 22930
rect 28920 22642 28948 22902
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28276 21690 28488 21706
rect 28264 21684 28488 21690
rect 28316 21678 28488 21684
rect 28264 21626 28316 21632
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27816 16590 27844 16934
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27632 10266 27660 10678
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27264 8634 27292 8774
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 27724 8498 27752 9930
rect 28092 9674 28120 18702
rect 28276 18222 28304 21626
rect 28736 21350 28764 22510
rect 28920 22234 28948 22578
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28920 22098 28948 22170
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 29012 21894 29040 23802
rect 29460 23316 29512 23322
rect 29460 23258 29512 23264
rect 29472 22778 29500 23258
rect 29460 22772 29512 22778
rect 29460 22714 29512 22720
rect 31024 22432 31076 22438
rect 31024 22374 31076 22380
rect 29828 21956 29880 21962
rect 29828 21898 29880 21904
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29840 21690 29868 21898
rect 30932 21888 30984 21894
rect 30932 21830 30984 21836
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29460 21548 29512 21554
rect 29460 21490 29512 21496
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28816 19916 28868 19922
rect 28954 19916 29006 19922
rect 28868 19876 28954 19904
rect 28816 19858 28868 19864
rect 28954 19858 29006 19864
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28632 19304 28684 19310
rect 28632 19246 28684 19252
rect 28644 18766 28672 19246
rect 28920 19242 28948 19654
rect 29104 19514 29132 19790
rect 29092 19508 29144 19514
rect 29092 19450 29144 19456
rect 28908 19236 28960 19242
rect 28908 19178 28960 19184
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28264 18216 28316 18222
rect 28264 18158 28316 18164
rect 29276 18148 29328 18154
rect 29276 18090 29328 18096
rect 28540 17060 28592 17066
rect 28540 17002 28592 17008
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 28184 16250 28212 16390
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28552 13530 28580 17002
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28552 12850 28580 13466
rect 28540 12844 28592 12850
rect 28540 12786 28592 12792
rect 28172 12776 28224 12782
rect 28172 12718 28224 12724
rect 28184 10470 28212 12718
rect 28540 11892 28592 11898
rect 28540 11834 28592 11840
rect 28552 11694 28580 11834
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 28920 11626 28948 14962
rect 29012 13841 29040 15302
rect 29184 14816 29236 14822
rect 29184 14758 29236 14764
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 29104 14074 29132 14214
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29196 13938 29224 14758
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 28998 13832 29054 13841
rect 28998 13767 29054 13776
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 29104 11898 29132 12786
rect 29288 12434 29316 18090
rect 29472 16182 29500 21490
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29748 20058 29776 20402
rect 30944 20398 30972 21830
rect 31036 21146 31064 22374
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30116 18222 30144 18702
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30116 17610 30144 18158
rect 30288 18148 30340 18154
rect 30288 18090 30340 18096
rect 29644 17604 29696 17610
rect 29644 17546 29696 17552
rect 30104 17604 30156 17610
rect 30104 17546 30156 17552
rect 29656 17202 29684 17546
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29748 16590 29776 16934
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29460 16176 29512 16182
rect 29460 16118 29512 16124
rect 29368 14340 29420 14346
rect 29368 14282 29420 14288
rect 29380 14074 29408 14282
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29472 12918 29500 16118
rect 29552 13320 29604 13326
rect 29552 13262 29604 13268
rect 29460 12912 29512 12918
rect 29460 12854 29512 12860
rect 29288 12406 29408 12434
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 29288 11354 29316 11698
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 28172 10464 28224 10470
rect 28172 10406 28224 10412
rect 28000 9646 28120 9674
rect 28000 8838 28028 9646
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28644 8906 28672 9522
rect 28632 8900 28684 8906
rect 28632 8842 28684 8848
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27448 7750 27476 8366
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27448 6338 27476 7686
rect 27724 7426 27752 8434
rect 28000 8430 28028 8774
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 28000 8022 28028 8366
rect 28644 8022 28672 8842
rect 27988 8016 28040 8022
rect 27988 7958 28040 7964
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 27724 7410 27844 7426
rect 27724 7404 27856 7410
rect 27724 7398 27804 7404
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27540 6934 27568 7142
rect 27528 6928 27580 6934
rect 27528 6870 27580 6876
rect 27448 6310 27568 6338
rect 27540 5642 27568 6310
rect 27724 5778 27752 7398
rect 27804 7346 27856 7352
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 29000 6180 29052 6186
rect 29000 6122 29052 6128
rect 29012 5914 29040 6122
rect 29000 5908 29052 5914
rect 29000 5850 29052 5856
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27434 5264 27490 5273
rect 27434 5199 27490 5208
rect 26790 4992 26846 5001
rect 26790 4927 26846 4936
rect 26804 4826 26832 4927
rect 27448 4826 27476 5199
rect 26792 4820 26844 4826
rect 26792 4762 26844 4768
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 26988 3194 27016 3470
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26608 2916 26660 2922
rect 26056 2644 26108 2650
rect 26056 2586 26108 2592
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 25872 2100 25924 2106
rect 25872 2042 25924 2048
rect 26068 800 26096 2246
rect 26160 1970 26188 2910
rect 26608 2858 26660 2864
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26252 2514 26280 2790
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26148 1964 26200 1970
rect 26148 1906 26200 1912
rect 26712 800 26740 2994
rect 26976 2916 27028 2922
rect 26976 2858 27028 2864
rect 26988 2378 27016 2858
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27356 800 27384 2246
rect 27540 1970 27568 5578
rect 27724 5302 27752 5714
rect 29012 5370 29040 5850
rect 29000 5364 29052 5370
rect 29000 5306 29052 5312
rect 27712 5296 27764 5302
rect 27712 5238 27764 5244
rect 27724 4622 27752 5238
rect 29104 5166 29132 6802
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 27804 5092 27856 5098
rect 27804 5034 27856 5040
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27816 2854 27844 5034
rect 28632 5024 28684 5030
rect 28632 4966 28684 4972
rect 28644 4622 28672 4966
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28552 4486 28580 4558
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 27896 4276 27948 4282
rect 27896 4218 27948 4224
rect 27908 3942 27936 4218
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27908 3466 27936 3878
rect 27896 3460 27948 3466
rect 27896 3402 27948 3408
rect 28552 3194 28580 4422
rect 28644 4282 28672 4558
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27724 2038 27752 2382
rect 28080 2304 28132 2310
rect 28080 2246 28132 2252
rect 27712 2032 27764 2038
rect 27712 1974 27764 1980
rect 27528 1964 27580 1970
rect 27528 1906 27580 1912
rect 28092 800 28120 2246
rect 28736 800 28764 3470
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28828 3126 28856 3334
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 28920 2378 28948 4082
rect 29012 4010 29040 4422
rect 29104 4214 29132 5102
rect 29184 5092 29236 5098
rect 29184 5034 29236 5040
rect 29196 4690 29224 5034
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29092 4208 29144 4214
rect 29092 4150 29144 4156
rect 29000 4004 29052 4010
rect 29000 3946 29052 3952
rect 29380 3738 29408 12406
rect 29564 12238 29592 13262
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29656 12850 29684 13194
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29656 12238 29684 12582
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29564 10538 29592 12174
rect 29748 10606 29776 16526
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30024 15502 30052 16390
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30116 14958 30144 17546
rect 30300 17338 30328 18090
rect 30656 17876 30708 17882
rect 30656 17818 30708 17824
rect 30472 17808 30524 17814
rect 30472 17750 30524 17756
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30392 17134 30420 17614
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30392 16658 30420 17070
rect 30484 16794 30512 17750
rect 30668 17270 30696 17818
rect 30944 17678 30972 20334
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 31128 17610 31156 18022
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 30760 16998 30788 17206
rect 30748 16992 30800 16998
rect 30748 16934 30800 16940
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 30472 16788 30524 16794
rect 30472 16730 30524 16736
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30104 14952 30156 14958
rect 30104 14894 30156 14900
rect 29920 14884 29972 14890
rect 29920 14826 29972 14832
rect 29932 14074 29960 14826
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 30012 13456 30064 13462
rect 30012 13398 30064 13404
rect 30024 12986 30052 13398
rect 30116 13394 30144 14894
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30196 14272 30248 14278
rect 30196 14214 30248 14220
rect 30208 14074 30236 14214
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30208 13938 30236 14010
rect 30196 13932 30248 13938
rect 30196 13874 30248 13880
rect 30104 13388 30156 13394
rect 30104 13330 30156 13336
rect 30300 13326 30328 14350
rect 30392 13802 30420 16594
rect 31220 16590 31248 16934
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30012 12980 30064 12986
rect 30012 12922 30064 12928
rect 30392 12782 30420 13738
rect 30576 13530 30604 13874
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30944 13326 30972 13670
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31220 12986 31248 13262
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 30392 11218 30420 12718
rect 30484 11558 30512 12922
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 30944 11762 30972 12038
rect 30932 11756 30984 11762
rect 30932 11698 30984 11704
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30564 11076 30616 11082
rect 30564 11018 30616 11024
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29552 10532 29604 10538
rect 29552 10474 29604 10480
rect 29564 10062 29592 10474
rect 30300 10198 30328 10950
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30576 10130 30604 11018
rect 31036 10742 31064 11698
rect 31024 10736 31076 10742
rect 31024 10678 31076 10684
rect 30564 10124 30616 10130
rect 30564 10066 30616 10072
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29564 8362 29592 9998
rect 30012 9988 30064 9994
rect 30012 9930 30064 9936
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29748 8634 29776 8774
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 30024 8430 30052 9930
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30668 9586 30696 9862
rect 30852 9722 30880 9930
rect 30840 9716 30892 9722
rect 30840 9658 30892 9664
rect 31312 9654 31340 25094
rect 32600 24614 32628 25298
rect 32784 25158 32812 25842
rect 32876 25838 32904 28154
rect 33232 28076 33284 28082
rect 33232 28018 33284 28024
rect 33244 27606 33272 28018
rect 33508 28008 33560 28014
rect 33508 27950 33560 27956
rect 33232 27600 33284 27606
rect 33232 27542 33284 27548
rect 33520 27470 33548 27950
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 36096 27606 36124 37198
rect 37280 37120 37332 37126
rect 37280 37062 37332 37068
rect 38016 37120 38068 37126
rect 38016 37062 38068 37068
rect 36912 36032 36964 36038
rect 36912 35974 36964 35980
rect 36084 27600 36136 27606
rect 36084 27542 36136 27548
rect 33508 27464 33560 27470
rect 33508 27406 33560 27412
rect 35348 27464 35400 27470
rect 35348 27406 35400 27412
rect 32956 27328 33008 27334
rect 32956 27270 33008 27276
rect 32968 25974 32996 27270
rect 33520 27062 33548 27406
rect 34152 27396 34204 27402
rect 34152 27338 34204 27344
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33692 27328 33744 27334
rect 33692 27270 33744 27276
rect 33612 27130 33640 27270
rect 33600 27124 33652 27130
rect 33600 27066 33652 27072
rect 33508 27056 33560 27062
rect 33508 26998 33560 27004
rect 33508 26920 33560 26926
rect 33508 26862 33560 26868
rect 33520 26790 33548 26862
rect 33508 26784 33560 26790
rect 33508 26726 33560 26732
rect 33140 26308 33192 26314
rect 33140 26250 33192 26256
rect 32956 25968 33008 25974
rect 32956 25910 33008 25916
rect 32864 25832 32916 25838
rect 32864 25774 32916 25780
rect 32876 25294 32904 25774
rect 33152 25770 33180 26250
rect 33520 26042 33548 26726
rect 33612 26382 33640 27066
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33508 26036 33560 26042
rect 33508 25978 33560 25984
rect 33140 25764 33192 25770
rect 33140 25706 33192 25712
rect 32864 25288 32916 25294
rect 32864 25230 32916 25236
rect 32772 25152 32824 25158
rect 32772 25094 32824 25100
rect 32784 24886 32812 25094
rect 32772 24880 32824 24886
rect 32772 24822 32824 24828
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 31392 24064 31444 24070
rect 31392 24006 31444 24012
rect 31404 23866 31432 24006
rect 31392 23860 31444 23866
rect 31392 23802 31444 23808
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 31404 22030 31432 23054
rect 31484 23044 31536 23050
rect 31484 22986 31536 22992
rect 31496 22778 31524 22986
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 32496 22568 32548 22574
rect 32496 22510 32548 22516
rect 32220 22500 32272 22506
rect 32220 22442 32272 22448
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 32232 21690 32260 22442
rect 32508 22094 32536 22510
rect 32324 22066 32536 22094
rect 32220 21684 32272 21690
rect 32220 21626 32272 21632
rect 32324 21486 32352 22066
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32312 21480 32364 21486
rect 32312 21422 32364 21428
rect 31944 21412 31996 21418
rect 31944 21354 31996 21360
rect 31956 21146 31984 21354
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31404 19922 31432 20742
rect 32324 20466 32352 21422
rect 32416 20942 32444 21830
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32416 18766 32444 19654
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 32600 18630 32628 24550
rect 33704 23322 33732 27270
rect 34164 27130 34192 27338
rect 34152 27124 34204 27130
rect 34152 27066 34204 27072
rect 34152 26988 34204 26994
rect 34152 26930 34204 26936
rect 34164 26586 34192 26930
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35360 25362 35388 27406
rect 35992 27056 36044 27062
rect 35992 26998 36044 27004
rect 36004 26586 36032 26998
rect 35992 26580 36044 26586
rect 35992 26522 36044 26528
rect 36096 26450 36124 27542
rect 36636 27124 36688 27130
rect 36636 27066 36688 27072
rect 36268 26580 36320 26586
rect 36268 26522 36320 26528
rect 36084 26444 36136 26450
rect 36084 26386 36136 26392
rect 36096 26234 36124 26386
rect 36280 26382 36308 26522
rect 36544 26444 36596 26450
rect 36544 26386 36596 26392
rect 36268 26376 36320 26382
rect 36268 26318 36320 26324
rect 36096 26206 36216 26234
rect 36084 25696 36136 25702
rect 36084 25638 36136 25644
rect 35348 25356 35400 25362
rect 35348 25298 35400 25304
rect 35360 24818 35388 25298
rect 35532 25220 35584 25226
rect 35532 25162 35584 25168
rect 35900 25220 35952 25226
rect 35900 25162 35952 25168
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34152 23724 34204 23730
rect 34152 23666 34204 23672
rect 33692 23316 33744 23322
rect 33692 23258 33744 23264
rect 32772 22976 32824 22982
rect 32772 22918 32824 22924
rect 32784 21690 32812 22918
rect 33968 22704 34020 22710
rect 33968 22646 34020 22652
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 32772 21684 32824 21690
rect 32772 21626 32824 21632
rect 32956 21480 33008 21486
rect 32956 21422 33008 21428
rect 32968 21010 32996 21422
rect 33520 21350 33548 21966
rect 33980 21554 34008 22646
rect 34060 22500 34112 22506
rect 34060 22442 34112 22448
rect 34072 21690 34100 22442
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 33968 21548 34020 21554
rect 33968 21490 34020 21496
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 34164 21146 34192 23666
rect 34532 22778 34560 24142
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35072 23248 35124 23254
rect 35072 23190 35124 23196
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 34532 22234 34560 22578
rect 34624 22574 34652 22986
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 34520 22228 34572 22234
rect 34520 22170 34572 22176
rect 34624 22030 34652 22510
rect 34704 22160 34756 22166
rect 34704 22102 34756 22108
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 32956 21004 33008 21010
rect 32956 20946 33008 20952
rect 32968 20058 32996 20946
rect 34164 20942 34192 21082
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 34716 20806 34744 22102
rect 34808 21486 34836 22510
rect 35084 22506 35112 23190
rect 35072 22500 35124 22506
rect 35072 22442 35124 22448
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35360 22098 35388 24754
rect 35544 24410 35572 25162
rect 35532 24404 35584 24410
rect 35532 24346 35584 24352
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 35820 22234 35848 22578
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35348 22092 35400 22098
rect 35348 22034 35400 22040
rect 35912 21622 35940 25162
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 36004 24410 36032 24754
rect 35992 24404 36044 24410
rect 35992 24346 36044 24352
rect 36096 23798 36124 25638
rect 36188 25498 36216 26206
rect 36280 25906 36308 26318
rect 36556 25906 36584 26386
rect 36268 25900 36320 25906
rect 36268 25842 36320 25848
rect 36544 25900 36596 25906
rect 36544 25842 36596 25848
rect 36268 25764 36320 25770
rect 36268 25706 36320 25712
rect 36176 25492 36228 25498
rect 36176 25434 36228 25440
rect 36280 24410 36308 25706
rect 36556 25226 36584 25842
rect 36544 25220 36596 25226
rect 36544 25162 36596 25168
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 36176 24200 36228 24206
rect 36176 24142 36228 24148
rect 36084 23792 36136 23798
rect 36084 23734 36136 23740
rect 36188 23322 36216 24142
rect 36176 23316 36228 23322
rect 36176 23258 36228 23264
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 35992 22228 36044 22234
rect 35992 22170 36044 22176
rect 35900 21616 35952 21622
rect 35900 21558 35952 21564
rect 34796 21480 34848 21486
rect 34796 21422 34848 21428
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 21010 35388 21422
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 36004 20806 36032 22170
rect 36096 22030 36124 22374
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 36084 21344 36136 21350
rect 36084 21286 36136 21292
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 33048 20392 33100 20398
rect 33048 20334 33100 20340
rect 32956 20052 33008 20058
rect 32956 19994 33008 20000
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 31864 17610 31892 18566
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 31852 17604 31904 17610
rect 31852 17546 31904 17552
rect 31576 17536 31628 17542
rect 31576 17478 31628 17484
rect 31588 17202 31616 17478
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31864 17105 31892 17546
rect 31850 17096 31906 17105
rect 31850 17031 31906 17040
rect 32324 16726 32352 18158
rect 32312 16720 32364 16726
rect 32312 16662 32364 16668
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 31760 14952 31812 14958
rect 31760 14894 31812 14900
rect 31772 14618 31800 14894
rect 31760 14612 31812 14618
rect 31760 14554 31812 14560
rect 31772 14074 31800 14554
rect 31760 14068 31812 14074
rect 31760 14010 31812 14016
rect 32036 13524 32088 13530
rect 32036 13466 32088 13472
rect 32048 12986 32076 13466
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31404 11762 31432 12582
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31760 11348 31812 11354
rect 31760 11290 31812 11296
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30300 8430 30328 9318
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30012 8424 30064 8430
rect 30012 8366 30064 8372
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29472 4826 29500 5102
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29564 4622 29592 8298
rect 30024 7954 30052 8366
rect 30104 8288 30156 8294
rect 30104 8230 30156 8236
rect 30116 8022 30144 8230
rect 30104 8016 30156 8022
rect 30104 7958 30156 7964
rect 30012 7948 30064 7954
rect 30012 7890 30064 7896
rect 30024 6866 30052 7890
rect 30300 7478 30328 8366
rect 30668 8022 30696 8910
rect 31024 8832 31076 8838
rect 31024 8774 31076 8780
rect 30656 8016 30708 8022
rect 30656 7958 30708 7964
rect 31036 7886 31064 8774
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 30288 7472 30340 7478
rect 30208 7420 30288 7426
rect 30208 7414 30340 7420
rect 30208 7398 30328 7414
rect 30472 7404 30524 7410
rect 30104 7200 30156 7206
rect 30104 7142 30156 7148
rect 30116 6934 30144 7142
rect 30104 6928 30156 6934
rect 30104 6870 30156 6876
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 30208 5166 30236 7398
rect 30472 7346 30524 7352
rect 30288 7336 30340 7342
rect 30288 7278 30340 7284
rect 30300 6730 30328 7278
rect 30484 6866 30512 7346
rect 30852 7002 30880 7822
rect 31116 7200 31168 7206
rect 31116 7142 31168 7148
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 30852 6866 30880 6938
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30840 6860 30892 6866
rect 30840 6802 30892 6808
rect 31128 6798 31156 7142
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 30288 6724 30340 6730
rect 30288 6666 30340 6672
rect 30196 5160 30248 5166
rect 30116 5108 30196 5114
rect 30116 5102 30248 5108
rect 30116 5086 30236 5102
rect 29826 4720 29882 4729
rect 29826 4655 29882 4664
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 29368 3732 29420 3738
rect 29368 3674 29420 3680
rect 29380 2446 29408 3674
rect 29472 3126 29500 3878
rect 29460 3120 29512 3126
rect 29460 3062 29512 3068
rect 29564 3058 29592 4558
rect 29840 4214 29868 4655
rect 29828 4208 29880 4214
rect 29828 4150 29880 4156
rect 29840 3738 29868 4150
rect 30116 4078 30144 5086
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 30208 4622 30236 4966
rect 31312 4690 31340 9590
rect 31772 9586 31800 11290
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31772 9042 31800 9522
rect 32128 9172 32180 9178
rect 32128 9114 32180 9120
rect 31760 9036 31812 9042
rect 31760 8978 31812 8984
rect 31772 8838 31800 8978
rect 32140 8974 32168 9114
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31760 8832 31812 8838
rect 31760 8774 31812 8780
rect 32232 5370 32260 16458
rect 32324 16454 32352 16662
rect 32312 16448 32364 16454
rect 32312 16390 32364 16396
rect 32496 11620 32548 11626
rect 32496 11562 32548 11568
rect 32508 11286 32536 11562
rect 32496 11280 32548 11286
rect 32496 11222 32548 11228
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 32324 8566 32352 10610
rect 32600 9654 32628 18566
rect 33060 16114 33088 20334
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 36096 19854 36124 21286
rect 36176 20800 36228 20806
rect 36176 20742 36228 20748
rect 36188 20641 36216 20742
rect 36174 20632 36230 20641
rect 36174 20567 36230 20576
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 34796 19168 34848 19174
rect 34796 19110 34848 19116
rect 34808 18630 34836 19110
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34796 18624 34848 18630
rect 34796 18566 34848 18572
rect 35716 18624 35768 18630
rect 35716 18566 35768 18572
rect 35728 18290 35756 18566
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 35716 18284 35768 18290
rect 35716 18226 35768 18232
rect 34428 17604 34480 17610
rect 34428 17546 34480 17552
rect 33968 17264 34020 17270
rect 33968 17206 34020 17212
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 33232 17128 33284 17134
rect 33232 17070 33284 17076
rect 33152 16726 33180 17070
rect 33140 16720 33192 16726
rect 33140 16662 33192 16668
rect 33048 16108 33100 16114
rect 33048 16050 33100 16056
rect 33060 11354 33088 16050
rect 33244 16046 33272 17070
rect 33980 16726 34008 17206
rect 34440 17066 34468 17546
rect 34532 17338 34560 18226
rect 34796 18080 34848 18086
rect 34796 18022 34848 18028
rect 34808 17610 34836 18022
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 35346 17640 35402 17649
rect 34796 17604 34848 17610
rect 35346 17575 35402 17584
rect 34796 17546 34848 17552
rect 35360 17338 35388 17575
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 35348 17332 35400 17338
rect 35348 17274 35400 17280
rect 35360 17134 35388 17274
rect 35348 17128 35400 17134
rect 35348 17070 35400 17076
rect 34428 17060 34480 17066
rect 34428 17002 34480 17008
rect 34060 16788 34112 16794
rect 34060 16730 34112 16736
rect 33968 16720 34020 16726
rect 33968 16662 34020 16668
rect 33232 16040 33284 16046
rect 33232 15982 33284 15988
rect 33416 15428 33468 15434
rect 33416 15370 33468 15376
rect 33048 11348 33100 11354
rect 33048 11290 33100 11296
rect 32680 11076 32732 11082
rect 32680 11018 32732 11024
rect 32692 10266 32720 11018
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32588 9648 32640 9654
rect 32588 9590 32640 9596
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 32324 8022 32352 8502
rect 32772 8084 32824 8090
rect 32772 8026 32824 8032
rect 32312 8016 32364 8022
rect 32312 7958 32364 7964
rect 32784 7002 32812 8026
rect 32772 6996 32824 7002
rect 32772 6938 32824 6944
rect 32220 5364 32272 5370
rect 32220 5306 32272 5312
rect 31668 4752 31720 4758
rect 31668 4694 31720 4700
rect 31300 4684 31352 4690
rect 31300 4626 31352 4632
rect 30196 4616 30248 4622
rect 30196 4558 30248 4564
rect 30288 4548 30340 4554
rect 30288 4490 30340 4496
rect 30300 4146 30328 4490
rect 31680 4282 31708 4694
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 32140 4146 32168 4422
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 30300 3738 30328 4082
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 31116 3460 31168 3466
rect 31116 3402 31168 3408
rect 31128 3194 31156 3402
rect 31220 3194 31248 3946
rect 31116 3188 31168 3194
rect 31116 3130 31168 3136
rect 31208 3188 31260 3194
rect 31208 3130 31260 3136
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 30748 2848 30800 2854
rect 30748 2790 30800 2796
rect 30760 2446 30788 2790
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 29460 2304 29512 2310
rect 29460 2246 29512 2252
rect 30104 2304 30156 2310
rect 30104 2246 30156 2252
rect 29472 800 29500 2246
rect 30116 800 30144 2246
rect 30760 800 30788 2382
rect 31484 2304 31536 2310
rect 31484 2246 31536 2252
rect 31496 800 31524 2246
rect 32140 800 32168 2518
rect 32232 2446 32260 5306
rect 32784 4146 32812 6938
rect 33428 5914 33456 15370
rect 34072 14618 34100 16730
rect 34440 16726 34468 17002
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34428 16720 34480 16726
rect 34428 16662 34480 16668
rect 34244 16040 34296 16046
rect 34244 15982 34296 15988
rect 34060 14612 34112 14618
rect 34060 14554 34112 14560
rect 34072 13954 34100 14554
rect 34256 14346 34284 15982
rect 34440 14634 34468 16662
rect 34796 16448 34848 16454
rect 34796 16390 34848 16396
rect 34808 15978 34836 16390
rect 35728 16046 35756 18226
rect 35808 18148 35860 18154
rect 35808 18090 35860 18096
rect 35716 16040 35768 16046
rect 35716 15982 35768 15988
rect 34796 15972 34848 15978
rect 34796 15914 34848 15920
rect 35624 15904 35676 15910
rect 35624 15846 35676 15852
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 35636 15502 35664 15846
rect 35728 15609 35756 15982
rect 35714 15600 35770 15609
rect 35714 15535 35770 15544
rect 35624 15496 35676 15502
rect 35624 15438 35676 15444
rect 35728 15162 35756 15535
rect 35716 15156 35768 15162
rect 35716 15098 35768 15104
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 34348 14606 34468 14634
rect 34716 14618 34744 14962
rect 34796 14816 34848 14822
rect 34796 14758 34848 14764
rect 34704 14612 34756 14618
rect 34244 14340 34296 14346
rect 34244 14282 34296 14288
rect 34072 13938 34192 13954
rect 34072 13932 34204 13938
rect 34072 13926 34152 13932
rect 33508 12844 33560 12850
rect 33508 12786 33560 12792
rect 33520 11150 33548 12786
rect 34072 12238 34100 13926
rect 34152 13874 34204 13880
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 34164 12782 34192 13330
rect 34256 13258 34284 14282
rect 34348 13802 34376 14606
rect 34704 14554 34756 14560
rect 34428 14544 34480 14550
rect 34428 14486 34480 14492
rect 34440 14074 34468 14486
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34808 14006 34836 14758
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34796 14000 34848 14006
rect 34796 13942 34848 13948
rect 34336 13796 34388 13802
rect 34336 13738 34388 13744
rect 34348 13394 34376 13738
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34336 13388 34388 13394
rect 34336 13330 34388 13336
rect 34244 13252 34296 13258
rect 34244 13194 34296 13200
rect 34152 12776 34204 12782
rect 34152 12718 34204 12724
rect 34060 12232 34112 12238
rect 34060 12174 34112 12180
rect 34256 12170 34284 13194
rect 34980 13184 35032 13190
rect 34980 13126 35032 13132
rect 34992 12850 35020 13126
rect 34980 12844 35032 12850
rect 34980 12786 35032 12792
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 35716 12640 35768 12646
rect 35716 12582 35768 12588
rect 34808 12374 34836 12582
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34796 12368 34848 12374
rect 34796 12310 34848 12316
rect 35728 12322 35756 12582
rect 35820 12434 35848 18090
rect 36096 17814 36124 19382
rect 36188 17882 36216 19790
rect 36280 18154 36308 24346
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36464 20806 36492 21490
rect 36452 20800 36504 20806
rect 36452 20742 36504 20748
rect 36360 19712 36412 19718
rect 36360 19654 36412 19660
rect 36372 19174 36400 19654
rect 36464 19378 36492 20742
rect 36452 19372 36504 19378
rect 36452 19314 36504 19320
rect 36360 19168 36412 19174
rect 36360 19110 36412 19116
rect 36372 18290 36400 19110
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36268 18148 36320 18154
rect 36268 18090 36320 18096
rect 36176 17876 36228 17882
rect 36176 17818 36228 17824
rect 36084 17808 36136 17814
rect 36084 17750 36136 17756
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 35912 15706 35940 17546
rect 36096 17270 36124 17750
rect 36084 17264 36136 17270
rect 36084 17206 36136 17212
rect 36372 17134 36400 18226
rect 36556 18170 36584 25162
rect 36648 21554 36676 27066
rect 36728 26240 36780 26246
rect 36728 26182 36780 26188
rect 36740 24274 36768 26182
rect 36924 25974 36952 35974
rect 37292 35894 37320 37062
rect 38028 36825 38056 37062
rect 38014 36816 38070 36825
rect 38014 36751 38070 36760
rect 38120 36378 38148 37431
rect 38212 36922 38240 38791
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 38200 36780 38252 36786
rect 38200 36722 38252 36728
rect 38108 36372 38160 36378
rect 38108 36314 38160 36320
rect 37372 36168 37424 36174
rect 37370 36136 37372 36145
rect 37424 36136 37426 36145
rect 37370 36071 37426 36080
rect 38212 35894 38240 36722
rect 37292 35866 37412 35894
rect 38212 35866 38424 35894
rect 37004 35692 37056 35698
rect 37004 35634 37056 35640
rect 37016 26926 37044 35634
rect 37280 27464 37332 27470
rect 37280 27406 37332 27412
rect 37188 27328 37240 27334
rect 37188 27270 37240 27276
rect 37200 26994 37228 27270
rect 37188 26988 37240 26994
rect 37188 26930 37240 26936
rect 37004 26920 37056 26926
rect 37004 26862 37056 26868
rect 37016 26382 37044 26862
rect 37096 26784 37148 26790
rect 37096 26726 37148 26732
rect 37108 26518 37136 26726
rect 37096 26512 37148 26518
rect 37096 26454 37148 26460
rect 37004 26376 37056 26382
rect 37004 26318 37056 26324
rect 36912 25968 36964 25974
rect 36912 25910 36964 25916
rect 37108 25906 37136 26454
rect 37096 25900 37148 25906
rect 37096 25842 37148 25848
rect 37004 25832 37056 25838
rect 37004 25774 37056 25780
rect 37016 25226 37044 25774
rect 37200 25537 37228 26930
rect 37186 25528 37242 25537
rect 37186 25463 37242 25472
rect 37292 25430 37320 27406
rect 37384 26926 37412 35866
rect 38016 35488 38068 35494
rect 38016 35430 38068 35436
rect 38028 35329 38056 35430
rect 38014 35320 38070 35329
rect 38014 35255 38070 35264
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 38028 34649 38056 34886
rect 38014 34640 38070 34649
rect 38014 34575 38070 34584
rect 38108 33992 38160 33998
rect 38106 33960 38108 33969
rect 38160 33960 38162 33969
rect 38106 33895 38162 33904
rect 38292 33856 38344 33862
rect 38292 33798 38344 33804
rect 37556 33516 37608 33522
rect 37556 33458 37608 33464
rect 37464 27396 37516 27402
rect 37464 27338 37516 27344
rect 37372 26920 37424 26926
rect 37372 26862 37424 26868
rect 37372 26784 37424 26790
rect 37372 26726 37424 26732
rect 37384 26586 37412 26726
rect 37372 26580 37424 26586
rect 37372 26522 37424 26528
rect 37370 26480 37426 26489
rect 37370 26415 37426 26424
rect 37384 26234 37412 26415
rect 37476 26382 37504 27338
rect 37464 26376 37516 26382
rect 37464 26318 37516 26324
rect 37384 26206 37504 26234
rect 37372 25696 37424 25702
rect 37372 25638 37424 25644
rect 37280 25424 37332 25430
rect 37280 25366 37332 25372
rect 37188 25288 37240 25294
rect 37188 25230 37240 25236
rect 37004 25220 37056 25226
rect 37004 25162 37056 25168
rect 37200 24614 37228 25230
rect 37280 25152 37332 25158
rect 37280 25094 37332 25100
rect 37188 24608 37240 24614
rect 37188 24550 37240 24556
rect 37200 24410 37228 24550
rect 37188 24404 37240 24410
rect 37188 24346 37240 24352
rect 37292 24342 37320 25094
rect 37280 24336 37332 24342
rect 37280 24278 37332 24284
rect 36728 24268 36780 24274
rect 36728 24210 36780 24216
rect 37384 24206 37412 25638
rect 37476 25294 37504 26206
rect 37568 26042 37596 33458
rect 38016 33312 38068 33318
rect 38014 33280 38016 33289
rect 38068 33280 38070 33289
rect 38014 33215 38070 33224
rect 38016 32768 38068 32774
rect 38016 32710 38068 32716
rect 38028 32609 38056 32710
rect 38014 32600 38070 32609
rect 38014 32535 38070 32544
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 37924 32224 37976 32230
rect 37924 32166 37976 32172
rect 37832 31340 37884 31346
rect 37832 31282 37884 31288
rect 37740 30048 37792 30054
rect 37740 29990 37792 29996
rect 37648 27872 37700 27878
rect 37648 27814 37700 27820
rect 37556 26036 37608 26042
rect 37556 25978 37608 25984
rect 37556 25900 37608 25906
rect 37556 25842 37608 25848
rect 37568 25770 37596 25842
rect 37556 25764 37608 25770
rect 37556 25706 37608 25712
rect 37464 25288 37516 25294
rect 37464 25230 37516 25236
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 37464 24744 37516 24750
rect 37464 24686 37516 24692
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 37476 22778 37504 24686
rect 37568 22982 37596 24754
rect 37556 22976 37608 22982
rect 37556 22918 37608 22924
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37372 22704 37424 22710
rect 37372 22646 37424 22652
rect 37188 22568 37240 22574
rect 37188 22510 37240 22516
rect 37200 22234 37228 22510
rect 37188 22228 37240 22234
rect 37188 22170 37240 22176
rect 37384 21690 37412 22646
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37372 21684 37424 21690
rect 37372 21626 37424 21632
rect 37476 21554 37504 22578
rect 37568 21554 37596 22918
rect 37660 22522 37688 27814
rect 37752 22642 37780 29990
rect 37844 25974 37872 31282
rect 37832 25968 37884 25974
rect 37832 25910 37884 25916
rect 37936 25906 37964 32166
rect 38120 31929 38148 32370
rect 38106 31920 38162 31929
rect 38106 31855 38162 31864
rect 38200 31816 38252 31822
rect 38200 31758 38252 31764
rect 38016 31136 38068 31142
rect 38014 31104 38016 31113
rect 38068 31104 38070 31113
rect 38014 31039 38070 31048
rect 38016 30592 38068 30598
rect 38016 30534 38068 30540
rect 38028 30433 38056 30534
rect 38014 30424 38070 30433
rect 38014 30359 38070 30368
rect 38108 30252 38160 30258
rect 38108 30194 38160 30200
rect 38120 29753 38148 30194
rect 38106 29744 38162 29753
rect 38106 29679 38162 29688
rect 38212 29594 38240 31758
rect 38120 29566 38240 29594
rect 38014 29064 38070 29073
rect 38014 28999 38016 29008
rect 38068 28999 38070 29008
rect 38016 28970 38068 28976
rect 38016 28416 38068 28422
rect 38014 28384 38016 28393
rect 38068 28384 38070 28393
rect 38014 28319 38070 28328
rect 38120 28234 38148 29566
rect 38200 29164 38252 29170
rect 38200 29106 38252 29112
rect 38028 28206 38148 28234
rect 38028 27554 38056 28206
rect 38108 28076 38160 28082
rect 38108 28018 38160 28024
rect 38120 27713 38148 28018
rect 38106 27704 38162 27713
rect 38106 27639 38162 27648
rect 38028 27526 38148 27554
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 38028 27033 38056 27270
rect 38014 27024 38070 27033
rect 38014 26959 38070 26968
rect 38016 26512 38068 26518
rect 38120 26489 38148 27526
rect 38016 26454 38068 26460
rect 38106 26480 38162 26489
rect 38028 26217 38056 26454
rect 38106 26415 38162 26424
rect 38212 26234 38240 29106
rect 38304 26382 38332 33798
rect 38396 27062 38424 35866
rect 38384 27056 38436 27062
rect 38384 26998 38436 27004
rect 38384 26784 38436 26790
rect 38384 26726 38436 26732
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38396 26234 38424 26726
rect 38014 26208 38070 26217
rect 38014 26143 38070 26152
rect 38120 26206 38240 26234
rect 38304 26206 38424 26234
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 37832 25764 37884 25770
rect 37832 25706 37884 25712
rect 37844 25294 37872 25706
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37844 24342 37872 25230
rect 38014 24848 38070 24857
rect 38014 24783 38070 24792
rect 38028 24682 38056 24783
rect 38120 24750 38148 26206
rect 38200 25968 38252 25974
rect 38200 25910 38252 25916
rect 38108 24744 38160 24750
rect 38108 24686 38160 24692
rect 38016 24676 38068 24682
rect 38016 24618 38068 24624
rect 37832 24336 37884 24342
rect 37832 24278 37884 24284
rect 38014 24168 38070 24177
rect 38014 24103 38070 24112
rect 38028 24070 38056 24103
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 38108 23724 38160 23730
rect 38108 23666 38160 23672
rect 37832 23520 37884 23526
rect 38120 23497 38148 23666
rect 37832 23462 37884 23468
rect 38106 23488 38162 23497
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 37660 22494 37780 22522
rect 37648 22092 37700 22098
rect 37648 22034 37700 22040
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 36912 21548 36964 21554
rect 36912 21490 36964 21496
rect 37004 21548 37056 21554
rect 37004 21490 37056 21496
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 36726 21312 36782 21321
rect 36726 21247 36782 21256
rect 36740 20602 36768 21247
rect 36924 21146 36952 21490
rect 37016 21418 37044 21490
rect 37004 21412 37056 21418
rect 37004 21354 37056 21360
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 37016 20942 37044 21354
rect 37372 21344 37424 21350
rect 37372 21286 37424 21292
rect 36820 20936 36872 20942
rect 36820 20878 36872 20884
rect 37004 20936 37056 20942
rect 37004 20878 37056 20884
rect 36728 20596 36780 20602
rect 36728 20538 36780 20544
rect 36556 18154 36676 18170
rect 36556 18148 36688 18154
rect 36556 18142 36636 18148
rect 36636 18090 36688 18096
rect 36360 17128 36412 17134
rect 36360 17070 36412 17076
rect 36084 16584 36136 16590
rect 36084 16526 36136 16532
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 35992 14408 36044 14414
rect 35992 14350 36044 14356
rect 35900 13932 35952 13938
rect 35900 13874 35952 13880
rect 35912 13530 35940 13874
rect 35900 13524 35952 13530
rect 35900 13466 35952 13472
rect 36004 13258 36032 14350
rect 36096 14074 36124 16526
rect 36176 16448 36228 16454
rect 36174 16416 36176 16425
rect 36228 16416 36230 16425
rect 36174 16351 36230 16360
rect 36174 14376 36230 14385
rect 36174 14311 36230 14320
rect 36188 14278 36216 14311
rect 36176 14272 36228 14278
rect 36176 14214 36228 14220
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 35820 12406 35940 12434
rect 35728 12294 35848 12322
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 34244 12164 34296 12170
rect 34244 12106 34296 12112
rect 34152 12096 34204 12102
rect 34152 12038 34204 12044
rect 34164 11830 34192 12038
rect 34152 11824 34204 11830
rect 34152 11766 34204 11772
rect 34440 11762 34468 12174
rect 35820 12170 35848 12294
rect 35808 12164 35860 12170
rect 35808 12106 35860 12112
rect 35912 12050 35940 12406
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 35820 12022 35940 12050
rect 34428 11756 34480 11762
rect 34428 11698 34480 11704
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 35820 10266 35848 12022
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 35820 9586 35848 10202
rect 34612 9580 34664 9586
rect 34612 9522 34664 9528
rect 35808 9580 35860 9586
rect 35808 9522 35860 9528
rect 34520 9376 34572 9382
rect 34520 9318 34572 9324
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33612 7546 33640 8298
rect 34072 7954 34100 8570
rect 34060 7948 34112 7954
rect 34060 7890 34112 7896
rect 33600 7540 33652 7546
rect 33600 7482 33652 7488
rect 34348 7478 34376 8910
rect 34428 8424 34480 8430
rect 34532 8378 34560 9318
rect 34480 8372 34560 8378
rect 34428 8366 34560 8372
rect 34440 8350 34560 8366
rect 34532 7818 34560 8350
rect 34520 7812 34572 7818
rect 34520 7754 34572 7760
rect 34336 7472 34388 7478
rect 34336 7414 34388 7420
rect 33416 5908 33468 5914
rect 33416 5850 33468 5856
rect 32864 5840 32916 5846
rect 32864 5782 32916 5788
rect 33428 5794 33456 5850
rect 32876 5370 32904 5782
rect 33428 5766 33548 5794
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32772 4140 32824 4146
rect 32772 4082 32824 4088
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 32324 3534 32352 3878
rect 32784 3738 32812 4082
rect 32876 3942 32904 5306
rect 33416 4616 33468 4622
rect 33416 4558 33468 4564
rect 33428 4078 33456 4558
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32784 800 32812 2994
rect 33520 2446 33548 5766
rect 34348 5370 34376 7414
rect 34532 6338 34560 7754
rect 34624 7546 34652 9522
rect 35440 9376 35492 9382
rect 35440 9318 35492 9324
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34704 9104 34756 9110
rect 34704 9046 34756 9052
rect 34716 7750 34744 9046
rect 35452 8498 35480 9318
rect 35808 8832 35860 8838
rect 35808 8774 35860 8780
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 34796 8288 34848 8294
rect 34796 8230 34848 8236
rect 34704 7744 34756 7750
rect 34704 7686 34756 7692
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34808 7274 34836 8230
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35360 8090 35388 8434
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 35360 7546 35388 8026
rect 35820 7886 35848 8774
rect 35808 7880 35860 7886
rect 35808 7822 35860 7828
rect 36096 7546 36124 11222
rect 36280 10266 36308 12174
rect 36452 11144 36504 11150
rect 36452 11086 36504 11092
rect 36464 10849 36492 11086
rect 36450 10840 36506 10849
rect 36450 10775 36506 10784
rect 36268 10260 36320 10266
rect 36268 10202 36320 10208
rect 36280 9058 36308 10202
rect 36648 10130 36676 18090
rect 36832 17882 36860 20878
rect 37016 20618 37044 20878
rect 37016 20590 37320 20618
rect 37384 20602 37412 21286
rect 37660 21010 37688 22034
rect 37648 21004 37700 21010
rect 37648 20946 37700 20952
rect 37648 20800 37700 20806
rect 37648 20742 37700 20748
rect 37292 20482 37320 20590
rect 37372 20596 37424 20602
rect 37372 20538 37424 20544
rect 37292 20466 37412 20482
rect 37660 20466 37688 20742
rect 37752 20466 37780 22494
rect 37844 21554 37872 23462
rect 38106 23423 38162 23432
rect 37924 23112 37976 23118
rect 37924 23054 37976 23060
rect 37936 22094 37964 23054
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 38028 22817 38056 22918
rect 38014 22808 38070 22817
rect 38014 22743 38070 22752
rect 38108 22636 38160 22642
rect 38108 22578 38160 22584
rect 38016 22094 38068 22098
rect 37936 22092 38068 22094
rect 37936 22066 38016 22092
rect 38016 22034 38068 22040
rect 37924 22024 37976 22030
rect 37924 21966 37976 21972
rect 38014 21992 38070 22001
rect 37936 21706 37964 21966
rect 38014 21927 38070 21936
rect 38028 21894 38056 21927
rect 38016 21888 38068 21894
rect 38016 21830 38068 21836
rect 37936 21678 38056 21706
rect 37832 21548 37884 21554
rect 37832 21490 37884 21496
rect 37924 21548 37976 21554
rect 37924 21490 37976 21496
rect 37936 21434 37964 21490
rect 37844 21406 37964 21434
rect 37844 21146 37872 21406
rect 37832 21140 37884 21146
rect 37832 21082 37884 21088
rect 37844 20942 37872 21082
rect 37832 20936 37884 20942
rect 37832 20878 37884 20884
rect 37844 20482 37872 20878
rect 37844 20466 37964 20482
rect 37292 20460 37424 20466
rect 37292 20454 37372 20460
rect 37372 20402 37424 20408
rect 37648 20460 37700 20466
rect 37648 20402 37700 20408
rect 37740 20460 37792 20466
rect 37740 20402 37792 20408
rect 37844 20460 37976 20466
rect 37844 20454 37924 20460
rect 37280 20256 37332 20262
rect 37280 20198 37332 20204
rect 37292 19990 37320 20198
rect 37280 19984 37332 19990
rect 37280 19926 37332 19932
rect 37280 19168 37332 19174
rect 37280 19110 37332 19116
rect 37292 18766 37320 19110
rect 37384 18834 37412 20402
rect 37844 18902 37872 20454
rect 37924 20402 37976 20408
rect 38028 20330 38056 21678
rect 38120 21554 38148 22578
rect 38212 22574 38240 25910
rect 38304 25770 38332 26206
rect 38292 25764 38344 25770
rect 38292 25706 38344 25712
rect 38292 24336 38344 24342
rect 38292 24278 38344 24284
rect 38200 22568 38252 22574
rect 38200 22510 38252 22516
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 38106 21312 38162 21321
rect 38106 21247 38162 21256
rect 38120 20942 38148 21247
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38016 20324 38068 20330
rect 38016 20266 38068 20272
rect 38016 19984 38068 19990
rect 38014 19952 38016 19961
rect 38068 19952 38070 19961
rect 38014 19887 38070 19896
rect 38108 19712 38160 19718
rect 38108 19654 38160 19660
rect 38120 19281 38148 19654
rect 38106 19272 38162 19281
rect 38106 19207 38162 19216
rect 38016 19168 38068 19174
rect 38016 19110 38068 19116
rect 37832 18896 37884 18902
rect 37832 18838 37884 18844
rect 37372 18828 37424 18834
rect 37372 18770 37424 18776
rect 37280 18760 37332 18766
rect 37280 18702 37332 18708
rect 37292 18086 37320 18702
rect 37372 18624 37424 18630
rect 38028 18601 38056 19110
rect 38120 18766 38148 19207
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 37372 18566 37424 18572
rect 38014 18592 38070 18601
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 36820 17876 36872 17882
rect 36820 17818 36872 17824
rect 36832 16590 36860 17818
rect 37096 17264 37148 17270
rect 37096 17206 37148 17212
rect 36820 16584 36872 16590
rect 36820 16526 36872 16532
rect 37004 16584 37056 16590
rect 37004 16526 37056 16532
rect 36820 16448 36872 16454
rect 36820 16390 36872 16396
rect 36832 14890 36860 16390
rect 37016 16114 37044 16526
rect 37004 16108 37056 16114
rect 37004 16050 37056 16056
rect 37016 15502 37044 16050
rect 37004 15496 37056 15502
rect 37004 15438 37056 15444
rect 36820 14884 36872 14890
rect 36820 14826 36872 14832
rect 37016 14414 37044 15438
rect 37108 15434 37136 17206
rect 37292 17202 37320 18022
rect 37188 17196 37240 17202
rect 37188 17138 37240 17144
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37200 16590 37228 17138
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 37200 15502 37228 16526
rect 37292 16046 37320 17138
rect 37384 16590 37412 18566
rect 38014 18527 38070 18536
rect 38016 18080 38068 18086
rect 38016 18022 38068 18028
rect 38028 17785 38056 18022
rect 38014 17776 38070 17785
rect 38014 17711 38070 17720
rect 38304 17270 38332 24278
rect 38384 22772 38436 22778
rect 38384 22714 38436 22720
rect 38396 20534 38424 22714
rect 38384 20528 38436 20534
rect 38384 20470 38436 20476
rect 38292 17264 38344 17270
rect 38292 17206 38344 17212
rect 38106 17096 38162 17105
rect 38106 17031 38162 17040
rect 38120 16590 38148 17031
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37648 16584 37700 16590
rect 37648 16526 37700 16532
rect 38108 16584 38160 16590
rect 38108 16526 38160 16532
rect 37372 16448 37424 16454
rect 37372 16390 37424 16396
rect 37280 16040 37332 16046
rect 37280 15982 37332 15988
rect 37188 15496 37240 15502
rect 37188 15438 37240 15444
rect 37096 15428 37148 15434
rect 37096 15370 37148 15376
rect 37200 14414 37228 15438
rect 37292 15094 37320 15982
rect 37384 15502 37412 16390
rect 37476 15978 37504 16526
rect 37464 15972 37516 15978
rect 37464 15914 37516 15920
rect 37476 15502 37504 15914
rect 37372 15496 37424 15502
rect 37372 15438 37424 15444
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37372 15360 37424 15366
rect 37372 15302 37424 15308
rect 37280 15088 37332 15094
rect 37280 15030 37332 15036
rect 37384 14414 37412 15302
rect 37476 14414 37504 15438
rect 37660 15162 37688 16526
rect 38014 15736 38070 15745
rect 38014 15671 38070 15680
rect 38028 15162 38056 15671
rect 38108 15496 38160 15502
rect 38108 15438 38160 15444
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 38120 15065 38148 15438
rect 38106 15056 38162 15065
rect 38106 14991 38162 15000
rect 38120 14618 38148 14991
rect 38108 14612 38160 14618
rect 38108 14554 38160 14560
rect 37004 14408 37056 14414
rect 37004 14350 37056 14356
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 37372 14408 37424 14414
rect 37372 14350 37424 14356
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 37016 13326 37044 14350
rect 37096 14340 37148 14346
rect 37096 14282 37148 14288
rect 37108 14074 37136 14282
rect 37096 14068 37148 14074
rect 37096 14010 37148 14016
rect 37200 13326 37228 14350
rect 37280 14340 37332 14346
rect 37280 14282 37332 14288
rect 37292 13394 37320 14282
rect 38016 13728 38068 13734
rect 38014 13696 38016 13705
rect 38068 13696 38070 13705
rect 38014 13631 38070 13640
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 37004 13320 37056 13326
rect 37188 13320 37240 13326
rect 37004 13262 37056 13268
rect 37108 13268 37188 13274
rect 37108 13262 37240 13268
rect 36820 13184 36872 13190
rect 36820 13126 36872 13132
rect 36912 13184 36964 13190
rect 36912 13126 36964 13132
rect 36832 12753 36860 13126
rect 36818 12744 36874 12753
rect 36818 12679 36874 12688
rect 36924 12442 36952 13126
rect 36912 12436 36964 12442
rect 36912 12378 36964 12384
rect 37016 11898 37044 13262
rect 37108 13246 37228 13262
rect 37004 11892 37056 11898
rect 37004 11834 37056 11840
rect 37108 11830 37136 13246
rect 37188 12776 37240 12782
rect 37188 12718 37240 12724
rect 37096 11824 37148 11830
rect 37096 11766 37148 11772
rect 37200 11694 37228 12718
rect 37292 11762 37320 13330
rect 38108 13320 38160 13326
rect 38108 13262 38160 13268
rect 38120 12986 38148 13262
rect 38108 12980 38160 12986
rect 38108 12922 38160 12928
rect 38120 12889 38148 12922
rect 38106 12880 38162 12889
rect 38106 12815 38162 12824
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 38028 12209 38056 12582
rect 38014 12200 38070 12209
rect 38014 12135 38070 12144
rect 37280 11756 37332 11762
rect 37280 11698 37332 11704
rect 37372 11756 37424 11762
rect 37372 11698 37424 11704
rect 37188 11688 37240 11694
rect 37188 11630 37240 11636
rect 37384 11354 37412 11698
rect 38014 11520 38070 11529
rect 38014 11455 38070 11464
rect 38028 11354 38056 11455
rect 37372 11348 37424 11354
rect 37372 11290 37424 11296
rect 38016 11348 38068 11354
rect 38016 11290 38068 11296
rect 37188 11280 37240 11286
rect 37188 11222 37240 11228
rect 37200 10169 37228 11222
rect 37648 11144 37700 11150
rect 37648 11086 37700 11092
rect 37280 10804 37332 10810
rect 37280 10746 37332 10752
rect 37186 10160 37242 10169
rect 36636 10124 36688 10130
rect 37186 10095 37242 10104
rect 36636 10066 36688 10072
rect 37292 9586 37320 10746
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37556 9512 37608 9518
rect 37556 9454 37608 9460
rect 37372 9444 37424 9450
rect 37372 9386 37424 9392
rect 36188 9030 36308 9058
rect 36188 8974 36216 9030
rect 36176 8968 36228 8974
rect 36176 8910 36228 8916
rect 36188 8566 36216 8910
rect 36360 8900 36412 8906
rect 36360 8842 36412 8848
rect 36176 8560 36228 8566
rect 36176 8502 36228 8508
rect 36372 8090 36400 8842
rect 37384 8634 37412 9386
rect 37464 9172 37516 9178
rect 37464 9114 37516 9120
rect 36728 8628 36780 8634
rect 36728 8570 36780 8576
rect 37372 8628 37424 8634
rect 37372 8570 37424 8576
rect 36360 8084 36412 8090
rect 36360 8026 36412 8032
rect 36740 7886 36768 8570
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 35348 7540 35400 7546
rect 35348 7482 35400 7488
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 36084 7540 36136 7546
rect 36084 7482 36136 7488
rect 34796 7268 34848 7274
rect 34796 7210 34848 7216
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34532 6310 34652 6338
rect 34520 6180 34572 6186
rect 34520 6122 34572 6128
rect 34532 5710 34560 6122
rect 34624 5778 34652 6310
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34612 5772 34664 5778
rect 34612 5714 34664 5720
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34428 5568 34480 5574
rect 34428 5510 34480 5516
rect 34336 5364 34388 5370
rect 34336 5306 34388 5312
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33612 4010 33640 4966
rect 34348 4690 34376 5306
rect 33876 4684 33928 4690
rect 33876 4626 33928 4632
rect 34336 4684 34388 4690
rect 34336 4626 34388 4632
rect 33888 4078 33916 4626
rect 34440 4486 34468 5510
rect 34624 5166 34652 5714
rect 34612 5160 34664 5166
rect 34612 5102 34664 5108
rect 34624 4690 34652 5102
rect 34612 4684 34664 4690
rect 34612 4626 34664 4632
rect 34612 4548 34664 4554
rect 34612 4490 34664 4496
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 34428 4480 34480 4486
rect 34428 4422 34480 4428
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33600 4004 33652 4010
rect 33600 3946 33652 3952
rect 33980 3534 34008 4422
rect 34440 4214 34468 4422
rect 34428 4208 34480 4214
rect 34428 4150 34480 4156
rect 34624 4146 34652 4490
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34152 3664 34204 3670
rect 34152 3606 34204 3612
rect 33968 3528 34020 3534
rect 33968 3470 34020 3476
rect 34164 3466 34192 3606
rect 34152 3460 34204 3466
rect 34152 3402 34204 3408
rect 34716 3058 34744 6190
rect 34808 4826 34836 6258
rect 35624 6112 35676 6118
rect 35624 6054 35676 6060
rect 35716 6112 35768 6118
rect 35716 6054 35768 6060
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35440 5568 35492 5574
rect 35440 5510 35492 5516
rect 35452 5098 35480 5510
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 35440 5092 35492 5098
rect 35440 5034 35492 5040
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34796 4820 34848 4826
rect 34796 4762 34848 4768
rect 35544 4282 35572 5170
rect 35532 4276 35584 4282
rect 35532 4218 35584 4224
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34704 3052 34756 3058
rect 34704 2994 34756 3000
rect 34808 2632 34836 3062
rect 35072 2984 35124 2990
rect 35256 2984 35308 2990
rect 35124 2944 35256 2972
rect 35072 2926 35124 2932
rect 35256 2926 35308 2932
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34808 2604 34928 2632
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 32876 1970 32904 2382
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 32864 1964 32916 1970
rect 32864 1906 32916 1912
rect 33520 800 33548 2246
rect 34164 800 34192 2246
rect 34900 800 34928 2604
rect 35636 2446 35664 6054
rect 35728 5710 35756 6054
rect 35716 5704 35768 5710
rect 35716 5646 35768 5652
rect 35728 4457 35756 5646
rect 35820 5522 35848 7482
rect 35820 5494 35940 5522
rect 35912 4690 35940 5494
rect 35900 4684 35952 4690
rect 35900 4626 35952 4632
rect 36096 4570 36124 7482
rect 37200 7478 37228 7822
rect 37188 7472 37240 7478
rect 37188 7414 37240 7420
rect 36636 7336 36688 7342
rect 36636 7278 36688 7284
rect 37370 7304 37426 7313
rect 36648 7002 36676 7278
rect 37370 7239 37372 7248
rect 37424 7239 37426 7248
rect 37372 7210 37424 7216
rect 36636 6996 36688 7002
rect 36636 6938 36688 6944
rect 36452 6792 36504 6798
rect 36452 6734 36504 6740
rect 37096 6792 37148 6798
rect 37096 6734 37148 6740
rect 36464 6633 36492 6734
rect 36450 6624 36506 6633
rect 36450 6559 36506 6568
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 36832 5914 36860 6394
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 37108 5710 37136 6734
rect 37280 6656 37332 6662
rect 37280 6598 37332 6604
rect 37188 6180 37240 6186
rect 37188 6122 37240 6128
rect 37096 5704 37148 5710
rect 36924 5652 37096 5658
rect 36924 5646 37148 5652
rect 36924 5642 37136 5646
rect 36912 5636 37136 5642
rect 36964 5630 37136 5636
rect 36912 5578 36964 5584
rect 36268 5024 36320 5030
rect 36268 4966 36320 4972
rect 36280 4622 36308 4966
rect 37108 4826 37136 5630
rect 37096 4820 37148 4826
rect 37096 4762 37148 4768
rect 36360 4684 36412 4690
rect 36360 4626 36412 4632
rect 36268 4616 36320 4622
rect 36096 4542 36216 4570
rect 36268 4558 36320 4564
rect 36084 4480 36136 4486
rect 35714 4448 35770 4457
rect 36084 4422 36136 4428
rect 35714 4383 35770 4392
rect 36096 4078 36124 4422
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 35716 3936 35768 3942
rect 35716 3878 35768 3884
rect 35728 3058 35756 3878
rect 36096 3738 36124 4014
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 35716 3052 35768 3058
rect 35716 2994 35768 3000
rect 36096 2446 36124 3674
rect 36188 3058 36216 4542
rect 36372 3738 36400 4626
rect 36636 3936 36688 3942
rect 36636 3878 36688 3884
rect 36648 3777 36676 3878
rect 36634 3768 36690 3777
rect 36360 3732 36412 3738
rect 36634 3703 36690 3712
rect 36360 3674 36412 3680
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 35532 2304 35584 2310
rect 35532 2246 35584 2252
rect 35544 800 35572 2246
rect 36188 800 36216 2790
rect 37200 2514 37228 6122
rect 37292 5953 37320 6598
rect 37278 5944 37334 5953
rect 37278 5879 37334 5888
rect 37370 5128 37426 5137
rect 37370 5063 37372 5072
rect 37424 5063 37426 5072
rect 37372 5034 37424 5040
rect 37370 4040 37426 4049
rect 37476 4026 37504 9114
rect 37568 8498 37596 9454
rect 37660 8838 37688 11086
rect 38304 10810 38332 17206
rect 38292 10804 38344 10810
rect 38292 10746 38344 10752
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 37740 10056 37792 10062
rect 37740 9998 37792 10004
rect 37648 8832 37700 8838
rect 37648 8774 37700 8780
rect 37660 8498 37688 8774
rect 37752 8566 37780 9998
rect 38028 9489 38056 10406
rect 38014 9480 38070 9489
rect 38014 9415 38070 9424
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 37924 8832 37976 8838
rect 37924 8774 37976 8780
rect 37740 8560 37792 8566
rect 37740 8502 37792 8508
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 37568 7410 37596 8434
rect 37660 7750 37688 8434
rect 37648 7744 37700 7750
rect 37648 7686 37700 7692
rect 37752 7478 37780 8502
rect 37936 8498 37964 8774
rect 38028 8498 38056 9318
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8673 38148 8910
rect 38106 8664 38162 8673
rect 38106 8599 38162 8608
rect 37924 8492 37976 8498
rect 37924 8434 37976 8440
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 38028 8242 38056 8434
rect 37936 8214 38056 8242
rect 37740 7472 37792 7478
rect 37740 7414 37792 7420
rect 37936 7426 37964 8214
rect 38016 8084 38068 8090
rect 38016 8026 38068 8032
rect 38028 7993 38056 8026
rect 38014 7984 38070 7993
rect 38120 7954 38148 8599
rect 38936 8016 38988 8022
rect 38936 7958 38988 7964
rect 38014 7919 38070 7928
rect 38108 7948 38160 7954
rect 38108 7890 38160 7896
rect 37556 7404 37608 7410
rect 37556 7346 37608 7352
rect 37568 5574 37596 7346
rect 37752 5642 37780 7414
rect 37936 7410 38056 7426
rect 37936 7404 38068 7410
rect 37936 7398 38016 7404
rect 37936 5710 37964 7398
rect 38016 7346 38068 7352
rect 38014 7304 38070 7313
rect 38014 7239 38070 7248
rect 38028 7002 38056 7239
rect 38016 6996 38068 7002
rect 38016 6938 38068 6944
rect 38108 6180 38160 6186
rect 38108 6122 38160 6128
rect 38016 6112 38068 6118
rect 38016 6054 38068 6060
rect 37924 5704 37976 5710
rect 37844 5652 37924 5658
rect 37844 5646 37976 5652
rect 37740 5636 37792 5642
rect 37740 5578 37792 5584
rect 37844 5630 37964 5646
rect 37556 5568 37608 5574
rect 37556 5510 37608 5516
rect 37568 5234 37596 5510
rect 37752 5302 37780 5578
rect 37844 5370 37872 5630
rect 37924 5568 37976 5574
rect 37924 5510 37976 5516
rect 37832 5364 37884 5370
rect 37832 5306 37884 5312
rect 37740 5296 37792 5302
rect 37740 5238 37792 5244
rect 37556 5228 37608 5234
rect 37556 5170 37608 5176
rect 37568 4146 37596 5170
rect 37752 4214 37780 5238
rect 37844 4282 37872 5306
rect 37936 5234 37964 5510
rect 38028 5273 38056 6054
rect 38120 5710 38148 6122
rect 38108 5704 38160 5710
rect 38108 5646 38160 5652
rect 38014 5264 38070 5273
rect 37924 5228 37976 5234
rect 38014 5199 38070 5208
rect 37924 5170 37976 5176
rect 37832 4276 37884 4282
rect 37832 4218 37884 4224
rect 37740 4208 37792 4214
rect 37740 4150 37792 4156
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37476 3998 37688 4026
rect 37370 3975 37372 3984
rect 37424 3975 37426 3984
rect 37372 3946 37424 3952
rect 37280 3392 37332 3398
rect 37280 3334 37332 3340
rect 37292 3097 37320 3334
rect 37278 3088 37334 3097
rect 37278 3023 37334 3032
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 37188 2508 37240 2514
rect 37188 2450 37240 2456
rect 36636 2304 36688 2310
rect 36636 2246 36688 2252
rect 36648 1737 36676 2246
rect 36634 1728 36690 1737
rect 36634 1663 36690 1672
rect 36924 800 36952 2450
rect 5724 264 5776 270
rect 5724 206 5776 212
rect 6366 0 6422 800
rect 7010 0 7066 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9770 0 9826 800
rect 10414 0 10470 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 13174 0 13230 800
rect 13818 0 13874 800
rect 14462 0 14518 800
rect 15198 0 15254 800
rect 15842 0 15898 800
rect 16486 0 16542 800
rect 17222 0 17278 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19246 0 19302 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22650 0 22706 800
rect 23294 0 23350 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 26054 0 26110 800
rect 26698 0 26754 800
rect 27342 0 27398 800
rect 28078 0 28134 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30102 0 30158 800
rect 30746 0 30802 800
rect 31482 0 31538 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34886 0 34942 800
rect 35530 0 35586 800
rect 36174 0 36230 800
rect 36910 0 36966 800
rect 37384 377 37412 2926
rect 37660 2922 37688 3998
rect 37844 3126 37872 4082
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 37832 3120 37884 3126
rect 37832 3062 37884 3068
rect 37464 2916 37516 2922
rect 37464 2858 37516 2864
rect 37648 2916 37700 2922
rect 37648 2858 37700 2864
rect 37476 1442 37504 2858
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37568 2106 37596 2382
rect 37556 2100 37608 2106
rect 37556 2042 37608 2048
rect 37476 1414 37596 1442
rect 37568 800 37596 1414
rect 38028 1057 38056 3334
rect 38120 2417 38148 5646
rect 38200 3188 38252 3194
rect 38200 3130 38252 3136
rect 38106 2408 38162 2417
rect 38106 2343 38162 2352
rect 38014 1048 38070 1057
rect 38014 983 38070 992
rect 38212 800 38240 3130
rect 38948 800 38976 7958
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 39592 800 39620 2994
rect 37370 368 37426 377
rect 37370 303 37426 312
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38934 0 38990 800
rect 39578 0 39634 800
<< via2 >>
rect 2870 39616 2926 39672
rect 2778 38800 2834 38856
rect 1490 37848 1546 37904
rect 1398 37032 1454 37088
rect 35714 39480 35770 39536
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 38198 38800 38254 38856
rect 35806 38120 35862 38176
rect 38106 37440 38162 37496
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 1398 36116 1400 36136
rect 1400 36116 1452 36136
rect 1452 36116 1454 36136
rect 1398 36080 1454 36116
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 1398 35264 1454 35320
rect 1398 34468 1454 34504
rect 1398 34448 1400 34468
rect 1400 34448 1452 34468
rect 1452 34448 1454 34468
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 1398 33496 1454 33552
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 1398 32680 1454 32736
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1490 31728 1546 31784
rect 1398 31320 1454 31376
rect 1398 30368 1454 30424
rect 1398 29996 1400 30016
rect 1400 29996 1452 30016
rect 1452 29996 1454 30016
rect 1398 29960 1454 29996
rect 1398 29144 1454 29200
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 1398 28736 1454 28792
rect 1398 27784 1454 27840
rect 1398 27412 1400 27432
rect 1400 27412 1452 27432
rect 1452 27412 1454 27432
rect 1398 27376 1454 27412
rect 1398 26424 1454 26480
rect 1490 26016 1546 26072
rect 1398 25608 1454 25664
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1490 24656 1546 24712
rect 1858 24248 1914 24304
rect 2134 23840 2190 23896
rect 1490 23468 1492 23488
rect 1492 23468 1544 23488
rect 1544 23468 1546 23488
rect 1490 23432 1546 23468
rect 1858 23044 1914 23080
rect 1858 23024 1860 23044
rect 1860 23024 1912 23044
rect 1912 23024 1914 23044
rect 2134 22480 2190 22536
rect 1490 22072 1546 22128
rect 1858 21664 1914 21720
rect 1398 21256 1454 21312
rect 1490 20748 1492 20768
rect 1492 20748 1544 20768
rect 1544 20748 1546 20768
rect 1490 20712 1546 20748
rect 1858 20304 1914 20360
rect 1490 19488 1546 19544
rect 1858 18944 1914 19000
rect 1398 18536 1454 18592
rect 2778 19896 2834 19952
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1490 18128 1546 18184
rect 1858 17720 1914 17776
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 2134 17332 2190 17368
rect 2134 17312 2136 17332
rect 2136 17312 2188 17332
rect 2188 17312 2190 17332
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 6274 17720 6330 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 1490 16768 1546 16824
rect 1858 16360 1914 16416
rect 1674 16108 1730 16144
rect 1674 16088 1676 16108
rect 1676 16088 1728 16108
rect 1728 16088 1730 16108
rect 2134 15952 2190 16008
rect 1490 15544 1546 15600
rect 1858 15000 1914 15056
rect 1398 14592 1454 14648
rect 1674 14456 1730 14512
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1398 13776 1454 13832
rect 1674 13368 1730 13424
rect 2134 13268 2136 13288
rect 2136 13268 2188 13288
rect 2188 13268 2190 13288
rect 2134 13232 2190 13268
rect 1490 12824 1546 12880
rect 1858 12416 1914 12472
rect 1398 12008 1454 12064
rect 1490 11620 1546 11656
rect 1490 11600 1492 11620
rect 1492 11600 1544 11620
rect 1544 11600 1546 11620
rect 1858 11092 1860 11112
rect 1860 11092 1912 11112
rect 1912 11092 1914 11112
rect 1858 11056 1914 11092
rect 1490 10240 1546 10296
rect 1858 9832 1914 9888
rect 2042 9288 2098 9344
rect 1490 8880 1546 8936
rect 1398 8064 1454 8120
rect 1490 7520 1546 7576
rect 1398 7112 1454 7168
rect 1490 6296 1546 6352
rect 1398 3168 1454 3224
rect 1674 5652 1676 5672
rect 1676 5652 1728 5672
rect 1728 5652 1730 5672
rect 1674 5616 1730 5652
rect 1582 4120 1638 4176
rect 2042 6740 2044 6760
rect 2044 6740 2096 6760
rect 2096 6740 2098 6760
rect 2042 6704 2098 6740
rect 1858 5888 1914 5944
rect 1858 4548 1914 4584
rect 1858 4528 1860 4548
rect 1860 4528 1912 4548
rect 1912 4528 1914 4548
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 2870 10648 2926 10704
rect 2778 8880 2834 8936
rect 2778 8472 2834 8528
rect 2962 8880 3018 8936
rect 1490 2352 1546 2408
rect 2870 5344 2926 5400
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 2962 4936 3018 4992
rect 3238 4664 3294 4720
rect 2778 3576 2834 3632
rect 2870 1808 2926 1864
rect 2778 1400 2834 1456
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4066 4664 4122 4720
rect 4250 4684 4306 4720
rect 4250 4664 4252 4684
rect 4252 4664 4304 4684
rect 4304 4664 4306 4684
rect 3514 2760 3570 2816
rect 3330 992 3386 1048
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3974 584 4030 640
rect 3974 212 3976 232
rect 3976 212 4028 232
rect 4028 212 4030 232
rect 3974 176 4030 212
rect 7010 16516 7066 16552
rect 7010 16496 7012 16516
rect 7012 16496 7064 16516
rect 7064 16496 7066 16516
rect 7562 17604 7618 17640
rect 7562 17584 7564 17604
rect 7564 17584 7616 17604
rect 7616 17584 7618 17604
rect 7746 17076 7748 17096
rect 7748 17076 7800 17096
rect 7800 17076 7802 17096
rect 7746 17040 7802 17076
rect 11150 17448 11206 17504
rect 10690 13268 10692 13288
rect 10692 13268 10744 13288
rect 10744 13268 10746 13288
rect 10690 13232 10746 13268
rect 9678 3304 9734 3360
rect 10322 3848 10378 3904
rect 10322 3460 10378 3496
rect 10322 3440 10324 3460
rect 10324 3440 10376 3460
rect 10376 3440 10378 3460
rect 10782 3304 10838 3360
rect 10966 3440 11022 3496
rect 11978 8916 11980 8936
rect 11980 8916 12032 8936
rect 12032 8916 12034 8936
rect 11978 8880 12034 8916
rect 12070 8744 12126 8800
rect 12806 15564 12862 15600
rect 12806 15544 12808 15564
rect 12808 15544 12860 15564
rect 12860 15544 12862 15564
rect 13726 19216 13782 19272
rect 13358 17448 13414 17504
rect 12254 5752 12310 5808
rect 12254 5228 12310 5264
rect 12254 5208 12256 5228
rect 12256 5208 12308 5228
rect 12308 5208 12310 5228
rect 14186 17720 14242 17776
rect 13358 13932 13414 13968
rect 13358 13912 13360 13932
rect 13360 13912 13412 13932
rect 13412 13912 13414 13932
rect 12806 7248 12862 7304
rect 13358 8916 13360 8936
rect 13360 8916 13412 8936
rect 13412 8916 13414 8936
rect 13358 8880 13414 8916
rect 12898 5616 12954 5672
rect 12714 5072 12770 5128
rect 13174 4936 13230 4992
rect 11794 3476 11796 3496
rect 11796 3476 11848 3496
rect 11848 3476 11850 3496
rect 11794 3440 11850 3476
rect 12898 3732 12954 3768
rect 12898 3712 12900 3732
rect 12900 3712 12952 3732
rect 12952 3712 12954 3732
rect 13358 3984 13414 4040
rect 14830 14320 14886 14376
rect 14462 6604 14464 6624
rect 14464 6604 14516 6624
rect 14516 6604 14518 6624
rect 14462 6568 14518 6604
rect 15474 13232 15530 13288
rect 15198 4528 15254 4584
rect 16302 6740 16304 6760
rect 16304 6740 16356 6760
rect 16356 6740 16358 6760
rect 16302 6704 16358 6740
rect 16210 4800 16266 4856
rect 17314 15000 17370 15056
rect 17406 14728 17462 14784
rect 17038 13368 17094 13424
rect 17774 14456 17830 14512
rect 18050 14864 18106 14920
rect 17958 14728 18014 14784
rect 17222 8744 17278 8800
rect 17498 6740 17500 6760
rect 17500 6740 17552 6760
rect 17552 6740 17554 6760
rect 17498 6704 17554 6740
rect 17774 14340 17830 14376
rect 17774 14320 17776 14340
rect 17776 14320 17828 14340
rect 17828 14320 17830 14340
rect 16854 4564 16856 4584
rect 16856 4564 16908 4584
rect 16908 4564 16910 4584
rect 16854 4528 16910 4564
rect 17866 13812 17868 13832
rect 17868 13812 17920 13832
rect 17920 13812 17922 13832
rect 17866 13776 17922 13812
rect 17866 12724 17868 12744
rect 17868 12724 17920 12744
rect 17920 12724 17922 12744
rect 17866 12688 17922 12724
rect 18510 16088 18566 16144
rect 17774 6568 17830 6624
rect 17958 6704 18014 6760
rect 18602 15000 18658 15056
rect 18786 14884 18842 14920
rect 18786 14864 18788 14884
rect 18788 14864 18840 14884
rect 18840 14864 18842 14884
rect 18510 13912 18566 13968
rect 19062 17186 19118 17232
rect 19062 17176 19064 17186
rect 19064 17176 19116 17186
rect 19116 17176 19118 17186
rect 18970 14728 19026 14784
rect 18602 4820 18658 4856
rect 18602 4800 18604 4820
rect 18604 4800 18656 4820
rect 18656 4800 18658 4820
rect 17774 3884 17776 3904
rect 17776 3884 17828 3904
rect 17828 3884 17830 3904
rect 17774 3848 17830 3884
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19982 18808 20038 18864
rect 19706 18692 19762 18728
rect 19706 18672 19708 18692
rect 19708 18672 19760 18692
rect 19760 18672 19762 18692
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19338 18028 19340 18048
rect 19340 18028 19392 18048
rect 19392 18028 19394 18048
rect 19338 17992 19394 18028
rect 19614 18164 19616 18184
rect 19616 18164 19668 18184
rect 19668 18164 19670 18184
rect 19614 18128 19670 18164
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19246 17212 19248 17232
rect 19248 17212 19300 17232
rect 19300 17212 19302 17232
rect 19246 17176 19302 17212
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 20166 18808 20222 18864
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20350 18672 20406 18728
rect 20626 17992 20682 18048
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19062 3712 19118 3768
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21454 18672 21510 18728
rect 21362 18128 21418 18184
rect 22466 16108 22522 16144
rect 22466 16088 22468 16108
rect 22468 16088 22520 16108
rect 22520 16088 22522 16108
rect 22926 19236 22982 19272
rect 22926 19216 22928 19236
rect 22928 19216 22980 19236
rect 22980 19216 22982 19236
rect 22834 16088 22890 16144
rect 24766 21936 24822 21992
rect 26146 5752 26202 5808
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 27802 21936 27858 21992
rect 27618 16496 27674 16552
rect 28998 13776 29054 13832
rect 27434 5208 27490 5264
rect 26790 4936 26846 4992
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 31850 17040 31906 17096
rect 29826 4664 29882 4720
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 36174 20576 36230 20632
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35346 17584 35402 17640
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35714 15544 35770 15600
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38014 36760 38070 36816
rect 37370 36116 37372 36136
rect 37372 36116 37424 36136
rect 37424 36116 37426 36136
rect 37370 36080 37426 36116
rect 37186 25472 37242 25528
rect 38014 35264 38070 35320
rect 38014 34584 38070 34640
rect 38106 33940 38108 33960
rect 38108 33940 38160 33960
rect 38160 33940 38162 33960
rect 38106 33904 38162 33940
rect 37370 26424 37426 26480
rect 38014 33260 38016 33280
rect 38016 33260 38068 33280
rect 38068 33260 38070 33280
rect 38014 33224 38070 33260
rect 38014 32544 38070 32600
rect 38106 31864 38162 31920
rect 38014 31084 38016 31104
rect 38016 31084 38068 31104
rect 38068 31084 38070 31104
rect 38014 31048 38070 31084
rect 38014 30368 38070 30424
rect 38106 29688 38162 29744
rect 38014 29028 38070 29064
rect 38014 29008 38016 29028
rect 38016 29008 38068 29028
rect 38068 29008 38070 29028
rect 38014 28364 38016 28384
rect 38016 28364 38068 28384
rect 38068 28364 38070 28384
rect 38014 28328 38070 28364
rect 38106 27648 38162 27704
rect 38014 26968 38070 27024
rect 38106 26424 38162 26480
rect 38014 26152 38070 26208
rect 38014 24792 38070 24848
rect 38014 24112 38070 24168
rect 36726 21256 36782 21312
rect 36174 16396 36176 16416
rect 36176 16396 36228 16416
rect 36228 16396 36230 16416
rect 36174 16360 36230 16396
rect 36174 14320 36230 14376
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 36450 10784 36506 10840
rect 38106 23432 38162 23488
rect 38014 22752 38070 22808
rect 38014 21936 38070 21992
rect 38106 21256 38162 21312
rect 38014 19932 38016 19952
rect 38016 19932 38068 19952
rect 38068 19932 38070 19952
rect 38014 19896 38070 19932
rect 38106 19216 38162 19272
rect 38014 18536 38070 18592
rect 38014 17720 38070 17776
rect 38106 17040 38162 17096
rect 38014 15680 38070 15736
rect 38106 15000 38162 15056
rect 38014 13676 38016 13696
rect 38016 13676 38068 13696
rect 38068 13676 38070 13696
rect 38014 13640 38070 13676
rect 36818 12688 36874 12744
rect 38106 12824 38162 12880
rect 38014 12144 38070 12200
rect 38014 11464 38070 11520
rect 37186 10104 37242 10160
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37370 7268 37426 7304
rect 37370 7248 37372 7268
rect 37372 7248 37424 7268
rect 37424 7248 37426 7268
rect 36450 6568 36506 6624
rect 35714 4392 35770 4448
rect 36634 3712 36690 3768
rect 37278 5888 37334 5944
rect 37370 5092 37426 5128
rect 37370 5072 37372 5092
rect 37372 5072 37424 5092
rect 37424 5072 37426 5092
rect 37370 4004 37426 4040
rect 37370 3984 37372 4004
rect 37372 3984 37424 4004
rect 37424 3984 37426 4004
rect 38014 9424 38070 9480
rect 38106 8608 38162 8664
rect 38014 7928 38070 7984
rect 38014 7248 38070 7304
rect 38014 5208 38070 5264
rect 37278 3032 37334 3088
rect 36634 1672 36690 1728
rect 38106 2352 38162 2408
rect 38014 992 38070 1048
rect 37370 312 37426 368
<< metal3 >>
rect 0 39674 800 39704
rect 2865 39674 2931 39677
rect 0 39672 2931 39674
rect 0 39616 2870 39672
rect 2926 39616 2931 39672
rect 0 39614 2931 39616
rect 0 39584 800 39614
rect 2865 39611 2931 39614
rect 35709 39538 35775 39541
rect 39200 39538 40000 39568
rect 35709 39536 40000 39538
rect 35709 39480 35714 39536
rect 35770 39480 40000 39536
rect 35709 39478 40000 39480
rect 35709 39475 35775 39478
rect 39200 39448 40000 39478
rect 0 39176 800 39296
rect 0 38858 800 38888
rect 2773 38858 2839 38861
rect 0 38856 2839 38858
rect 0 38800 2778 38856
rect 2834 38800 2839 38856
rect 0 38798 2839 38800
rect 0 38768 800 38798
rect 2773 38795 2839 38798
rect 38193 38858 38259 38861
rect 39200 38858 40000 38888
rect 38193 38856 40000 38858
rect 38193 38800 38198 38856
rect 38254 38800 40000 38856
rect 38193 38798 40000 38800
rect 38193 38795 38259 38798
rect 39200 38768 40000 38798
rect 0 38360 800 38480
rect 35801 38178 35867 38181
rect 39200 38178 40000 38208
rect 35801 38176 40000 38178
rect 35801 38120 35806 38176
rect 35862 38120 40000 38176
rect 35801 38118 40000 38120
rect 35801 38115 35867 38118
rect 39200 38088 40000 38118
rect 0 37906 800 37936
rect 1485 37906 1551 37909
rect 0 37904 1551 37906
rect 0 37848 1490 37904
rect 1546 37848 1551 37904
rect 0 37846 1551 37848
rect 0 37816 800 37846
rect 1485 37843 1551 37846
rect 4208 37568 4528 37569
rect 0 37408 800 37528
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 38101 37498 38167 37501
rect 39200 37498 40000 37528
rect 38101 37496 40000 37498
rect 38101 37440 38106 37496
rect 38162 37440 40000 37496
rect 38101 37438 40000 37440
rect 38101 37435 38167 37438
rect 39200 37408 40000 37438
rect 0 37090 800 37120
rect 1393 37090 1459 37093
rect 0 37088 1459 37090
rect 0 37032 1398 37088
rect 1454 37032 1459 37088
rect 0 37030 1459 37032
rect 0 37000 800 37030
rect 1393 37027 1459 37030
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 38009 36818 38075 36821
rect 39200 36818 40000 36848
rect 38009 36816 40000 36818
rect 38009 36760 38014 36816
rect 38070 36760 40000 36816
rect 38009 36758 40000 36760
rect 38009 36755 38075 36758
rect 39200 36728 40000 36758
rect 0 36592 800 36712
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 1393 36138 1459 36141
rect 0 36136 1459 36138
rect 0 36080 1398 36136
rect 1454 36080 1459 36136
rect 0 36078 1459 36080
rect 0 36048 800 36078
rect 1393 36075 1459 36078
rect 37365 36138 37431 36141
rect 39200 36138 40000 36168
rect 37365 36136 40000 36138
rect 37365 36080 37370 36136
rect 37426 36080 40000 36136
rect 37365 36078 40000 36080
rect 37365 36075 37431 36078
rect 39200 36048 40000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35640 800 35760
rect 4208 35392 4528 35393
rect 0 35322 800 35352
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 1393 35322 1459 35325
rect 0 35320 1459 35322
rect 0 35264 1398 35320
rect 1454 35264 1459 35320
rect 0 35262 1459 35264
rect 0 35232 800 35262
rect 1393 35259 1459 35262
rect 38009 35322 38075 35325
rect 39200 35322 40000 35352
rect 38009 35320 40000 35322
rect 38009 35264 38014 35320
rect 38070 35264 40000 35320
rect 38009 35262 40000 35264
rect 38009 35259 38075 35262
rect 39200 35232 40000 35262
rect 0 34824 800 34944
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 38009 34642 38075 34645
rect 39200 34642 40000 34672
rect 38009 34640 40000 34642
rect 38009 34584 38014 34640
rect 38070 34584 40000 34640
rect 38009 34582 40000 34584
rect 38009 34579 38075 34582
rect 39200 34552 40000 34582
rect 0 34506 800 34536
rect 1393 34506 1459 34509
rect 0 34504 1459 34506
rect 0 34448 1398 34504
rect 1454 34448 1459 34504
rect 0 34446 1459 34448
rect 0 34416 800 34446
rect 1393 34443 1459 34446
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33872 800 33992
rect 38101 33962 38167 33965
rect 39200 33962 40000 33992
rect 38101 33960 40000 33962
rect 38101 33904 38106 33960
rect 38162 33904 40000 33960
rect 38101 33902 40000 33904
rect 38101 33899 38167 33902
rect 39200 33872 40000 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33554 800 33584
rect 1393 33554 1459 33557
rect 0 33552 1459 33554
rect 0 33496 1398 33552
rect 1454 33496 1459 33552
rect 0 33494 1459 33496
rect 0 33464 800 33494
rect 1393 33491 1459 33494
rect 38009 33282 38075 33285
rect 39200 33282 40000 33312
rect 38009 33280 40000 33282
rect 38009 33224 38014 33280
rect 38070 33224 40000 33280
rect 38009 33222 40000 33224
rect 38009 33219 38075 33222
rect 4208 33216 4528 33217
rect 0 33056 800 33176
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 39200 33192 40000 33222
rect 34928 33151 35248 33152
rect 0 32738 800 32768
rect 1393 32738 1459 32741
rect 0 32736 1459 32738
rect 0 32680 1398 32736
rect 1454 32680 1459 32736
rect 0 32678 1459 32680
rect 0 32648 800 32678
rect 1393 32675 1459 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 38009 32602 38075 32605
rect 39200 32602 40000 32632
rect 38009 32600 40000 32602
rect 38009 32544 38014 32600
rect 38070 32544 40000 32600
rect 38009 32542 40000 32544
rect 38009 32539 38075 32542
rect 39200 32512 40000 32542
rect 0 32104 800 32224
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 38101 31922 38167 31925
rect 39200 31922 40000 31952
rect 38101 31920 40000 31922
rect 38101 31864 38106 31920
rect 38162 31864 40000 31920
rect 38101 31862 40000 31864
rect 38101 31859 38167 31862
rect 39200 31832 40000 31862
rect 0 31786 800 31816
rect 1485 31786 1551 31789
rect 0 31784 1551 31786
rect 0 31728 1490 31784
rect 1546 31728 1551 31784
rect 0 31726 1551 31728
rect 0 31696 800 31726
rect 1485 31723 1551 31726
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 38009 31106 38075 31109
rect 39200 31106 40000 31136
rect 38009 31104 40000 31106
rect 38009 31048 38014 31104
rect 38070 31048 40000 31104
rect 38009 31046 40000 31048
rect 38009 31043 38075 31046
rect 4208 31040 4528 31041
rect 0 30880 800 31000
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 39200 31016 40000 31046
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 0 30426 800 30456
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 1393 30426 1459 30429
rect 0 30424 1459 30426
rect 0 30368 1398 30424
rect 1454 30368 1459 30424
rect 0 30366 1459 30368
rect 0 30336 800 30366
rect 1393 30363 1459 30366
rect 38009 30426 38075 30429
rect 39200 30426 40000 30456
rect 38009 30424 40000 30426
rect 38009 30368 38014 30424
rect 38070 30368 40000 30424
rect 38009 30366 40000 30368
rect 38009 30363 38075 30366
rect 39200 30336 40000 30366
rect 0 30018 800 30048
rect 1393 30018 1459 30021
rect 0 30016 1459 30018
rect 0 29960 1398 30016
rect 1454 29960 1459 30016
rect 0 29958 1459 29960
rect 0 29928 800 29958
rect 1393 29955 1459 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 38101 29746 38167 29749
rect 39200 29746 40000 29776
rect 38101 29744 40000 29746
rect 38101 29688 38106 29744
rect 38162 29688 40000 29744
rect 38101 29686 40000 29688
rect 38101 29683 38167 29686
rect 39200 29656 40000 29686
rect 0 29520 800 29640
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 0 29202 800 29232
rect 1393 29202 1459 29205
rect 0 29200 1459 29202
rect 0 29144 1398 29200
rect 1454 29144 1459 29200
rect 0 29142 1459 29144
rect 0 29112 800 29142
rect 1393 29139 1459 29142
rect 38009 29066 38075 29069
rect 39200 29066 40000 29096
rect 38009 29064 40000 29066
rect 38009 29008 38014 29064
rect 38070 29008 40000 29064
rect 38009 29006 40000 29008
rect 38009 29003 38075 29006
rect 39200 28976 40000 29006
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 1393 28794 1459 28797
rect 0 28792 1459 28794
rect 0 28736 1398 28792
rect 1454 28736 1459 28792
rect 0 28734 1459 28736
rect 0 28704 800 28734
rect 1393 28731 1459 28734
rect 38009 28386 38075 28389
rect 39200 28386 40000 28416
rect 38009 28384 40000 28386
rect 38009 28328 38014 28384
rect 38070 28328 40000 28384
rect 38009 28326 40000 28328
rect 38009 28323 38075 28326
rect 19568 28320 19888 28321
rect 0 28160 800 28280
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 39200 28296 40000 28326
rect 19568 28255 19888 28256
rect 0 27842 800 27872
rect 1393 27842 1459 27845
rect 0 27840 1459 27842
rect 0 27784 1398 27840
rect 1454 27784 1459 27840
rect 0 27782 1459 27784
rect 0 27752 800 27782
rect 1393 27779 1459 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 38101 27706 38167 27709
rect 39200 27706 40000 27736
rect 38101 27704 40000 27706
rect 38101 27648 38106 27704
rect 38162 27648 40000 27704
rect 38101 27646 40000 27648
rect 38101 27643 38167 27646
rect 39200 27616 40000 27646
rect 0 27434 800 27464
rect 1393 27434 1459 27437
rect 0 27432 1459 27434
rect 0 27376 1398 27432
rect 1454 27376 1459 27432
rect 0 27374 1459 27376
rect 0 27344 800 27374
rect 1393 27371 1459 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 0 26936 800 27056
rect 38009 27026 38075 27029
rect 39200 27026 40000 27056
rect 38009 27024 40000 27026
rect 38009 26968 38014 27024
rect 38070 26968 40000 27024
rect 38009 26966 40000 26968
rect 38009 26963 38075 26966
rect 39200 26936 40000 26966
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 0 26482 800 26512
rect 1393 26482 1459 26485
rect 0 26480 1459 26482
rect 0 26424 1398 26480
rect 1454 26424 1459 26480
rect 0 26422 1459 26424
rect 0 26392 800 26422
rect 1393 26419 1459 26422
rect 37365 26482 37431 26485
rect 38101 26482 38167 26485
rect 37365 26480 38167 26482
rect 37365 26424 37370 26480
rect 37426 26424 38106 26480
rect 38162 26424 38167 26480
rect 37365 26422 38167 26424
rect 37365 26419 37431 26422
rect 38101 26419 38167 26422
rect 38009 26210 38075 26213
rect 39200 26210 40000 26240
rect 38009 26208 40000 26210
rect 38009 26152 38014 26208
rect 38070 26152 40000 26208
rect 38009 26150 40000 26152
rect 38009 26147 38075 26150
rect 19568 26144 19888 26145
rect 0 26074 800 26104
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 39200 26120 40000 26150
rect 19568 26079 19888 26080
rect 1485 26074 1551 26077
rect 0 26072 1551 26074
rect 0 26016 1490 26072
rect 1546 26016 1551 26072
rect 0 26014 1551 26016
rect 0 25984 800 26014
rect 1485 26011 1551 26014
rect 0 25666 800 25696
rect 1393 25666 1459 25669
rect 0 25664 1459 25666
rect 0 25608 1398 25664
rect 1454 25608 1459 25664
rect 0 25606 1459 25608
rect 0 25576 800 25606
rect 1393 25603 1459 25606
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 37181 25530 37247 25533
rect 39200 25530 40000 25560
rect 37181 25528 40000 25530
rect 37181 25472 37186 25528
rect 37242 25472 40000 25528
rect 37181 25470 40000 25472
rect 37181 25467 37247 25470
rect 39200 25440 40000 25470
rect 0 25258 800 25288
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25168 800 25198
rect 1393 25195 1459 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 38009 24850 38075 24853
rect 39200 24850 40000 24880
rect 38009 24848 40000 24850
rect 38009 24792 38014 24848
rect 38070 24792 40000 24848
rect 38009 24790 40000 24792
rect 38009 24787 38075 24790
rect 39200 24760 40000 24790
rect 0 24714 800 24744
rect 1485 24714 1551 24717
rect 0 24712 1551 24714
rect 0 24656 1490 24712
rect 1546 24656 1551 24712
rect 0 24654 1551 24656
rect 0 24624 800 24654
rect 1485 24651 1551 24654
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 0 24306 800 24336
rect 1853 24306 1919 24309
rect 0 24304 1919 24306
rect 0 24248 1858 24304
rect 1914 24248 1919 24304
rect 0 24246 1919 24248
rect 0 24216 800 24246
rect 1853 24243 1919 24246
rect 38009 24170 38075 24173
rect 39200 24170 40000 24200
rect 38009 24168 40000 24170
rect 38009 24112 38014 24168
rect 38070 24112 40000 24168
rect 38009 24110 40000 24112
rect 38009 24107 38075 24110
rect 39200 24080 40000 24110
rect 19568 23968 19888 23969
rect 0 23898 800 23928
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 2129 23898 2195 23901
rect 0 23896 2195 23898
rect 0 23840 2134 23896
rect 2190 23840 2195 23896
rect 0 23838 2195 23840
rect 0 23808 800 23838
rect 2129 23835 2195 23838
rect 0 23490 800 23520
rect 1485 23490 1551 23493
rect 0 23488 1551 23490
rect 0 23432 1490 23488
rect 1546 23432 1551 23488
rect 0 23430 1551 23432
rect 0 23400 800 23430
rect 1485 23427 1551 23430
rect 38101 23490 38167 23493
rect 39200 23490 40000 23520
rect 38101 23488 40000 23490
rect 38101 23432 38106 23488
rect 38162 23432 40000 23488
rect 38101 23430 40000 23432
rect 38101 23427 38167 23430
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 39200 23400 40000 23430
rect 34928 23359 35248 23360
rect 0 23082 800 23112
rect 1853 23082 1919 23085
rect 0 23080 1919 23082
rect 0 23024 1858 23080
rect 1914 23024 1919 23080
rect 0 23022 1919 23024
rect 0 22992 800 23022
rect 1853 23019 1919 23022
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 38009 22810 38075 22813
rect 39200 22810 40000 22840
rect 38009 22808 40000 22810
rect 38009 22752 38014 22808
rect 38070 22752 40000 22808
rect 38009 22750 40000 22752
rect 38009 22747 38075 22750
rect 39200 22720 40000 22750
rect 0 22538 800 22568
rect 2129 22538 2195 22541
rect 0 22536 2195 22538
rect 0 22480 2134 22536
rect 2190 22480 2195 22536
rect 0 22478 2195 22480
rect 0 22448 800 22478
rect 2129 22475 2195 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 22130 800 22160
rect 1485 22130 1551 22133
rect 0 22128 1551 22130
rect 0 22072 1490 22128
rect 1546 22072 1551 22128
rect 0 22070 1551 22072
rect 0 22040 800 22070
rect 1485 22067 1551 22070
rect 24761 21994 24827 21997
rect 27797 21994 27863 21997
rect 24761 21992 27863 21994
rect 24761 21936 24766 21992
rect 24822 21936 27802 21992
rect 27858 21936 27863 21992
rect 24761 21934 27863 21936
rect 24761 21931 24827 21934
rect 27797 21931 27863 21934
rect 38009 21994 38075 21997
rect 39200 21994 40000 22024
rect 38009 21992 40000 21994
rect 38009 21936 38014 21992
rect 38070 21936 40000 21992
rect 38009 21934 40000 21936
rect 38009 21931 38075 21934
rect 39200 21904 40000 21934
rect 19568 21792 19888 21793
rect 0 21722 800 21752
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 1853 21722 1919 21725
rect 0 21720 1919 21722
rect 0 21664 1858 21720
rect 1914 21664 1919 21720
rect 0 21662 1919 21664
rect 0 21632 800 21662
rect 1853 21659 1919 21662
rect 0 21314 800 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 800 21254
rect 1393 21251 1459 21254
rect 36721 21314 36787 21317
rect 38101 21314 38167 21317
rect 39200 21314 40000 21344
rect 36721 21312 40000 21314
rect 36721 21256 36726 21312
rect 36782 21256 38106 21312
rect 38162 21256 40000 21312
rect 36721 21254 40000 21256
rect 36721 21251 36787 21254
rect 38101 21251 38167 21254
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 39200 21224 40000 21254
rect 34928 21183 35248 21184
rect 0 20770 800 20800
rect 1485 20770 1551 20773
rect 0 20768 1551 20770
rect 0 20712 1490 20768
rect 1546 20712 1551 20768
rect 0 20710 1551 20712
rect 0 20680 800 20710
rect 1485 20707 1551 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 36169 20634 36235 20637
rect 39200 20634 40000 20664
rect 36169 20632 40000 20634
rect 36169 20576 36174 20632
rect 36230 20576 40000 20632
rect 36169 20574 40000 20576
rect 36169 20571 36235 20574
rect 39200 20544 40000 20574
rect 0 20362 800 20392
rect 1853 20362 1919 20365
rect 0 20360 1919 20362
rect 0 20304 1858 20360
rect 1914 20304 1919 20360
rect 0 20302 1919 20304
rect 0 20272 800 20302
rect 1853 20299 1919 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19954 800 19984
rect 2773 19954 2839 19957
rect 0 19952 2839 19954
rect 0 19896 2778 19952
rect 2834 19896 2839 19952
rect 0 19894 2839 19896
rect 0 19864 800 19894
rect 2773 19891 2839 19894
rect 38009 19954 38075 19957
rect 39200 19954 40000 19984
rect 38009 19952 40000 19954
rect 38009 19896 38014 19952
rect 38070 19896 40000 19952
rect 38009 19894 40000 19896
rect 38009 19891 38075 19894
rect 39200 19864 40000 19894
rect 19568 19616 19888 19617
rect 0 19546 800 19576
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 1485 19546 1551 19549
rect 0 19544 1551 19546
rect 0 19488 1490 19544
rect 1546 19488 1551 19544
rect 0 19486 1551 19488
rect 0 19456 800 19486
rect 1485 19483 1551 19486
rect 13721 19274 13787 19277
rect 22921 19274 22987 19277
rect 13721 19272 22987 19274
rect 13721 19216 13726 19272
rect 13782 19216 22926 19272
rect 22982 19216 22987 19272
rect 13721 19214 22987 19216
rect 13721 19211 13787 19214
rect 22921 19211 22987 19214
rect 38101 19274 38167 19277
rect 39200 19274 40000 19304
rect 38101 19272 40000 19274
rect 38101 19216 38106 19272
rect 38162 19216 40000 19272
rect 38101 19214 40000 19216
rect 38101 19211 38167 19214
rect 39200 19184 40000 19214
rect 4208 19072 4528 19073
rect 0 19002 800 19032
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 1853 19002 1919 19005
rect 0 19000 1919 19002
rect 0 18944 1858 19000
rect 1914 18944 1919 19000
rect 0 18942 1919 18944
rect 0 18912 800 18942
rect 1853 18939 1919 18942
rect 19977 18866 20043 18869
rect 20161 18866 20227 18869
rect 19977 18864 20227 18866
rect 19977 18808 19982 18864
rect 20038 18808 20166 18864
rect 20222 18808 20227 18864
rect 19977 18806 20227 18808
rect 19977 18803 20043 18806
rect 20161 18803 20227 18806
rect 19701 18730 19767 18733
rect 20345 18730 20411 18733
rect 21449 18730 21515 18733
rect 19701 18728 21515 18730
rect 19701 18672 19706 18728
rect 19762 18672 20350 18728
rect 20406 18672 21454 18728
rect 21510 18672 21515 18728
rect 19701 18670 21515 18672
rect 19701 18667 19767 18670
rect 20345 18667 20411 18670
rect 21449 18667 21515 18670
rect 0 18594 800 18624
rect 1393 18594 1459 18597
rect 0 18592 1459 18594
rect 0 18536 1398 18592
rect 1454 18536 1459 18592
rect 0 18534 1459 18536
rect 0 18504 800 18534
rect 1393 18531 1459 18534
rect 38009 18594 38075 18597
rect 39200 18594 40000 18624
rect 38009 18592 40000 18594
rect 38009 18536 38014 18592
rect 38070 18536 40000 18592
rect 38009 18534 40000 18536
rect 38009 18531 38075 18534
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 39200 18504 40000 18534
rect 19568 18463 19888 18464
rect 0 18186 800 18216
rect 1485 18186 1551 18189
rect 0 18184 1551 18186
rect 0 18128 1490 18184
rect 1546 18128 1551 18184
rect 0 18126 1551 18128
rect 0 18096 800 18126
rect 1485 18123 1551 18126
rect 19609 18186 19675 18189
rect 21357 18186 21423 18189
rect 19609 18184 21423 18186
rect 19609 18128 19614 18184
rect 19670 18128 21362 18184
rect 21418 18128 21423 18184
rect 19609 18126 21423 18128
rect 19609 18123 19675 18126
rect 21357 18123 21423 18126
rect 19333 18050 19399 18053
rect 20621 18050 20687 18053
rect 19333 18048 20687 18050
rect 19333 17992 19338 18048
rect 19394 17992 20626 18048
rect 20682 17992 20687 18048
rect 19333 17990 20687 17992
rect 19333 17987 19399 17990
rect 20621 17987 20687 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 1853 17778 1919 17781
rect 0 17776 1919 17778
rect 0 17720 1858 17776
rect 1914 17720 1919 17776
rect 0 17718 1919 17720
rect 0 17688 800 17718
rect 1853 17715 1919 17718
rect 6269 17778 6335 17781
rect 14181 17778 14247 17781
rect 6269 17776 14247 17778
rect 6269 17720 6274 17776
rect 6330 17720 14186 17776
rect 14242 17720 14247 17776
rect 6269 17718 14247 17720
rect 6269 17715 6335 17718
rect 14181 17715 14247 17718
rect 38009 17778 38075 17781
rect 39200 17778 40000 17808
rect 38009 17776 40000 17778
rect 38009 17720 38014 17776
rect 38070 17720 40000 17776
rect 38009 17718 40000 17720
rect 38009 17715 38075 17718
rect 39200 17688 40000 17718
rect 7557 17642 7623 17645
rect 35341 17642 35407 17645
rect 7557 17640 35407 17642
rect 7557 17584 7562 17640
rect 7618 17584 35346 17640
rect 35402 17584 35407 17640
rect 7557 17582 35407 17584
rect 7557 17579 7623 17582
rect 35341 17579 35407 17582
rect 11145 17506 11211 17509
rect 13353 17506 13419 17509
rect 11145 17504 13419 17506
rect 11145 17448 11150 17504
rect 11206 17448 13358 17504
rect 13414 17448 13419 17504
rect 11145 17446 13419 17448
rect 11145 17443 11211 17446
rect 13353 17443 13419 17446
rect 19568 17440 19888 17441
rect 0 17370 800 17400
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 2129 17370 2195 17373
rect 0 17368 2195 17370
rect 0 17312 2134 17368
rect 2190 17312 2195 17368
rect 0 17310 2195 17312
rect 0 17280 800 17310
rect 2129 17307 2195 17310
rect 19057 17234 19123 17237
rect 19241 17234 19307 17237
rect 19057 17232 19307 17234
rect 19057 17176 19062 17232
rect 19118 17176 19246 17232
rect 19302 17176 19307 17232
rect 19057 17174 19307 17176
rect 19057 17171 19123 17174
rect 19241 17171 19307 17174
rect 7741 17098 7807 17101
rect 31845 17098 31911 17101
rect 7741 17096 31911 17098
rect 7741 17040 7746 17096
rect 7802 17040 31850 17096
rect 31906 17040 31911 17096
rect 7741 17038 31911 17040
rect 7741 17035 7807 17038
rect 31845 17035 31911 17038
rect 38101 17098 38167 17101
rect 39200 17098 40000 17128
rect 38101 17096 40000 17098
rect 38101 17040 38106 17096
rect 38162 17040 40000 17096
rect 38101 17038 40000 17040
rect 38101 17035 38167 17038
rect 39200 17008 40000 17038
rect 4208 16896 4528 16897
rect 0 16826 800 16856
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 7005 16554 7071 16557
rect 27613 16554 27679 16557
rect 7005 16552 27679 16554
rect 7005 16496 7010 16552
rect 7066 16496 27618 16552
rect 27674 16496 27679 16552
rect 7005 16494 27679 16496
rect 7005 16491 7071 16494
rect 27613 16491 27679 16494
rect 0 16418 800 16448
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16328 800 16358
rect 1853 16355 1919 16358
rect 36169 16418 36235 16421
rect 39200 16418 40000 16448
rect 36169 16416 40000 16418
rect 36169 16360 36174 16416
rect 36230 16360 40000 16416
rect 36169 16358 40000 16360
rect 36169 16355 36235 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 39200 16328 40000 16358
rect 19568 16287 19888 16288
rect 1669 16146 1735 16149
rect 18505 16146 18571 16149
rect 1669 16144 18571 16146
rect 1669 16088 1674 16144
rect 1730 16088 18510 16144
rect 18566 16088 18571 16144
rect 1669 16086 18571 16088
rect 1669 16083 1735 16086
rect 18505 16083 18571 16086
rect 22461 16146 22527 16149
rect 22829 16146 22895 16149
rect 22461 16144 22895 16146
rect 22461 16088 22466 16144
rect 22522 16088 22834 16144
rect 22890 16088 22895 16144
rect 22461 16086 22895 16088
rect 22461 16083 22527 16086
rect 22829 16083 22895 16086
rect 0 16010 800 16040
rect 2129 16010 2195 16013
rect 0 16008 2195 16010
rect 0 15952 2134 16008
rect 2190 15952 2195 16008
rect 0 15950 2195 15952
rect 0 15920 800 15950
rect 2129 15947 2195 15950
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 38009 15738 38075 15741
rect 39200 15738 40000 15768
rect 38009 15736 40000 15738
rect 38009 15680 38014 15736
rect 38070 15680 40000 15736
rect 38009 15678 40000 15680
rect 38009 15675 38075 15678
rect 39200 15648 40000 15678
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 12801 15602 12867 15605
rect 35709 15602 35775 15605
rect 12801 15600 35775 15602
rect 12801 15544 12806 15600
rect 12862 15544 35714 15600
rect 35770 15544 35775 15600
rect 12801 15542 35775 15544
rect 12801 15539 12867 15542
rect 35709 15539 35775 15542
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15088
rect 1853 15058 1919 15061
rect 0 15056 1919 15058
rect 0 15000 1858 15056
rect 1914 15000 1919 15056
rect 0 14998 1919 15000
rect 0 14968 800 14998
rect 1853 14995 1919 14998
rect 17309 15058 17375 15061
rect 18597 15058 18663 15061
rect 17309 15056 18663 15058
rect 17309 15000 17314 15056
rect 17370 15000 18602 15056
rect 18658 15000 18663 15056
rect 17309 14998 18663 15000
rect 17309 14995 17375 14998
rect 18597 14995 18663 14998
rect 38101 15058 38167 15061
rect 39200 15058 40000 15088
rect 38101 15056 40000 15058
rect 38101 15000 38106 15056
rect 38162 15000 40000 15056
rect 38101 14998 40000 15000
rect 38101 14995 38167 14998
rect 39200 14968 40000 14998
rect 18045 14922 18111 14925
rect 18781 14922 18847 14925
rect 18045 14920 18847 14922
rect 18045 14864 18050 14920
rect 18106 14864 18786 14920
rect 18842 14864 18847 14920
rect 18045 14862 18847 14864
rect 18045 14859 18111 14862
rect 18781 14859 18847 14862
rect 17401 14786 17467 14789
rect 17953 14786 18019 14789
rect 18965 14786 19031 14789
rect 17401 14784 19031 14786
rect 17401 14728 17406 14784
rect 17462 14728 17958 14784
rect 18014 14728 18970 14784
rect 19026 14728 19031 14784
rect 17401 14726 19031 14728
rect 17401 14723 17467 14726
rect 17953 14723 18019 14726
rect 18965 14723 19031 14726
rect 4208 14720 4528 14721
rect 0 14650 800 14680
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 1393 14650 1459 14653
rect 0 14648 1459 14650
rect 0 14592 1398 14648
rect 1454 14592 1459 14648
rect 0 14590 1459 14592
rect 0 14560 800 14590
rect 1393 14587 1459 14590
rect 1669 14514 1735 14517
rect 17769 14514 17835 14517
rect 1669 14512 17835 14514
rect 1669 14456 1674 14512
rect 1730 14456 17774 14512
rect 17830 14456 17835 14512
rect 1669 14454 17835 14456
rect 1669 14451 1735 14454
rect 17769 14451 17835 14454
rect 14825 14378 14891 14381
rect 17769 14378 17835 14381
rect 14825 14376 17835 14378
rect 14825 14320 14830 14376
rect 14886 14320 17774 14376
rect 17830 14320 17835 14376
rect 14825 14318 17835 14320
rect 14825 14315 14891 14318
rect 17769 14315 17835 14318
rect 36169 14378 36235 14381
rect 39200 14378 40000 14408
rect 36169 14376 40000 14378
rect 36169 14320 36174 14376
rect 36230 14320 40000 14376
rect 36169 14318 40000 14320
rect 36169 14315 36235 14318
rect 39200 14288 40000 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 13353 13970 13419 13973
rect 18505 13970 18571 13973
rect 13353 13968 18571 13970
rect 13353 13912 13358 13968
rect 13414 13912 18510 13968
rect 18566 13912 18571 13968
rect 13353 13910 18571 13912
rect 13353 13907 13419 13910
rect 18505 13907 18571 13910
rect 0 13834 800 13864
rect 1393 13834 1459 13837
rect 0 13832 1459 13834
rect 0 13776 1398 13832
rect 1454 13776 1459 13832
rect 0 13774 1459 13776
rect 0 13744 800 13774
rect 1393 13771 1459 13774
rect 17861 13834 17927 13837
rect 28993 13834 29059 13837
rect 17861 13832 29059 13834
rect 17861 13776 17866 13832
rect 17922 13776 28998 13832
rect 29054 13776 29059 13832
rect 17861 13774 29059 13776
rect 17861 13771 17927 13774
rect 28993 13771 29059 13774
rect 38009 13698 38075 13701
rect 39200 13698 40000 13728
rect 38009 13696 40000 13698
rect 38009 13640 38014 13696
rect 38070 13640 40000 13696
rect 38009 13638 40000 13640
rect 38009 13635 38075 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 39200 13608 40000 13638
rect 34928 13567 35248 13568
rect 1669 13426 1735 13429
rect 17033 13426 17099 13429
rect 1669 13424 17099 13426
rect 1669 13368 1674 13424
rect 1730 13368 17038 13424
rect 17094 13368 17099 13424
rect 1669 13366 17099 13368
rect 1669 13363 1735 13366
rect 17033 13363 17099 13366
rect 0 13290 800 13320
rect 2129 13290 2195 13293
rect 0 13288 2195 13290
rect 0 13232 2134 13288
rect 2190 13232 2195 13288
rect 0 13230 2195 13232
rect 0 13200 800 13230
rect 2129 13227 2195 13230
rect 10685 13290 10751 13293
rect 15469 13290 15535 13293
rect 10685 13288 15535 13290
rect 10685 13232 10690 13288
rect 10746 13232 15474 13288
rect 15530 13232 15535 13288
rect 10685 13230 15535 13232
rect 10685 13227 10751 13230
rect 15469 13227 15535 13230
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 0 12882 800 12912
rect 1485 12882 1551 12885
rect 0 12880 1551 12882
rect 0 12824 1490 12880
rect 1546 12824 1551 12880
rect 0 12822 1551 12824
rect 0 12792 800 12822
rect 1485 12819 1551 12822
rect 38101 12882 38167 12885
rect 39200 12882 40000 12912
rect 38101 12880 40000 12882
rect 38101 12824 38106 12880
rect 38162 12824 40000 12880
rect 38101 12822 40000 12824
rect 38101 12819 38167 12822
rect 39200 12792 40000 12822
rect 17861 12746 17927 12749
rect 36813 12746 36879 12749
rect 17861 12744 36879 12746
rect 17861 12688 17866 12744
rect 17922 12688 36818 12744
rect 36874 12688 36879 12744
rect 17861 12686 36879 12688
rect 17861 12683 17927 12686
rect 36813 12683 36879 12686
rect 4208 12544 4528 12545
rect 0 12474 800 12504
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 1853 12474 1919 12477
rect 0 12472 1919 12474
rect 0 12416 1858 12472
rect 1914 12416 1919 12472
rect 0 12414 1919 12416
rect 0 12384 800 12414
rect 1853 12411 1919 12414
rect 38009 12202 38075 12205
rect 39200 12202 40000 12232
rect 38009 12200 40000 12202
rect 38009 12144 38014 12200
rect 38070 12144 40000 12200
rect 38009 12142 40000 12144
rect 38009 12139 38075 12142
rect 39200 12112 40000 12142
rect 0 12066 800 12096
rect 1393 12066 1459 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 800 12006
rect 1393 12003 1459 12006
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 38009 11522 38075 11525
rect 39200 11522 40000 11552
rect 38009 11520 40000 11522
rect 38009 11464 38014 11520
rect 38070 11464 40000 11520
rect 38009 11462 40000 11464
rect 38009 11459 38075 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 39200 11432 40000 11462
rect 34928 11391 35248 11392
rect 0 11114 800 11144
rect 1853 11114 1919 11117
rect 0 11112 1919 11114
rect 0 11056 1858 11112
rect 1914 11056 1919 11112
rect 0 11054 1919 11056
rect 0 11024 800 11054
rect 1853 11051 1919 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 36445 10842 36511 10845
rect 39200 10842 40000 10872
rect 36445 10840 40000 10842
rect 36445 10784 36450 10840
rect 36506 10784 40000 10840
rect 36445 10782 40000 10784
rect 36445 10779 36511 10782
rect 39200 10752 40000 10782
rect 0 10706 800 10736
rect 2865 10706 2931 10709
rect 0 10704 2931 10706
rect 0 10648 2870 10704
rect 2926 10648 2931 10704
rect 0 10646 2931 10648
rect 0 10616 800 10646
rect 2865 10643 2931 10646
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 37181 10162 37247 10165
rect 39200 10162 40000 10192
rect 37181 10160 40000 10162
rect 37181 10104 37186 10160
rect 37242 10104 40000 10160
rect 37181 10102 40000 10104
rect 37181 10099 37247 10102
rect 39200 10072 40000 10102
rect 0 9890 800 9920
rect 1853 9890 1919 9893
rect 0 9888 1919 9890
rect 0 9832 1858 9888
rect 1914 9832 1919 9888
rect 0 9830 1919 9832
rect 0 9800 800 9830
rect 1853 9827 1919 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 38009 9482 38075 9485
rect 39200 9482 40000 9512
rect 38009 9480 40000 9482
rect 38009 9424 38014 9480
rect 38070 9424 40000 9480
rect 38009 9422 40000 9424
rect 38009 9419 38075 9422
rect 39200 9392 40000 9422
rect 0 9346 800 9376
rect 2037 9346 2103 9349
rect 0 9344 2103 9346
rect 0 9288 2042 9344
rect 2098 9288 2103 9344
rect 0 9286 2103 9288
rect 0 9256 800 9286
rect 2037 9283 2103 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 2773 8938 2839 8941
rect 2957 8938 3023 8941
rect 2773 8936 3023 8938
rect 2773 8880 2778 8936
rect 2834 8880 2962 8936
rect 3018 8880 3023 8936
rect 2773 8878 3023 8880
rect 2773 8875 2839 8878
rect 2957 8875 3023 8878
rect 11973 8938 12039 8941
rect 13353 8938 13419 8941
rect 11973 8936 13419 8938
rect 11973 8880 11978 8936
rect 12034 8880 13358 8936
rect 13414 8880 13419 8936
rect 11973 8878 13419 8880
rect 11973 8875 12039 8878
rect 13353 8875 13419 8878
rect 12065 8802 12131 8805
rect 17217 8802 17283 8805
rect 12065 8800 17283 8802
rect 12065 8744 12070 8800
rect 12126 8744 17222 8800
rect 17278 8744 17283 8800
rect 12065 8742 17283 8744
rect 12065 8739 12131 8742
rect 17217 8739 17283 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 38101 8666 38167 8669
rect 39200 8666 40000 8696
rect 38101 8664 40000 8666
rect 38101 8608 38106 8664
rect 38162 8608 40000 8664
rect 38101 8606 40000 8608
rect 38101 8603 38167 8606
rect 39200 8576 40000 8606
rect 0 8530 800 8560
rect 2773 8530 2839 8533
rect 0 8528 2839 8530
rect 0 8472 2778 8528
rect 2834 8472 2839 8528
rect 0 8470 2839 8472
rect 0 8440 800 8470
rect 2773 8467 2839 8470
rect 4208 8192 4528 8193
rect 0 8122 800 8152
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 38009 7986 38075 7989
rect 39200 7986 40000 8016
rect 38009 7984 40000 7986
rect 38009 7928 38014 7984
rect 38070 7928 40000 7984
rect 38009 7926 40000 7928
rect 38009 7923 38075 7926
rect 39200 7896 40000 7926
rect 19568 7648 19888 7649
rect 0 7578 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 12801 7306 12867 7309
rect 37365 7306 37431 7309
rect 12801 7304 37431 7306
rect 12801 7248 12806 7304
rect 12862 7248 37370 7304
rect 37426 7248 37431 7304
rect 12801 7246 37431 7248
rect 12801 7243 12867 7246
rect 37365 7243 37431 7246
rect 38009 7306 38075 7309
rect 39200 7306 40000 7336
rect 38009 7304 40000 7306
rect 38009 7248 38014 7304
rect 38070 7248 40000 7304
rect 38009 7246 40000 7248
rect 38009 7243 38075 7246
rect 39200 7216 40000 7246
rect 0 7170 800 7200
rect 1393 7170 1459 7173
rect 0 7168 1459 7170
rect 0 7112 1398 7168
rect 1454 7112 1459 7168
rect 0 7110 1459 7112
rect 0 7080 800 7110
rect 1393 7107 1459 7110
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6762 800 6792
rect 2037 6762 2103 6765
rect 0 6760 2103 6762
rect 0 6704 2042 6760
rect 2098 6704 2103 6760
rect 0 6702 2103 6704
rect 0 6672 800 6702
rect 2037 6699 2103 6702
rect 16297 6762 16363 6765
rect 17493 6762 17559 6765
rect 17953 6762 18019 6765
rect 16297 6760 18019 6762
rect 16297 6704 16302 6760
rect 16358 6704 17498 6760
rect 17554 6704 17958 6760
rect 18014 6704 18019 6760
rect 16297 6702 18019 6704
rect 16297 6699 16363 6702
rect 17493 6699 17559 6702
rect 17953 6699 18019 6702
rect 14457 6626 14523 6629
rect 17769 6626 17835 6629
rect 14457 6624 17835 6626
rect 14457 6568 14462 6624
rect 14518 6568 17774 6624
rect 17830 6568 17835 6624
rect 14457 6566 17835 6568
rect 14457 6563 14523 6566
rect 17769 6563 17835 6566
rect 36445 6626 36511 6629
rect 39200 6626 40000 6656
rect 36445 6624 40000 6626
rect 36445 6568 36450 6624
rect 36506 6568 40000 6624
rect 36445 6566 40000 6568
rect 36445 6563 36511 6566
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 39200 6536 40000 6566
rect 19568 6495 19888 6496
rect 0 6354 800 6384
rect 1485 6354 1551 6357
rect 0 6352 1551 6354
rect 0 6296 1490 6352
rect 1546 6296 1551 6352
rect 0 6294 1551 6296
rect 0 6264 800 6294
rect 1485 6291 1551 6294
rect 4208 6016 4528 6017
rect 0 5946 800 5976
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 1853 5946 1919 5949
rect 0 5944 1919 5946
rect 0 5888 1858 5944
rect 1914 5888 1919 5944
rect 0 5886 1919 5888
rect 0 5856 800 5886
rect 1853 5883 1919 5886
rect 37273 5946 37339 5949
rect 39200 5946 40000 5976
rect 37273 5944 40000 5946
rect 37273 5888 37278 5944
rect 37334 5888 40000 5944
rect 37273 5886 40000 5888
rect 37273 5883 37339 5886
rect 39200 5856 40000 5886
rect 12249 5810 12315 5813
rect 26141 5810 26207 5813
rect 12249 5808 26207 5810
rect 12249 5752 12254 5808
rect 12310 5752 26146 5808
rect 26202 5752 26207 5808
rect 12249 5750 26207 5752
rect 12249 5747 12315 5750
rect 26141 5747 26207 5750
rect 1669 5674 1735 5677
rect 12893 5674 12959 5677
rect 1669 5672 12959 5674
rect 1669 5616 1674 5672
rect 1730 5616 12898 5672
rect 12954 5616 12959 5672
rect 1669 5614 12959 5616
rect 1669 5611 1735 5614
rect 12893 5611 12959 5614
rect 19568 5472 19888 5473
rect 0 5402 800 5432
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 2865 5402 2931 5405
rect 0 5400 2931 5402
rect 0 5344 2870 5400
rect 2926 5344 2931 5400
rect 0 5342 2931 5344
rect 0 5312 800 5342
rect 2865 5339 2931 5342
rect 12249 5266 12315 5269
rect 27429 5266 27495 5269
rect 12249 5264 27495 5266
rect 12249 5208 12254 5264
rect 12310 5208 27434 5264
rect 27490 5208 27495 5264
rect 12249 5206 27495 5208
rect 12249 5203 12315 5206
rect 27429 5203 27495 5206
rect 38009 5266 38075 5269
rect 39200 5266 40000 5296
rect 38009 5264 40000 5266
rect 38009 5208 38014 5264
rect 38070 5208 40000 5264
rect 38009 5206 40000 5208
rect 38009 5203 38075 5206
rect 39200 5176 40000 5206
rect 12709 5130 12775 5133
rect 37365 5130 37431 5133
rect 12709 5128 37431 5130
rect 12709 5072 12714 5128
rect 12770 5072 37370 5128
rect 37426 5072 37431 5128
rect 12709 5070 37431 5072
rect 12709 5067 12775 5070
rect 37365 5067 37431 5070
rect 0 4994 800 5024
rect 2957 4994 3023 4997
rect 0 4992 3023 4994
rect 0 4936 2962 4992
rect 3018 4936 3023 4992
rect 0 4934 3023 4936
rect 0 4904 800 4934
rect 2957 4931 3023 4934
rect 13169 4994 13235 4997
rect 26785 4994 26851 4997
rect 13169 4992 26851 4994
rect 13169 4936 13174 4992
rect 13230 4936 26790 4992
rect 26846 4936 26851 4992
rect 13169 4934 26851 4936
rect 13169 4931 13235 4934
rect 26785 4931 26851 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 16205 4858 16271 4861
rect 18597 4858 18663 4861
rect 16205 4856 18663 4858
rect 16205 4800 16210 4856
rect 16266 4800 18602 4856
rect 18658 4800 18663 4856
rect 16205 4798 18663 4800
rect 16205 4795 16271 4798
rect 18597 4795 18663 4798
rect 3233 4722 3299 4725
rect 4061 4722 4127 4725
rect 4245 4722 4311 4725
rect 29821 4722 29887 4725
rect 3233 4720 29887 4722
rect 3233 4664 3238 4720
rect 3294 4664 4066 4720
rect 4122 4664 4250 4720
rect 4306 4664 29826 4720
rect 29882 4664 29887 4720
rect 3233 4662 29887 4664
rect 3233 4659 3299 4662
rect 4061 4659 4127 4662
rect 4245 4659 4311 4662
rect 29821 4659 29887 4662
rect 0 4586 800 4616
rect 1853 4586 1919 4589
rect 0 4584 1919 4586
rect 0 4528 1858 4584
rect 1914 4528 1919 4584
rect 0 4526 1919 4528
rect 0 4496 800 4526
rect 1853 4523 1919 4526
rect 15193 4586 15259 4589
rect 16849 4586 16915 4589
rect 15193 4584 16915 4586
rect 15193 4528 15198 4584
rect 15254 4528 16854 4584
rect 16910 4528 16915 4584
rect 15193 4526 16915 4528
rect 15193 4523 15259 4526
rect 16849 4523 16915 4526
rect 35709 4450 35775 4453
rect 39200 4450 40000 4480
rect 35709 4448 40000 4450
rect 35709 4392 35714 4448
rect 35770 4392 40000 4448
rect 35709 4390 40000 4392
rect 35709 4387 35775 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 39200 4360 40000 4390
rect 19568 4319 19888 4320
rect 0 4178 800 4208
rect 1577 4178 1643 4181
rect 0 4176 1643 4178
rect 0 4120 1582 4176
rect 1638 4120 1643 4176
rect 0 4118 1643 4120
rect 0 4088 800 4118
rect 1577 4115 1643 4118
rect 13353 4042 13419 4045
rect 37365 4042 37431 4045
rect 13353 4040 37431 4042
rect 13353 3984 13358 4040
rect 13414 3984 37370 4040
rect 37426 3984 37431 4040
rect 13353 3982 37431 3984
rect 13353 3979 13419 3982
rect 37365 3979 37431 3982
rect 10317 3906 10383 3909
rect 17769 3906 17835 3909
rect 10317 3904 17835 3906
rect 10317 3848 10322 3904
rect 10378 3848 17774 3904
rect 17830 3848 17835 3904
rect 10317 3846 17835 3848
rect 10317 3843 10383 3846
rect 17769 3843 17835 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 12893 3770 12959 3773
rect 19057 3770 19123 3773
rect 12893 3768 19123 3770
rect 12893 3712 12898 3768
rect 12954 3712 19062 3768
rect 19118 3712 19123 3768
rect 12893 3710 19123 3712
rect 12893 3707 12959 3710
rect 19057 3707 19123 3710
rect 36629 3770 36695 3773
rect 39200 3770 40000 3800
rect 36629 3768 40000 3770
rect 36629 3712 36634 3768
rect 36690 3712 40000 3768
rect 36629 3710 40000 3712
rect 36629 3707 36695 3710
rect 39200 3680 40000 3710
rect 0 3634 800 3664
rect 2773 3634 2839 3637
rect 0 3632 2839 3634
rect 0 3576 2778 3632
rect 2834 3576 2839 3632
rect 0 3574 2839 3576
rect 0 3544 800 3574
rect 2773 3571 2839 3574
rect 10317 3498 10383 3501
rect 10961 3498 11027 3501
rect 11789 3498 11855 3501
rect 10317 3496 11855 3498
rect 10317 3440 10322 3496
rect 10378 3440 10966 3496
rect 11022 3440 11794 3496
rect 11850 3440 11855 3496
rect 10317 3438 11855 3440
rect 10317 3435 10383 3438
rect 10961 3435 11027 3438
rect 11789 3435 11855 3438
rect 9673 3362 9739 3365
rect 10777 3362 10843 3365
rect 9673 3360 10843 3362
rect 9673 3304 9678 3360
rect 9734 3304 10782 3360
rect 10838 3304 10843 3360
rect 9673 3302 10843 3304
rect 9673 3299 9739 3302
rect 10777 3299 10843 3302
rect 19568 3296 19888 3297
rect 0 3226 800 3256
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 1393 3226 1459 3229
rect 0 3224 1459 3226
rect 0 3168 1398 3224
rect 1454 3168 1459 3224
rect 0 3166 1459 3168
rect 0 3136 800 3166
rect 1393 3163 1459 3166
rect 37273 3090 37339 3093
rect 39200 3090 40000 3120
rect 37273 3088 40000 3090
rect 37273 3032 37278 3088
rect 37334 3032 40000 3088
rect 37273 3030 40000 3032
rect 37273 3027 37339 3030
rect 39200 3000 40000 3030
rect 0 2818 800 2848
rect 3509 2818 3575 2821
rect 0 2816 3575 2818
rect 0 2760 3514 2816
rect 3570 2760 3575 2816
rect 0 2758 3575 2760
rect 0 2728 800 2758
rect 3509 2755 3575 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 0 2410 800 2440
rect 1485 2410 1551 2413
rect 0 2408 1551 2410
rect 0 2352 1490 2408
rect 1546 2352 1551 2408
rect 0 2350 1551 2352
rect 0 2320 800 2350
rect 1485 2347 1551 2350
rect 38101 2410 38167 2413
rect 39200 2410 40000 2440
rect 38101 2408 40000 2410
rect 38101 2352 38106 2408
rect 38162 2352 40000 2408
rect 38101 2350 40000 2352
rect 38101 2347 38167 2350
rect 39200 2320 40000 2350
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 0 1866 800 1896
rect 2865 1866 2931 1869
rect 0 1864 2931 1866
rect 0 1808 2870 1864
rect 2926 1808 2931 1864
rect 0 1806 2931 1808
rect 0 1776 800 1806
rect 2865 1803 2931 1806
rect 36629 1730 36695 1733
rect 39200 1730 40000 1760
rect 36629 1728 40000 1730
rect 36629 1672 36634 1728
rect 36690 1672 40000 1728
rect 36629 1670 40000 1672
rect 36629 1667 36695 1670
rect 39200 1640 40000 1670
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 0 1050 800 1080
rect 3325 1050 3391 1053
rect 0 1048 3391 1050
rect 0 992 3330 1048
rect 3386 992 3391 1048
rect 0 990 3391 992
rect 0 960 800 990
rect 3325 987 3391 990
rect 38009 1050 38075 1053
rect 39200 1050 40000 1080
rect 38009 1048 40000 1050
rect 38009 992 38014 1048
rect 38070 992 40000 1048
rect 38009 990 40000 992
rect 38009 987 38075 990
rect 39200 960 40000 990
rect 0 642 800 672
rect 3969 642 4035 645
rect 0 640 4035 642
rect 0 584 3974 640
rect 4030 584 4035 640
rect 0 582 4035 584
rect 0 552 800 582
rect 3969 579 4035 582
rect 37365 370 37431 373
rect 39200 370 40000 400
rect 37365 368 40000 370
rect 37365 312 37370 368
rect 37426 312 40000 368
rect 37365 310 40000 312
rect 37365 307 37431 310
rect 39200 280 40000 310
rect 0 234 800 264
rect 3969 234 4035 237
rect 0 232 4035 234
rect 0 176 3974 232
rect 4030 176 4035 232
rect 0 174 4035 176
rect 0 144 800 174
rect 3969 171 4035 174
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__A PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10856 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__B
timestamp 1644511149
transform 1 0 4416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__A_N
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__C
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__A
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__A
timestamp 1644511149
transform -1 0 20056 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__A
timestamp 1644511149
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__A
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__B
timestamp 1644511149
transform 1 0 6256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1644511149
transform -1 0 36340 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__A
timestamp 1644511149
transform 1 0 34776 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1644511149
transform 1 0 35696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__A
timestamp 1644511149
transform -1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__B
timestamp 1644511149
transform -1 0 26404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A2
timestamp 1644511149
transform -1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__B1
timestamp 1644511149
transform -1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__C1
timestamp 1644511149
transform -1 0 10948 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__A
timestamp 1644511149
transform 1 0 19596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__C
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A2
timestamp 1644511149
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A3
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A2
timestamp 1644511149
transform -1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A1
timestamp 1644511149
transform -1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__A
timestamp 1644511149
transform 1 0 25668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__A
timestamp 1644511149
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__A
timestamp 1644511149
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A2
timestamp 1644511149
transform -1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A2
timestamp 1644511149
transform -1 0 13248 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A2
timestamp 1644511149
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A2
timestamp 1644511149
transform -1 0 13064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1644511149
transform -1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1644511149
transform -1 0 35512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A
timestamp 1644511149
transform -1 0 35880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A2
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A
timestamp 1644511149
transform -1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1644511149
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A2
timestamp 1644511149
transform -1 0 17940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1644511149
transform -1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A2
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1644511149
transform -1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A2
timestamp 1644511149
transform -1 0 17940 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A2
timestamp 1644511149
transform -1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 1644511149
transform -1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1644511149
transform 1 0 35328 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A
timestamp 1644511149
transform -1 0 34960 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A2
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A
timestamp 1644511149
transform 1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A
timestamp 1644511149
transform -1 0 21252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1644511149
transform -1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1644511149
transform -1 0 25300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1644511149
transform -1 0 25300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1644511149
transform 1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A2
timestamp 1644511149
transform -1 0 37536 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__C1
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1644511149
transform 1 0 24472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1644511149
transform 1 0 23736 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A2
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A2
timestamp 1644511149
transform 1 0 36156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__C1
timestamp 1644511149
transform -1 0 36708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__B
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A2
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A3
timestamp 1644511149
transform 1 0 22264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1644511149
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B
timestamp 1644511149
transform -1 0 23460 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A3
timestamp 1644511149
transform -1 0 22816 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp 1644511149
transform -1 0 35696 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__C1
timestamp 1644511149
transform -1 0 35144 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1644511149
transform -1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1644511149
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A2
timestamp 1644511149
transform -1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A3
timestamp 1644511149
transform -1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A1
timestamp 1644511149
transform 1 0 24104 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B
timestamp 1644511149
transform -1 0 23368 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A3
timestamp 1644511149
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__B1
timestamp 1644511149
transform -1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A2
timestamp 1644511149
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__C1
timestamp 1644511149
transform 1 0 36708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1644511149
transform -1 0 24748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A2
timestamp 1644511149
transform 1 0 25208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A3
timestamp 1644511149
transform -1 0 25944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A3
timestamp 1644511149
transform -1 0 22632 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B1
timestamp 1644511149
transform -1 0 22816 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1644511149
transform 1 0 32200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1644511149
transform 1 0 31832 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1644511149
transform -1 0 33212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A0
timestamp 1644511149
transform 1 0 34040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A0
timestamp 1644511149
transform 1 0 33396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A0
timestamp 1644511149
transform 1 0 34500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A0
timestamp 1644511149
transform 1 0 33580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A0
timestamp 1644511149
transform 1 0 34040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1644511149
transform 1 0 32936 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A0
timestamp 1644511149
transform 1 0 33488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A0
timestamp 1644511149
transform -1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A0
timestamp 1644511149
transform 1 0 33120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A0
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A0
timestamp 1644511149
transform 1 0 33396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1644511149
transform -1 0 32476 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A0
timestamp 1644511149
transform -1 0 31556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A0
timestamp 1644511149
transform -1 0 33488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A0
timestamp 1644511149
transform 1 0 34040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A0
timestamp 1644511149
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A0
timestamp 1644511149
transform 1 0 34040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A0
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__S
timestamp 1644511149
transform 1 0 33304 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A_N
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A0
timestamp 1644511149
transform -1 0 32936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__S
timestamp 1644511149
transform 1 0 33304 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A_N
timestamp 1644511149
transform -1 0 29992 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A0
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__S
timestamp 1644511149
transform 1 0 32384 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A_N
timestamp 1644511149
transform 1 0 30452 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A0
timestamp 1644511149
transform -1 0 34040 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S
timestamp 1644511149
transform -1 0 34868 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A_N
timestamp 1644511149
transform -1 0 33672 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1644511149
transform -1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A0
timestamp 1644511149
transform 1 0 30176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A_N
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1644511149
transform 1 0 28520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A
timestamp 1644511149
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A0
timestamp 1644511149
transform 1 0 27784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A0
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A0
timestamp 1644511149
transform 1 0 29256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A0
timestamp 1644511149
transform -1 0 29900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A
timestamp 1644511149
transform 1 0 28152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A0
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A0
timestamp 1644511149
transform 1 0 30176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A0
timestamp 1644511149
transform -1 0 29808 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A0
timestamp 1644511149
transform 1 0 29532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A0
timestamp 1644511149
transform -1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1644511149
transform 1 0 27048 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A0
timestamp 1644511149
transform 1 0 27508 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A0
timestamp 1644511149
transform 1 0 26772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A0
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A1
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A0
timestamp 1644511149
transform -1 0 28336 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1644511149
transform 1 0 28704 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A0
timestamp 1644511149
transform 1 0 26312 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1644511149
transform 1 0 27784 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A0
timestamp 1644511149
transform 1 0 28152 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1
timestamp 1644511149
transform 1 0 28704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__S
timestamp 1644511149
transform -1 0 28520 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A0
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A1
timestamp 1644511149
transform 1 0 25576 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__S
timestamp 1644511149
transform -1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A_N
timestamp 1644511149
transform -1 0 24564 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A0
timestamp 1644511149
transform -1 0 21804 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1644511149
transform 1 0 24932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S
timestamp 1644511149
transform 1 0 26128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A_N
timestamp 1644511149
transform -1 0 21988 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A0
timestamp 1644511149
transform 1 0 21160 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1
timestamp 1644511149
transform 1 0 24932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__S
timestamp 1644511149
transform -1 0 25944 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A_N
timestamp 1644511149
transform 1 0 22080 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B
timestamp 1644511149
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B1_N
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A1
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1_N
timestamp 1644511149
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A1
timestamp 1644511149
transform 1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1644511149
transform -1 0 20148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A1
timestamp 1644511149
transform 1 0 6256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1
timestamp 1644511149
transform 1 0 6808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1
timestamp 1644511149
transform -1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A1
timestamp 1644511149
transform -1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A1
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A1
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1
timestamp 1644511149
transform -1 0 20516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A1
timestamp 1644511149
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A1
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1644511149
transform 1 0 23736 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A1
timestamp 1644511149
transform 1 0 23736 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1644511149
transform -1 0 27140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1644511149
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A1
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A2
timestamp 1644511149
transform -1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1644511149
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A2
timestamp 1644511149
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1644511149
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1_N
timestamp 1644511149
transform -1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1644511149
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B1_N
timestamp 1644511149
transform -1 0 23276 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A1
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A2
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1644511149
transform -1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__B1_N
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A1
timestamp 1644511149
transform -1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B1_N
timestamp 1644511149
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A1
timestamp 1644511149
transform -1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1_N
timestamp 1644511149
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A1
timestamp 1644511149
transform 1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1644511149
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A1
timestamp 1644511149
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A1
timestamp 1644511149
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A1
timestamp 1644511149
transform -1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1644511149
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A1
timestamp 1644511149
transform 1 0 7360 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1644511149
transform -1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A1
timestamp 1644511149
transform 1 0 9844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A1
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A1
timestamp 1644511149
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A1
timestamp 1644511149
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1644511149
transform -1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A1
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1644511149
transform -1 0 15732 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A1
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1644511149
transform -1 0 13616 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A1
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1644511149
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A1
timestamp 1644511149
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A1
timestamp 1644511149
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A1
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A2
timestamp 1644511149
transform 1 0 26772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A2
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A1
timestamp 1644511149
transform 1 0 27324 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A2
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A1
timestamp 1644511149
transform 1 0 25576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A2
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1644511149
transform 1 0 24472 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A1
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1644511149
transform -1 0 24656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A1
timestamp 1644511149
transform 1 0 30728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A2
timestamp 1644511149
transform 1 0 28520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1644511149
transform 1 0 28152 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1644511149
transform 1 0 28520 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__CLK
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__CLK
timestamp 1644511149
transform 1 0 32844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__CLK
timestamp 1644511149
transform -1 0 36708 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__CLK
timestamp 1644511149
transform 1 0 35328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__CLK
timestamp 1644511149
transform 1 0 36248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__CLK
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__CLK
timestamp 1644511149
transform 1 0 35604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__CLK
timestamp 1644511149
transform 1 0 34040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__CLK
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__CLK
timestamp 1644511149
transform 1 0 32660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__CLK
timestamp 1644511149
transform 1 0 32752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__CLK
timestamp 1644511149
transform -1 0 32936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__CLK
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__CLK
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__CLK
timestamp 1644511149
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__CLK
timestamp 1644511149
transform -1 0 26220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__CLK
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__CLK
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__CLK
timestamp 1644511149
transform 1 0 17296 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1644511149
transform -1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 36800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 37536 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 37444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 37536 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 37536 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 37536 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 37536 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 36800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 36248 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 37444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 36524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 36064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 37444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 36064 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 37444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 38180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 36800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 37444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 23552 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 25852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 27784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 31648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 35972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform -1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 13984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 2852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 2208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 2944 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 2944 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 2208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 2208 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 2208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 2208 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 2208 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 2208 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 2208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 2944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1644511149
transform -1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1644511149
transform -1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1644511149
transform -1 0 2852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1644511149
transform -1 0 2300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1644511149
transform -1 0 2852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1644511149
transform -1 0 2852 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1644511149
transform -1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1644511149
transform -1 0 2484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1644511149
transform -1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1644511149
transform -1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1644511149
transform -1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1644511149
transform -1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1644511149
transform -1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1644511149
transform -1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1644511149
transform -1 0 3220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1644511149
transform -1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1644511149
transform -1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1644511149
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1644511149
transform -1 0 6440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1644511149
transform -1 0 30452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1644511149
transform -1 0 36892 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1644511149
transform -1 0 37444 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1644511149
transform -1 0 37444 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1644511149
transform -1 0 37444 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1644511149
transform -1 0 37444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1644511149
transform -1 0 37444 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1644511149
transform -1 0 26404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1644511149
transform -1 0 26588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1644511149
transform -1 0 27140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1644511149
transform -1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 1644511149
transform -1 0 29716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output129_A
timestamp 1644511149
transform -1 0 32292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output130_A
timestamp 1644511149
transform 1 0 33396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1644511149
transform 1 0 35236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output132_A
timestamp 1644511149
transform 1 0 36248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output140_A
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1644511149
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1644511149
transform 1 0 32844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output163_A
timestamp 1644511149
transform -1 0 2852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1644511149
transform -1 0 3404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1644511149
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output166_A
timestamp 1644511149
transform -1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1644511149
transform 1 0 3312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1644511149
transform 1 0 3496 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1644511149
transform -1 0 2760 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1644511149
transform -1 0 2300 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_158
timestamp 1644511149
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1644511149
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1644511149
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_210
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1644511149
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_263
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1644511149
transform 1 0 28520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1644511149
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_341
timestamp 1644511149
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1644511149
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_379
timestamp 1644511149
transform 1 0 35972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_383
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 1644511149
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_83
timestamp 1644511149
transform 1 0 8740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp 1644511149
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1644511149
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1644511149
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_140
timestamp 1644511149
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_155
timestamp 1644511149
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_171
timestamp 1644511149
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_182
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1644511149
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_227
timestamp 1644511149
transform 1 0 21988 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1644511149
transform 1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_252
timestamp 1644511149
transform 1 0 24288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_263
timestamp 1644511149
transform 1 0 25300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1644511149
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_290
timestamp 1644511149
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_310
timestamp 1644511149
transform 1 0 29624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_316
timestamp 1644511149
transform 1 0 30176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1644511149
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1644511149
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_341
timestamp 1644511149
transform 1 0 32476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_348
timestamp 1644511149
transform 1 0 33120 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_357
timestamp 1644511149
transform 1 0 33948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_364
timestamp 1644511149
transform 1 0 34592 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_372
timestamp 1644511149
transform 1 0 35328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_380
timestamp 1644511149
transform 1 0 36064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_395
timestamp 1644511149
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1644511149
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_45
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1644511149
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_107
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_149 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1644511149
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1644511149
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_222
timestamp 1644511149
transform 1 0 21528 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_260
timestamp 1644511149
transform 1 0 25024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1644511149
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_283
timestamp 1644511149
transform 1 0 27140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_311
timestamp 1644511149
transform 1 0 29716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_315
timestamp 1644511149
transform 1 0 30084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_318
timestamp 1644511149
transform 1 0 30360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_324
timestamp 1644511149
transform 1 0 30912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_341
timestamp 1644511149
transform 1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_347
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_381
timestamp 1644511149
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_387
timestamp 1644511149
transform 1 0 36708 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1644511149
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1644511149
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_98
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_146
timestamp 1644511149
transform 1 0 14536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1644511149
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_176
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_254
timestamp 1644511149
transform 1 0 24472 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_265
timestamp 1644511149
transform 1 0 25484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1644511149
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_289
timestamp 1644511149
transform 1 0 27692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_292
timestamp 1644511149
transform 1 0 27968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_302
timestamp 1644511149
transform 1 0 28888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_309
timestamp 1644511149
transform 1 0 29532 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_327
timestamp 1644511149
transform 1 0 31188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_340
timestamp 1644511149
transform 1 0 32384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_344
timestamp 1644511149
transform 1 0 32752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_347
timestamp 1644511149
transform 1 0 33028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_357
timestamp 1644511149
transform 1 0 33948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_377
timestamp 1644511149
transform 1 0 35788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_383
timestamp 1644511149
transform 1 0 36340 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_402
timestamp 1644511149
transform 1 0 38088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_406
timestamp 1644511149
transform 1 0 38456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1644511149
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_35
timestamp 1644511149
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1644511149
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1644511149
transform 1 0 9108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_99
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_117
timestamp 1644511149
transform 1 0 11868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_148
timestamp 1644511149
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_156
timestamp 1644511149
transform 1 0 15456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1644511149
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_207
timestamp 1644511149
transform 1 0 20148 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_234
timestamp 1644511149
transform 1 0 22632 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_260
timestamp 1644511149
transform 1 0 25024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1644511149
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_280
timestamp 1644511149
transform 1 0 26864 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1644511149
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_325
timestamp 1644511149
transform 1 0 31004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1644511149
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_341
timestamp 1644511149
transform 1 0 32476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1644511149
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 1644511149
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_374
timestamp 1644511149
transform 1 0 35512 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_382
timestamp 1644511149
transform 1 0 36248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_399
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1644511149
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_31
timestamp 1644511149
transform 1 0 3956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1644511149
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_64
timestamp 1644511149
transform 1 0 6992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_76
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1644511149
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1644511149
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_142
timestamp 1644511149
transform 1 0 14168 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_150
timestamp 1644511149
transform 1 0 14904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_155
timestamp 1644511149
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1644511149
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_241
timestamp 1644511149
transform 1 0 23276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1644511149
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_255
timestamp 1644511149
transform 1 0 24564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_264
timestamp 1644511149
transform 1 0 25392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1644511149
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1644511149
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_289
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_299
timestamp 1644511149
transform 1 0 28612 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1644511149
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_319
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1644511149
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_339
timestamp 1644511149
transform 1 0 32292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_347
timestamp 1644511149
transform 1 0 33028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_353
timestamp 1644511149
transform 1 0 33580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_366
timestamp 1644511149
transform 1 0 34776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_376
timestamp 1644511149
transform 1 0 35696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_383
timestamp 1644511149
transform 1 0 36340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1644511149
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_38
timestamp 1644511149
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_49
timestamp 1644511149
transform 1 0 5612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1644511149
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1644511149
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1644511149
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_112
timestamp 1644511149
transform 1 0 11408 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_124
timestamp 1644511149
transform 1 0 12512 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_130
timestamp 1644511149
transform 1 0 13064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1644511149
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1644511149
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_169
timestamp 1644511149
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1644511149
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1644511149
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_204
timestamp 1644511149
transform 1 0 19872 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_216
timestamp 1644511149
transform 1 0 20976 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1644511149
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_225
timestamp 1644511149
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_237
timestamp 1644511149
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_260
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_266
timestamp 1644511149
transform 1 0 25576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1644511149
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_283
timestamp 1644511149
transform 1 0 27140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_295
timestamp 1644511149
transform 1 0 28244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1644511149
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1644511149
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1644511149
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_374
timestamp 1644511149
transform 1 0 35512 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_383
timestamp 1644511149
transform 1 0 36340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_396
timestamp 1644511149
transform 1 0 37536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_29
timestamp 1644511149
transform 1 0 3772 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1644511149
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1644511149
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1644511149
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_64
timestamp 1644511149
transform 1 0 6992 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1644511149
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1644511149
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1644511149
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1644511149
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_121
timestamp 1644511149
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1644511149
transform 1 0 12696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1644511149
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_138
timestamp 1644511149
transform 1 0 13800 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1644511149
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1644511149
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_203
timestamp 1644511149
transform 1 0 19780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_211
timestamp 1644511149
transform 1 0 20516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1644511149
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 1644511149
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_252
timestamp 1644511149
transform 1 0 24288 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_264
timestamp 1644511149
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_365
timestamp 1644511149
transform 1 0 34684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_379
timestamp 1644511149
transform 1 0 35972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_395
timestamp 1644511149
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1644511149
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1644511149
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1644511149
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1644511149
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1644511149
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1644511149
transform 1 0 6440 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_113
timestamp 1644511149
transform 1 0 11500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1644511149
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_128
timestamp 1644511149
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1644511149
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_181
timestamp 1644511149
transform 1 0 17756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1644511149
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_214
timestamp 1644511149
transform 1 0 20792 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_226
timestamp 1644511149
transform 1 0 21896 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_238
timestamp 1644511149
transform 1 0 23000 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1644511149
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_255
timestamp 1644511149
transform 1 0 24564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_267
timestamp 1644511149
transform 1 0 25668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_279
timestamp 1644511149
transform 1 0 26772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_291
timestamp 1644511149
transform 1 0 27876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1644511149
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_318
timestamp 1644511149
transform 1 0 30360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_322
timestamp 1644511149
transform 1 0 30728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1644511149
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_380
timestamp 1644511149
transform 1 0 36064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_387
timestamp 1644511149
transform 1 0 36708 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 1644511149
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_17
timestamp 1644511149
transform 1 0 2668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1644511149
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1644511149
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1644511149
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1644511149
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_59
timestamp 1644511149
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1644511149
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_75
timestamp 1644511149
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1644511149
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_95
timestamp 1644511149
transform 1 0 9844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1644511149
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_133
timestamp 1644511149
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_145
timestamp 1644511149
transform 1 0 14444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1644511149
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1644511149
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_175
timestamp 1644511149
transform 1 0 17204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_187
timestamp 1644511149
transform 1 0 18308 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_207
timestamp 1644511149
transform 1 0 20148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1644511149
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_233
timestamp 1644511149
transform 1 0 22540 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_236
timestamp 1644511149
transform 1 0 22816 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_248
timestamp 1644511149
transform 1 0 23920 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_260
timestamp 1644511149
transform 1 0 25024 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1644511149
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_292
timestamp 1644511149
transform 1 0 27968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_304
timestamp 1644511149
transform 1 0 29072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_308
timestamp 1644511149
transform 1 0 29440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_321
timestamp 1644511149
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1644511149
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_368
timestamp 1644511149
transform 1 0 34960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_374
timestamp 1644511149
transform 1 0 35512 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_384
timestamp 1644511149
transform 1 0 36432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1644511149
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_406
timestamp 1644511149
transform 1 0 38456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1644511149
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1644511149
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_47
timestamp 1644511149
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_59
timestamp 1644511149
transform 1 0 6532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_71
timestamp 1644511149
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1644511149
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1644511149
transform 1 0 10212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1644511149
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_123
timestamp 1644511149
transform 1 0 12420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1644511149
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_169
timestamp 1644511149
transform 1 0 16652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_181
timestamp 1644511149
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1644511149
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_238
timestamp 1644511149
transform 1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1644511149
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_269
timestamp 1644511149
transform 1 0 25852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_286
timestamp 1644511149
transform 1 0 27416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_294
timestamp 1644511149
transform 1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_300
timestamp 1644511149
transform 1 0 28704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_318
timestamp 1644511149
transform 1 0 30360 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_340
timestamp 1644511149
transform 1 0 32384 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_346
timestamp 1644511149
transform 1 0 32936 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1644511149
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_374
timestamp 1644511149
transform 1 0 35512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_381
timestamp 1644511149
transform 1 0 36156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1644511149
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1644511149
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_33
timestamp 1644511149
transform 1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_61
timestamp 1644511149
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1644511149
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_101
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1644511149
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1644511149
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_144
timestamp 1644511149
transform 1 0 14352 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_156
timestamp 1644511149
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_208
timestamp 1644511149
transform 1 0 20240 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1644511149
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1644511149
transform 1 0 22632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_255
timestamp 1644511149
transform 1 0 24564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1644511149
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1644511149
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_290
timestamp 1644511149
transform 1 0 27784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_304
timestamp 1644511149
transform 1 0 29072 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_312
timestamp 1644511149
transform 1 0 29808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1644511149
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_355
timestamp 1644511149
transform 1 0 33764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_368
timestamp 1644511149
transform 1 0 34960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1644511149
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_402
timestamp 1644511149
transform 1 0 38088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1644511149
transform 1 0 38456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1644511149
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_45
timestamp 1644511149
transform 1 0 5244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_57
timestamp 1644511149
transform 1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1644511149
transform 1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_113
timestamp 1644511149
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_124
timestamp 1644511149
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp 1644511149
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1644511149
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_151
timestamp 1644511149
transform 1 0 14996 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_175
timestamp 1644511149
transform 1 0 17204 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_211
timestamp 1644511149
transform 1 0 20516 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1644511149
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1644511149
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_266
timestamp 1644511149
transform 1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_286
timestamp 1644511149
transform 1 0 27416 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_294
timestamp 1644511149
transform 1 0 28152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1644511149
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_313
timestamp 1644511149
transform 1 0 29900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_324
timestamp 1644511149
transform 1 0 30912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_334
timestamp 1644511149
transform 1 0 31832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_340
timestamp 1644511149
transform 1 0 32384 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1644511149
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_371
timestamp 1644511149
transform 1 0 35236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_379
timestamp 1644511149
transform 1 0 35972 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_396
timestamp 1644511149
transform 1 0 37536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1644511149
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1644511149
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_17
timestamp 1644511149
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1644511149
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_46
timestamp 1644511149
transform 1 0 5336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1644511149
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1644511149
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_94
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1644511149
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1644511149
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_143
timestamp 1644511149
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_155
timestamp 1644511149
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1644511149
transform 1 0 19780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_211
timestamp 1644511149
transform 1 0 20516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_233
timestamp 1644511149
transform 1 0 22540 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_243
timestamp 1644511149
transform 1 0 23460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_251
timestamp 1644511149
transform 1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_257
timestamp 1644511149
transform 1 0 24748 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1644511149
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_283
timestamp 1644511149
transform 1 0 27140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_291
timestamp 1644511149
transform 1 0 27876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_299
timestamp 1644511149
transform 1 0 28612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_311
timestamp 1644511149
transform 1 0 29716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_319
timestamp 1644511149
transform 1 0 30452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_324
timestamp 1644511149
transform 1 0 30912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_345
timestamp 1644511149
transform 1 0 32844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_357
timestamp 1644511149
transform 1 0 33948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_369
timestamp 1644511149
transform 1 0 35052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_377
timestamp 1644511149
transform 1 0 35788 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1644511149
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1644511149
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1644511149
transform 1 0 7452 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1644511149
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1644511149
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_117
timestamp 1644511149
transform 1 0 11868 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1644511149
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1644511149
transform 1 0 12972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1644511149
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1644511149
transform 1 0 14260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_151
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_164
timestamp 1644511149
transform 1 0 16192 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1644511149
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1644511149
transform 1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1644511149
transform 1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1644511149
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_235
timestamp 1644511149
transform 1 0 22724 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_241
timestamp 1644511149
transform 1 0 23276 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_256
timestamp 1644511149
transform 1 0 24656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_264
timestamp 1644511149
transform 1 0 25392 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1644511149
transform 1 0 26036 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_285
timestamp 1644511149
transform 1 0 27324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_293
timestamp 1644511149
transform 1 0 28060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1644511149
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_313
timestamp 1644511149
transform 1 0 29900 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_320
timestamp 1644511149
transform 1 0 30544 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_326
timestamp 1644511149
transform 1 0 31096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_343
timestamp 1644511149
transform 1 0 32660 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1644511149
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_373
timestamp 1644511149
transform 1 0 35420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_378
timestamp 1644511149
transform 1 0 35880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_384
timestamp 1644511149
transform 1 0 36432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_400
timestamp 1644511149
transform 1 0 37904 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1644511149
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_19
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_25
timestamp 1644511149
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1644511149
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1644511149
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_92
timestamp 1644511149
transform 1 0 9568 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1644511149
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_119
timestamp 1644511149
transform 1 0 12052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_136
timestamp 1644511149
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_148
timestamp 1644511149
transform 1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_175
timestamp 1644511149
transform 1 0 17204 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1644511149
transform 1 0 18032 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_192
timestamp 1644511149
transform 1 0 18768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_199
timestamp 1644511149
transform 1 0 19412 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_207
timestamp 1644511149
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1644511149
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_235
timestamp 1644511149
transform 1 0 22724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_247
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_263
timestamp 1644511149
transform 1 0 25300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1644511149
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1644511149
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_309
timestamp 1644511149
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_314
timestamp 1644511149
transform 1 0 29992 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1644511149
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1644511149
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_395
timestamp 1644511149
transform 1 0 37444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1644511149
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1644511149
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1644511149
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1644511149
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_129
timestamp 1644511149
transform 1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1644511149
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_161
timestamp 1644511149
transform 1 0 15916 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1644511149
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_172
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1644511149
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_267
timestamp 1644511149
transform 1 0 25668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_273
timestamp 1644511149
transform 1 0 26220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_285
timestamp 1644511149
transform 1 0 27324 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_297
timestamp 1644511149
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1644511149
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_311
timestamp 1644511149
transform 1 0 29716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_324
timestamp 1644511149
transform 1 0 30912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_336
timestamp 1644511149
transform 1 0 32016 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_348
timestamp 1644511149
transform 1 0 33120 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_380
timestamp 1644511149
transform 1 0 36064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_387
timestamp 1644511149
transform 1 0 36708 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1644511149
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_23
timestamp 1644511149
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1644511149
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1644511149
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp 1644511149
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_96
timestamp 1644511149
transform 1 0 9936 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_124
timestamp 1644511149
transform 1 0 12512 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1644511149
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1644511149
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_141
timestamp 1644511149
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_153
timestamp 1644511149
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1644511149
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_209
timestamp 1644511149
transform 1 0 20332 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1644511149
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_312
timestamp 1644511149
transform 1 0 29808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1644511149
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_324
timestamp 1644511149
transform 1 0 30912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_345
timestamp 1644511149
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_359
timestamp 1644511149
transform 1 0 34132 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1644511149
transform 1 0 35972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_402
timestamp 1644511149
transform 1 0 38088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_406
timestamp 1644511149
transform 1 0 38456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_12
timestamp 1644511149
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_20
timestamp 1644511149
transform 1 0 2944 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_38
timestamp 1644511149
transform 1 0 4600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_50
timestamp 1644511149
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_62
timestamp 1644511149
transform 1 0 6808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1644511149
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1644511149
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1644511149
transform 1 0 10764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_117
timestamp 1644511149
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1644511149
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_169
timestamp 1644511149
transform 1 0 16652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_181
timestamp 1644511149
transform 1 0 17756 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1644511149
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1644511149
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_204
timestamp 1644511149
transform 1 0 19872 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_232
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_244
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_259
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1644511149
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1644511149
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_326
timestamp 1644511149
transform 1 0 31096 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_338
timestamp 1644511149
transform 1 0 32200 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_350
timestamp 1644511149
transform 1 0 33304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_356
timestamp 1644511149
transform 1 0 33856 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1644511149
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_371
timestamp 1644511149
transform 1 0 35236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_397
timestamp 1644511149
transform 1 0 37628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_405
timestamp 1644511149
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_25
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_35
timestamp 1644511149
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1644511149
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_88
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1644511149
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1644511149
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1644511149
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1644511149
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1644511149
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_145
timestamp 1644511149
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_177
timestamp 1644511149
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_183
timestamp 1644511149
transform 1 0 17940 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_195
timestamp 1644511149
transform 1 0 19044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_203
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1644511149
transform 1 0 25484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1644511149
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_283
timestamp 1644511149
transform 1 0 27140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_291
timestamp 1644511149
transform 1 0 27876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_296
timestamp 1644511149
transform 1 0 28336 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_306
timestamp 1644511149
transform 1 0 29256 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_323
timestamp 1644511149
transform 1 0 30820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1644511149
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_354
timestamp 1644511149
transform 1 0 33672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_367
timestamp 1644511149
transform 1 0 34868 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_377
timestamp 1644511149
transform 1 0 35788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1644511149
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_395
timestamp 1644511149
transform 1 0 37444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1644511149
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1644511149
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_37
timestamp 1644511149
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_49
timestamp 1644511149
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1644511149
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1644511149
transform 1 0 9660 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1644511149
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_111
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1644511149
transform 1 0 12328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_126
timestamp 1644511149
transform 1 0 12696 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1644511149
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_143
timestamp 1644511149
transform 1 0 14260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_155
timestamp 1644511149
transform 1 0 15364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1644511149
transform 1 0 16468 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_179
timestamp 1644511149
transform 1 0 17572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1644511149
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1644511149
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1644511149
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1644511149
transform 1 0 22080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_234
timestamp 1644511149
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1644511149
transform 1 0 25760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_297
timestamp 1644511149
transform 1 0 28428 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1644511149
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_337
timestamp 1644511149
transform 1 0 32108 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_349
timestamp 1644511149
transform 1 0 33212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_353
timestamp 1644511149
transform 1 0 33580 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1644511149
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_374
timestamp 1644511149
transform 1 0 35512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_380
timestamp 1644511149
transform 1 0 36064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_386
timestamp 1644511149
transform 1 0 36616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_396
timestamp 1644511149
transform 1 0 37536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_9
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_21
timestamp 1644511149
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_33
timestamp 1644511149
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1644511149
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1644511149
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1644511149
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1644511149
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1644511149
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1644511149
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1644511149
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_130
timestamp 1644511149
transform 1 0 13064 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1644511149
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1644511149
transform 1 0 17296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1644511149
transform 1 0 17664 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_183
timestamp 1644511149
transform 1 0 17940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_195
timestamp 1644511149
transform 1 0 19044 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_207
timestamp 1644511149
transform 1 0 20148 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1644511149
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_227
timestamp 1644511149
transform 1 0 21988 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_239
timestamp 1644511149
transform 1 0 23092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_251
timestamp 1644511149
transform 1 0 24196 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1644511149
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1644511149
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1644511149
transform 1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_328
timestamp 1644511149
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_345
timestamp 1644511149
transform 1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_350
timestamp 1644511149
transform 1 0 33304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_363
timestamp 1644511149
transform 1 0 34500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_383
timestamp 1644511149
transform 1 0 36340 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1644511149
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_13
timestamp 1644511149
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1644511149
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_90
timestamp 1644511149
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_102
timestamp 1644511149
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1644511149
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_120
timestamp 1644511149
transform 1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1644511149
transform 1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_166
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1644511149
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1644511149
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1644511149
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_312
timestamp 1644511149
transform 1 0 29808 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_334
timestamp 1644511149
transform 1 0 31832 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_346
timestamp 1644511149
transform 1 0 32936 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1644511149
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_371
timestamp 1644511149
transform 1 0 35236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_383
timestamp 1644511149
transform 1 0 36340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_396
timestamp 1644511149
transform 1 0 37536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_400
timestamp 1644511149
transform 1 0 37904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_6
timestamp 1644511149
transform 1 0 1656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_24
timestamp 1644511149
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1644511149
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_48
timestamp 1644511149
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1644511149
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_122
timestamp 1644511149
transform 1 0 12328 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_130
timestamp 1644511149
transform 1 0 13064 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1644511149
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1644511149
transform 1 0 14076 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_157
timestamp 1644511149
transform 1 0 15548 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1644511149
transform 1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_195
timestamp 1644511149
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1644511149
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_214
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_257
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_262
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_268
timestamp 1644511149
transform 1 0 25760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_272
timestamp 1644511149
transform 1 0 26128 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1644511149
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_311
timestamp 1644511149
transform 1 0 29716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_318
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1644511149
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_368
timestamp 1644511149
transform 1 0 34960 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_378
timestamp 1644511149
transform 1 0 35880 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_395
timestamp 1644511149
transform 1 0 37444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1644511149
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1644511149
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1644511149
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_91
timestamp 1644511149
transform 1 0 9476 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1644511149
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1644511149
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_113
timestamp 1644511149
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1644511149
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1644511149
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_167
timestamp 1644511149
transform 1 0 16468 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_175
timestamp 1644511149
transform 1 0 17204 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_180
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_237
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_256
timestamp 1644511149
transform 1 0 24656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_262
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_271
timestamp 1644511149
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1644511149
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_373
timestamp 1644511149
transform 1 0 35420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_378
timestamp 1644511149
transform 1 0 35880 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_386
timestamp 1644511149
transform 1 0 36616 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_396
timestamp 1644511149
transform 1 0 37536 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_7
timestamp 1644511149
transform 1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_14
timestamp 1644511149
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1644511149
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1644511149
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1644511149
transform 1 0 7636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_91
timestamp 1644511149
transform 1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_97
timestamp 1644511149
transform 1 0 10028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1644511149
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_127
timestamp 1644511149
transform 1 0 12788 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1644511149
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_147
timestamp 1644511149
transform 1 0 14628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1644511149
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1644511149
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_180
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_232
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1644511149
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_248
timestamp 1644511149
transform 1 0 23920 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_256
timestamp 1644511149
transform 1 0 24656 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_265
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_269
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1644511149
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1644511149
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_301
timestamp 1644511149
transform 1 0 28796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_309
timestamp 1644511149
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_321
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1644511149
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_345
timestamp 1644511149
transform 1 0 32844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_358
timestamp 1644511149
transform 1 0 34040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_362
timestamp 1644511149
transform 1 0 34408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_369
timestamp 1644511149
transform 1 0 35052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_377
timestamp 1644511149
transform 1 0 35788 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1644511149
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1644511149
transform 1 0 38180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1644511149
transform 1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_73
timestamp 1644511149
transform 1 0 7820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_93
timestamp 1644511149
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_111
timestamp 1644511149
transform 1 0 11316 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_119
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_181
timestamp 1644511149
transform 1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1644511149
transform 1 0 20884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_230
timestamp 1644511149
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1644511149
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_242
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1644511149
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1644511149
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_320
timestamp 1644511149
transform 1 0 30544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1644511149
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_346
timestamp 1644511149
transform 1 0 32936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_350
timestamp 1644511149
transform 1 0 33304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1644511149
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_374
timestamp 1644511149
transform 1 0 35512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_378
timestamp 1644511149
transform 1 0 35880 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_383
timestamp 1644511149
transform 1 0 36340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_396
timestamp 1644511149
transform 1 0 37536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1644511149
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1644511149
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_25
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_37
timestamp 1644511149
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1644511149
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_94
timestamp 1644511149
transform 1 0 9752 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_138
timestamp 1644511149
transform 1 0 13800 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_146
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_177
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1644511149
transform 1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1644511149
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_242
timestamp 1644511149
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1644511149
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1644511149
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_292
timestamp 1644511149
transform 1 0 27968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_304
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_308
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_315
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1644511149
transform 1 0 31004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_355
timestamp 1644511149
transform 1 0 33764 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_368
timestamp 1644511149
transform 1 0 34960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_374
timestamp 1644511149
transform 1 0 35512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_401
timestamp 1644511149
transform 1 0 37996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_14
timestamp 1644511149
transform 1 0 2392 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_20
timestamp 1644511149
transform 1 0 2944 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_38
timestamp 1644511149
transform 1 0 4600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_50
timestamp 1644511149
transform 1 0 5704 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1644511149
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_71
timestamp 1644511149
transform 1 0 7636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1644511149
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_114
timestamp 1644511149
transform 1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1644511149
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1644511149
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_143
timestamp 1644511149
transform 1 0 14260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_155
timestamp 1644511149
transform 1 0 15364 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_161
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_164
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_181
timestamp 1644511149
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1644511149
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_199
timestamp 1644511149
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1644511149
transform 1 0 20884 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1644511149
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1644511149
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_257
timestamp 1644511149
transform 1 0 24748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_263
timestamp 1644511149
transform 1 0 25300 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_288
timestamp 1644511149
transform 1 0 27600 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_296
timestamp 1644511149
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_311
timestamp 1644511149
transform 1 0 29716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_341
timestamp 1644511149
transform 1 0 32476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_348
timestamp 1644511149
transform 1 0 33120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_356
timestamp 1644511149
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_381
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1644511149
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_85
timestamp 1644511149
transform 1 0 8924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_100
timestamp 1644511149
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_116
timestamp 1644511149
transform 1 0 11776 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_126
timestamp 1644511149
transform 1 0 12696 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_136
timestamp 1644511149
transform 1 0 13616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_148
timestamp 1644511149
transform 1 0 14720 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1644511149
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_199
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1644511149
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_253
timestamp 1644511149
transform 1 0 24380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_264
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_285
timestamp 1644511149
transform 1 0 27324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_309
timestamp 1644511149
transform 1 0 29532 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_313
timestamp 1644511149
transform 1 0 29900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_320
timestamp 1644511149
transform 1 0 30544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1644511149
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_366
timestamp 1644511149
transform 1 0 34776 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_374
timestamp 1644511149
transform 1 0 35512 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_379
timestamp 1644511149
transform 1 0 35972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1644511149
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_395
timestamp 1644511149
transform 1 0 37444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1644511149
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_35
timestamp 1644511149
transform 1 0 4324 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_47
timestamp 1644511149
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_59
timestamp 1644511149
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1644511149
transform 1 0 7636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_117
timestamp 1644511149
transform 1 0 11868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_120
timestamp 1644511149
transform 1 0 12144 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1644511149
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1644511149
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_230
timestamp 1644511149
transform 1 0 22264 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1644511149
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1644511149
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_281
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_287
timestamp 1644511149
transform 1 0 27508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1644511149
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_336
timestamp 1644511149
transform 1 0 32016 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_344
timestamp 1644511149
transform 1 0 32752 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1644511149
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_368
timestamp 1644511149
transform 1 0 34960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_382
timestamp 1644511149
transform 1 0 36248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1644511149
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_22
timestamp 1644511149
transform 1 0 3128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1644511149
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1644511149
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1644511149
transform 1 0 16836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_183
timestamp 1644511149
transform 1 0 17940 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_191
timestamp 1644511149
transform 1 0 18676 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_202
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1644511149
transform 1 0 20424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_246
timestamp 1644511149
transform 1 0 23736 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_258
timestamp 1644511149
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1644511149
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1644511149
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_284
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_292
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_365
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_368
timestamp 1644511149
transform 1 0 34960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1644511149
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_395
timestamp 1644511149
transform 1 0 37444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1644511149
transform 1 0 38180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_13
timestamp 1644511149
transform 1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1644511149
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_31
timestamp 1644511149
transform 1 0 3956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_43
timestamp 1644511149
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_55
timestamp 1644511149
transform 1 0 6164 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_67
timestamp 1644511149
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1644511149
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_127
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_171
timestamp 1644511149
transform 1 0 16836 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_203
timestamp 1644511149
transform 1 0 19780 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1644511149
transform 1 0 20884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1644511149
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_256
timestamp 1644511149
transform 1 0 24656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_268
timestamp 1644511149
transform 1 0 25760 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_280
timestamp 1644511149
transform 1 0 26864 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_286
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1644511149
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_312
timestamp 1644511149
transform 1 0 29808 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_324
timestamp 1644511149
transform 1 0 30912 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_336
timestamp 1644511149
transform 1 0 32016 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_349
timestamp 1644511149
transform 1 0 33212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_383
timestamp 1644511149
transform 1 0 36340 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_391
timestamp 1644511149
transform 1 0 37076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_395
timestamp 1644511149
transform 1 0 37444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1644511149
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1644511149
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_26
timestamp 1644511149
transform 1 0 3496 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_38
timestamp 1644511149
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1644511149
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_133
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1644511149
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_211
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_246
timestamp 1644511149
transform 1 0 23736 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_257
timestamp 1644511149
transform 1 0 24748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1644511149
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_290
timestamp 1644511149
transform 1 0 27784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_302
timestamp 1644511149
transform 1 0 28888 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_308
timestamp 1644511149
transform 1 0 29440 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_348
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_360
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_372
timestamp 1644511149
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_384
timestamp 1644511149
transform 1 0 36432 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_401
timestamp 1644511149
transform 1 0 37996 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1644511149
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1644511149
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1644511149
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_159
timestamp 1644511149
transform 1 0 15732 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1644511149
transform 1 0 24840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_270
timestamp 1644511149
transform 1 0 25944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_278
timestamp 1644511149
transform 1 0 26680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_281
timestamp 1644511149
transform 1 0 26956 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_293
timestamp 1644511149
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1644511149
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_331
timestamp 1644511149
transform 1 0 31556 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_344
timestamp 1644511149
transform 1 0 32752 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_356
timestamp 1644511149
transform 1 0 33856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_374
timestamp 1644511149
transform 1 0 35512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_378
timestamp 1644511149
transform 1 0 35880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_383
timestamp 1644511149
transform 1 0 36340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_396
timestamp 1644511149
transform 1 0 37536 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1644511149
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_12
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_24
timestamp 1644511149
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_36
timestamp 1644511149
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1644511149
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_139
timestamp 1644511149
transform 1 0 13892 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_175
timestamp 1644511149
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1644511149
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_257
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_263
timestamp 1644511149
transform 1 0 25300 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_271
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1644511149
transform 1 0 28520 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_310
timestamp 1644511149
transform 1 0 29624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_315
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_323
timestamp 1644511149
transform 1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_346
timestamp 1644511149
transform 1 0 32936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_360
timestamp 1644511149
transform 1 0 34224 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_379
timestamp 1644511149
transform 1 0 35972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_401
timestamp 1644511149
transform 1 0 37996 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 1644511149
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_241
timestamp 1644511149
transform 1 0 23276 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1644511149
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_258
timestamp 1644511149
transform 1 0 24840 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_264
timestamp 1644511149
transform 1 0 25392 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_326
timestamp 1644511149
transform 1 0 31096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_346
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_371
timestamp 1644511149
transform 1 0 35236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_393
timestamp 1644511149
transform 1 0 37260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1644511149
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_20
timestamp 1644511149
transform 1 0 2944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_26
timestamp 1644511149
transform 1 0 3496 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_38
timestamp 1644511149
transform 1 0 4600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_50
timestamp 1644511149
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_233
timestamp 1644511149
transform 1 0 22540 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_260
timestamp 1644511149
transform 1 0 25024 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_266
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_269
timestamp 1644511149
transform 1 0 25852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_291
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_304
timestamp 1644511149
transform 1 0 29072 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1644511149
transform 1 0 29624 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_322
timestamp 1644511149
transform 1 0 30728 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1644511149
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_343
timestamp 1644511149
transform 1 0 32660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_351
timestamp 1644511149
transform 1 0 33396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_360
timestamp 1644511149
transform 1 0 34224 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_380
timestamp 1644511149
transform 1 0 36064 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_401
timestamp 1644511149
transform 1 0 37996 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_19
timestamp 1644511149
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_229
timestamp 1644511149
transform 1 0 22172 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_238
timestamp 1644511149
transform 1 0 23000 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_256
timestamp 1644511149
transform 1 0 24656 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_268
timestamp 1644511149
transform 1 0 25760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_276
timestamp 1644511149
transform 1 0 26496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_284
timestamp 1644511149
transform 1 0 27232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_371
timestamp 1644511149
transform 1 0 35236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_383
timestamp 1644511149
transform 1 0 36340 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_395
timestamp 1644511149
transform 1 0 37444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_22
timestamp 1644511149
transform 1 0 3128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_28
timestamp 1644511149
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_40
timestamp 1644511149
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1644511149
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_235
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_246
timestamp 1644511149
transform 1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_264
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_272
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_290
timestamp 1644511149
transform 1 0 27784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_296
timestamp 1644511149
transform 1 0 28336 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_302
timestamp 1644511149
transform 1 0 28888 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_314
timestamp 1644511149
transform 1 0 29992 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_326
timestamp 1644511149
transform 1 0 31096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1644511149
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_396
timestamp 1644511149
transform 1 0 37536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1644511149
transform 1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_14
timestamp 1644511149
transform 1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1644511149
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_227
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1644511149
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_261
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_273
timestamp 1644511149
transform 1 0 26220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_284
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1644511149
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_298
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1644511149
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_371
timestamp 1644511149
transform 1 0 35236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_375
timestamp 1644511149
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_382
timestamp 1644511149
transform 1 0 36248 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_386
timestamp 1644511149
transform 1 0 36616 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1644511149
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_13
timestamp 1644511149
transform 1 0 2300 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_31
timestamp 1644511149
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_43
timestamp 1644511149
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_245
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_251
timestamp 1644511149
transform 1 0 24196 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1644511149
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_263
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_271
timestamp 1644511149
transform 1 0 26036 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_290
timestamp 1644511149
transform 1 0 27784 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_296
timestamp 1644511149
transform 1 0 28336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_302
timestamp 1644511149
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_314
timestamp 1644511149
transform 1 0 29992 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_326
timestamp 1644511149
transform 1 0 31096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1644511149
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_342
timestamp 1644511149
transform 1 0 32568 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_354
timestamp 1644511149
transform 1 0 33672 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_366
timestamp 1644511149
transform 1 0 34776 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_395
timestamp 1644511149
transform 1 0 37444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1644511149
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_6
timestamp 1644511149
transform 1 0 1656 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_12
timestamp 1644511149
transform 1 0 2208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_18
timestamp 1644511149
transform 1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1644511149
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_225
timestamp 1644511149
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_235
timestamp 1644511149
transform 1 0 22724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_262
timestamp 1644511149
transform 1 0 25208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_268
timestamp 1644511149
transform 1 0 25760 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_274
timestamp 1644511149
transform 1 0 26312 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_298
timestamp 1644511149
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1644511149
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_317
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_327
timestamp 1644511149
transform 1 0 31188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_340
timestamp 1644511149
transform 1 0 32384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_352
timestamp 1644511149
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_373
timestamp 1644511149
transform 1 0 35420 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_390
timestamp 1644511149
transform 1 0 36984 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_402
timestamp 1644511149
transform 1 0 38088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1644511149
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_9
timestamp 1644511149
transform 1 0 1932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_248
timestamp 1644511149
transform 1 0 23920 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_254
timestamp 1644511149
transform 1 0 24472 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_270
timestamp 1644511149
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1644511149
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_287
timestamp 1644511149
transform 1 0 27508 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_294
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_306
timestamp 1644511149
transform 1 0 29256 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_314
timestamp 1644511149
transform 1 0 29992 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_319
timestamp 1644511149
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_346
timestamp 1644511149
transform 1 0 32936 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_352
timestamp 1644511149
transform 1 0 33488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_358
timestamp 1644511149
transform 1 0 34040 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_366
timestamp 1644511149
transform 1 0 34776 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_370
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_376
timestamp 1644511149
transform 1 0 35696 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_402
timestamp 1644511149
transform 1 0 38088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1644511149
transform 1 0 38456 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_13
timestamp 1644511149
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1644511149
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_234
timestamp 1644511149
transform 1 0 22632 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1644511149
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_255
timestamp 1644511149
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_276
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_296
timestamp 1644511149
transform 1 0 28336 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_319
timestamp 1644511149
transform 1 0 30452 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1644511149
transform 1 0 31372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_336
timestamp 1644511149
transform 1 0 32016 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_349
timestamp 1644511149
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_367
timestamp 1644511149
transform 1 0 34868 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_379
timestamp 1644511149
transform 1 0 35972 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_383
timestamp 1644511149
transform 1 0 36340 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_395
timestamp 1644511149
transform 1 0 37444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1644511149
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_12
timestamp 1644511149
transform 1 0 2208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_24
timestamp 1644511149
transform 1 0 3312 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_36
timestamp 1644511149
transform 1 0 4416 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1644511149
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_229
timestamp 1644511149
transform 1 0 22172 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_254
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_310
timestamp 1644511149
transform 1 0 29624 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_314
timestamp 1644511149
transform 1 0 29992 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_321
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1644511149
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_353
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_372
timestamp 1644511149
transform 1 0 35328 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_384
timestamp 1644511149
transform 1 0 36432 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1644511149
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_396
timestamp 1644511149
transform 1 0 37536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1644511149
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_6
timestamp 1644511149
transform 1 0 1656 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_18
timestamp 1644511149
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1644511149
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_229
timestamp 1644511149
transform 1 0 22172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1644511149
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1644511149
transform 1 0 27048 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_294
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1644511149
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_341
timestamp 1644511149
transform 1 0 32476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_348
timestamp 1644511149
transform 1 0 33120 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_354
timestamp 1644511149
transform 1 0 33672 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1644511149
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_381
timestamp 1644511149
transform 1 0 36156 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1644511149
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1644511149
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_6
timestamp 1644511149
transform 1 0 1656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_12
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_24
timestamp 1644511149
transform 1 0 3312 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_36
timestamp 1644511149
transform 1 0 4416 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 1644511149
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_353
timestamp 1644511149
transform 1 0 33580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_365
timestamp 1644511149
transform 1 0 34684 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_377
timestamp 1644511149
transform 1 0 35788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1644511149
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_395
timestamp 1644511149
transform 1 0 37444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1644511149
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_6
timestamp 1644511149
transform 1 0 1656 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_14
timestamp 1644511149
transform 1 0 2392 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_22
timestamp 1644511149
transform 1 0 3128 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_34
timestamp 1644511149
transform 1 0 4232 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_46
timestamp 1644511149
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1644511149
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1644511149
transform 1 0 38180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_12
timestamp 1644511149
transform 1 0 2208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_6
timestamp 1644511149
transform 1 0 1656 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_18
timestamp 1644511149
transform 1 0 2760 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1644511149
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1644511149
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1644511149
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_396
timestamp 1644511149
transform 1 0 37536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_6
timestamp 1644511149
transform 1 0 1656 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_12
timestamp 1644511149
transform 1 0 2208 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_395
timestamp 1644511149
transform 1 0 37444 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1644511149
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_6
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_12
timestamp 1644511149
transform 1 0 2208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_24
timestamp 1644511149
transform 1 0 3312 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_36
timestamp 1644511149
transform 1 0 4416 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_48
timestamp 1644511149
transform 1 0 5520 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1644511149
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1644511149
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_396
timestamp 1644511149
transform 1 0 37536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1644511149
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1644511149
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1644511149
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_395
timestamp 1644511149
transform 1 0 37444 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_393
timestamp 1644511149
transform 1 0 37260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_396
timestamp 1644511149
transform 1 0 37536 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_18
timestamp 1644511149
transform 1 0 2760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1644511149
transform 1 0 3864 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1644511149
transform 1 0 4968 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1644511149
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_395
timestamp 1644511149
transform 1 0 37444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_6
timestamp 1644511149
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_18
timestamp 1644511149
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_200
timestamp 1644511149
transform 1 0 19504 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_206
timestamp 1644511149
transform 1 0 20056 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_218
timestamp 1644511149
transform 1 0 21160 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_230
timestamp 1644511149
transform 1 0 22264 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_242
timestamp 1644511149
transform 1 0 23368 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1644511149
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1644511149
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_388
timestamp 1644511149
transform 1 0 36800 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1644511149
transform 1 0 37444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_6
timestamp 1644511149
transform 1 0 1656 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_18
timestamp 1644511149
transform 1 0 2760 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1644511149
transform 1 0 3864 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1644511149
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1644511149
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_379
timestamp 1644511149
transform 1 0 35972 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_382
timestamp 1644511149
transform 1 0 36248 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1644511149
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1644511149
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1644511149
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_6
timestamp 1644511149
transform 1 0 1656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_13
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1644511149
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_181
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1644511149
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_210
timestamp 1644511149
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1644511149
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1644511149
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_380
timestamp 1644511149
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_388
timestamp 1644511149
transform 1 0 36800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1644511149
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__nand2b_4  _0454_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  _0455_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0456_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _0457_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0458_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0459_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0460_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0461_
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0462_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0463_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0464_
timestamp 1644511149
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0465_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0466_
timestamp 1644511149
transform 1 0 14260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0467_
timestamp 1644511149
transform -1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0468_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _0469_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_4  _0470_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3956 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__and3b_1  _0471_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11684 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0472_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13524 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0473_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0474_
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0475_
timestamp 1644511149
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _0476_
timestamp 1644511149
transform 1 0 12788 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0477_
timestamp 1644511149
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0478_
timestamp 1644511149
transform -1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _0479_
timestamp 1644511149
transform 1 0 12788 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0480_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19504 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1644511149
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0482_
timestamp 1644511149
transform 1 0 2668 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0483_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0484_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _0485_
timestamp 1644511149
transform 1 0 37628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0486_
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0487_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0488_
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0489_
timestamp 1644511149
transform 1 0 6808 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0490_
timestamp 1644511149
transform 1 0 36340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0491_
timestamp 1644511149
transform 1 0 36984 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_4  _0492_
timestamp 1644511149
transform -1 0 13340 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _0493_
timestamp 1644511149
transform 1 0 35604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0494_
timestamp 1644511149
transform -1 0 36800 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_2  _0495_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 38088 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0496_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0497_
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0498_
timestamp 1644511149
transform 1 0 26404 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0500_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11868 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0501_
timestamp 1644511149
transform -1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0502_
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0503_
timestamp 1644511149
transform -1 0 14996 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0504_
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0505_
timestamp 1644511149
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0506_
timestamp 1644511149
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0507_
timestamp 1644511149
transform -1 0 14260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0508_
timestamp 1644511149
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0509_
timestamp 1644511149
transform 1 0 12604 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0510_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13616 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0511_
timestamp 1644511149
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0512_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0513_
timestamp 1644511149
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0514_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0515_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0516_
timestamp 1644511149
transform -1 0 38088 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0517_
timestamp 1644511149
transform 1 0 26220 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0518_
timestamp 1644511149
transform -1 0 27876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0519_
timestamp 1644511149
transform -1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0520_
timestamp 1644511149
transform 1 0 12052 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0521_
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0522_
timestamp 1644511149
transform -1 0 12880 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0523_
timestamp 1644511149
transform -1 0 10948 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0524_
timestamp 1644511149
transform -1 0 11132 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0525_
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0526_
timestamp 1644511149
transform -1 0 16192 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1644511149
transform 1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0529_
timestamp 1644511149
transform 1 0 11316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0530_
timestamp 1644511149
transform 1 0 11868 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0531_
timestamp 1644511149
transform -1 0 12512 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0532_
timestamp 1644511149
transform -1 0 37536 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0533_
timestamp 1644511149
transform -1 0 27692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0534_
timestamp 1644511149
transform -1 0 10948 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0535_
timestamp 1644511149
transform -1 0 11040 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0536_
timestamp 1644511149
transform 1 0 10488 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0537_
timestamp 1644511149
transform 1 0 11868 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0538_
timestamp 1644511149
transform -1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0539_
timestamp 1644511149
transform -1 0 38088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0540_
timestamp 1644511149
transform -1 0 27968 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0541_
timestamp 1644511149
transform -1 0 9936 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0542_
timestamp 1644511149
transform -1 0 10948 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0543_
timestamp 1644511149
transform -1 0 12052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0544_
timestamp 1644511149
transform -1 0 11500 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0545_
timestamp 1644511149
transform -1 0 12328 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0546_
timestamp 1644511149
transform -1 0 38088 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1644511149
transform -1 0 27784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0548_
timestamp 1644511149
transform 1 0 17020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0549_
timestamp 1644511149
transform -1 0 11040 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0550_
timestamp 1644511149
transform -1 0 11408 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0551_
timestamp 1644511149
transform -1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0552_
timestamp 1644511149
transform 1 0 10396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0553_
timestamp 1644511149
transform 1 0 12880 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0554_
timestamp 1644511149
transform 1 0 11868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0555_
timestamp 1644511149
transform 1 0 20516 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0556_
timestamp 1644511149
transform -1 0 20148 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0557_
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0558_
timestamp 1644511149
transform -1 0 36800 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0559_
timestamp 1644511149
transform 1 0 35880 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_2  _0560_
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0561_
timestamp 1644511149
transform -1 0 28060 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0562_
timestamp 1644511149
transform -1 0 12144 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0563_
timestamp 1644511149
transform 1 0 17940 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0564_
timestamp 1644511149
transform 1 0 15548 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0565_
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1644511149
transform 1 0 14168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0567_
timestamp 1644511149
transform -1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0568_
timestamp 1644511149
transform -1 0 15180 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0569_
timestamp 1644511149
transform -1 0 16192 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0570_
timestamp 1644511149
transform -1 0 37536 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1644511149
transform -1 0 24748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0572_
timestamp 1644511149
transform 1 0 26128 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0573_
timestamp 1644511149
transform -1 0 19320 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0574_
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0575_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0576_
timestamp 1644511149
transform 1 0 17112 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0577_
timestamp 1644511149
transform 1 0 16560 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0578_
timestamp 1644511149
transform 1 0 16744 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1644511149
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1644511149
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0581_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0582_
timestamp 1644511149
transform -1 0 16192 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0583_
timestamp 1644511149
transform -1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0584_
timestamp 1644511149
transform -1 0 37536 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0585_
timestamp 1644511149
transform -1 0 26128 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0586_
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0587_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0588_
timestamp 1644511149
transform 1 0 15272 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0589_
timestamp 1644511149
transform -1 0 17296 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0590_
timestamp 1644511149
transform -1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0591_
timestamp 1644511149
transform -1 0 37536 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0592_
timestamp 1644511149
transform -1 0 26036 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0593_
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0594_
timestamp 1644511149
transform 1 0 17572 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0595_
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0596_
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0597_
timestamp 1644511149
transform 1 0 17020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0598_
timestamp 1644511149
transform -1 0 37536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0599_
timestamp 1644511149
transform -1 0 26036 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0600_
timestamp 1644511149
transform 1 0 19228 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0601_
timestamp 1644511149
transform -1 0 19044 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0602_
timestamp 1644511149
transform -1 0 19872 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0603_
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0604_
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0605_
timestamp 1644511149
transform -1 0 17388 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0606_
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0607_
timestamp 1644511149
transform -1 0 20148 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0608_
timestamp 1644511149
transform -1 0 37536 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0609_
timestamp 1644511149
transform -1 0 36800 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0610_
timestamp 1644511149
transform -1 0 36248 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_2  _0611_
timestamp 1644511149
transform -1 0 37536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0612_
timestamp 1644511149
transform -1 0 26128 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0613_
timestamp 1644511149
transform -1 0 20056 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0614_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0615_
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0616_
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0617_
timestamp 1644511149
transform 1 0 14536 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0618_
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0619_
timestamp 1644511149
transform -1 0 17756 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0620_
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0621_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 37996 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1644511149
transform -1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0623_
timestamp 1644511149
transform -1 0 24840 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0624_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0625_
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0626_
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0627_
timestamp 1644511149
transform 1 0 22172 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0628_
timestamp 1644511149
transform -1 0 22632 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0629_
timestamp 1644511149
transform 1 0 19596 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1644511149
transform 1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0631_
timestamp 1644511149
transform 1 0 16836 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0632_
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0633_
timestamp 1644511149
transform -1 0 21252 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _0634_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0635_
timestamp 1644511149
transform -1 0 36800 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0636_
timestamp 1644511149
transform -1 0 24748 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0637_
timestamp 1644511149
transform -1 0 25024 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0638_
timestamp 1644511149
transform -1 0 25024 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0639_
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0640_
timestamp 1644511149
transform -1 0 21344 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _0641_
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0642_
timestamp 1644511149
transform -1 0 37996 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0643_
timestamp 1644511149
transform -1 0 24748 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0644_
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0645_
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0646_
timestamp 1644511149
transform 1 0 19688 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0647_
timestamp 1644511149
transform -1 0 21252 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _0648_
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0649_
timestamp 1644511149
transform -1 0 37996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0650_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0651_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0652_
timestamp 1644511149
transform 1 0 24656 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0653_
timestamp 1644511149
transform 1 0 23920 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0654_
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0655_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0656_
timestamp 1644511149
transform -1 0 22264 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _0657_
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _0658_
timestamp 1644511149
transform -1 0 38088 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0659_
timestamp 1644511149
transform -1 0 24472 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0660_
timestamp 1644511149
transform 1 0 24840 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0661_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0662_
timestamp 1644511149
transform 1 0 12880 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0663_
timestamp 1644511149
transform 1 0 22816 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0664_
timestamp 1644511149
transform -1 0 22080 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0665_
timestamp 1644511149
transform -1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0666_
timestamp 1644511149
transform -1 0 37444 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0667_
timestamp 1644511149
transform -1 0 23920 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0668_
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0669_
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0670_
timestamp 1644511149
transform 1 0 14444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0671_
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0672_
timestamp 1644511149
transform -1 0 22264 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0673_
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0674_
timestamp 1644511149
transform -1 0 36800 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0675_
timestamp 1644511149
transform -1 0 23736 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0676_
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0677_
timestamp 1644511149
transform 1 0 22264 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0678_
timestamp 1644511149
transform 1 0 22816 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0679_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0680_
timestamp 1644511149
transform -1 0 22724 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0681_
timestamp 1644511149
transform 1 0 37352 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0682_
timestamp 1644511149
transform -1 0 23644 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0683_
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0684_
timestamp 1644511149
transform 1 0 23092 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0685_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0686_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _0687_
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0688_
timestamp 1644511149
transform -1 0 31832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0689_
timestamp 1644511149
transform 1 0 33120 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_2  _0690_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2668 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0691_
timestamp 1644511149
transform 1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0692_
timestamp 1644511149
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0693_
timestamp 1644511149
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0694_
timestamp 1644511149
transform 1 0 33580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0695_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0696_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33580 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform -1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1644511149
transform 1 0 33948 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0699_
timestamp 1644511149
transform -1 0 33948 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1644511149
transform -1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1644511149
transform -1 0 35512 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0702_
timestamp 1644511149
transform 1 0 35144 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 1644511149
transform -1 0 36340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1644511149
transform -1 0 34960 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0705_
timestamp 1644511149
transform 1 0 34408 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1644511149
transform -1 0 35420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0708_
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1644511149
transform -1 0 36156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0710_
timestamp 1644511149
transform 1 0 33120 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0711_
timestamp 1644511149
transform 1 0 33488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1644511149
transform -1 0 34868 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0713_
timestamp 1644511149
transform -1 0 35236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 1644511149
transform -1 0 34224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0716_
timestamp 1644511149
transform 1 0 33672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0717_
timestamp 1644511149
transform -1 0 35788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1644511149
transform -1 0 34500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0719_
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1644511149
transform -1 0 34960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1644511149
transform 1 0 34132 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0722_
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1644511149
transform -1 0 34776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0725_
timestamp 1644511149
transform 1 0 34500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0726_
timestamp 1644511149
transform -1 0 35880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0727_
timestamp 1644511149
transform -1 0 33120 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0728_
timestamp 1644511149
transform -1 0 33212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1644511149
transform 1 0 31924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0730_
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 1644511149
transform 1 0 33304 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0733_
timestamp 1644511149
transform -1 0 32660 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0734_
timestamp 1644511149
transform -1 0 31556 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1644511149
transform 1 0 34592 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0736_
timestamp 1644511149
transform 1 0 33672 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 1644511149
transform -1 0 35604 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1644511149
transform -1 0 35420 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0739_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0740_
timestamp 1644511149
transform 1 0 35972 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0742_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1644511149
transform -1 0 36064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0744_
timestamp 1644511149
transform 1 0 31280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0745_
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0746_
timestamp 1644511149
transform -1 0 31372 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 1644511149
transform -1 0 30636 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0749_
timestamp 1644511149
transform 1 0 31004 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0750_
timestamp 1644511149
transform -1 0 32016 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1644511149
transform 1 0 31556 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0752_
timestamp 1644511149
transform 1 0 29900 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1644511149
transform -1 0 33120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1644511149
transform -1 0 33212 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0755_
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0756_
timestamp 1644511149
transform -1 0 34224 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0757_
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0758_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0759_
timestamp 1644511149
transform 1 0 28244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1644511149
transform -1 0 31188 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0761_
timestamp 1644511149
transform 1 0 31372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1644511149
transform -1 0 32384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0763_
timestamp 1644511149
transform 1 0 27784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0764_
timestamp 1644511149
transform 1 0 28152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1644511149
transform -1 0 29072 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0766_
timestamp 1644511149
transform 1 0 28336 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0767_
timestamp 1644511149
transform -1 0 29532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1644511149
transform 1 0 28980 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0769_
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0770_
timestamp 1644511149
transform 1 0 30176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1644511149
transform 1 0 29808 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0772_
timestamp 1644511149
transform 1 0 29808 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0773_
timestamp 1644511149
transform -1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1644511149
transform 1 0 29900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0775_
timestamp 1644511149
transform 1 0 29808 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 1644511149
transform -1 0 30912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1644511149
transform 1 0 30084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0779_
timestamp 1644511149
transform 1 0 29992 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1644511149
transform -1 0 30912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0781_
timestamp 1644511149
transform 1 0 28152 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1644511149
transform 1 0 29992 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0783_
timestamp 1644511149
transform 1 0 29716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1644511149
transform 1 0 29808 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0786_
timestamp 1644511149
transform -1 0 30360 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0787_
timestamp 1644511149
transform -1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1644511149
transform -1 0 30544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0789_
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1644511149
transform 1 0 30176 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0792_
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0793_
timestamp 1644511149
transform -1 0 31188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0794_
timestamp 1644511149
transform -1 0 27968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1644511149
transform -1 0 28888 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0796_
timestamp 1644511149
transform 1 0 28612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0797_
timestamp 1644511149
transform -1 0 29808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0798_
timestamp 1644511149
transform -1 0 27232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0800_
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1644511149
transform -1 0 26496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1644511149
transform -1 0 27876 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 1644511149
transform -1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 1644511149
transform -1 0 26496 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1644511149
transform 1 0 28244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0806_
timestamp 1644511149
transform 1 0 26680 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1644511149
transform 1 0 27876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0809_
timestamp 1644511149
transform -1 0 27232 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1644511149
transform -1 0 26496 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0812_
timestamp 1644511149
transform -1 0 27508 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1644511149
transform -1 0 26496 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0814_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0816_
timestamp 1644511149
transform 1 0 23000 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0817_
timestamp 1644511149
transform 1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0819_
timestamp 1644511149
transform -1 0 22724 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 1644511149
transform -1 0 22540 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0822_
timestamp 1644511149
transform 1 0 22172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0823_
timestamp 1644511149
transform 1 0 22356 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0824_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0825_
timestamp 1644511149
transform -1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0826_
timestamp 1644511149
transform -1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0827_
timestamp 1644511149
transform -1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0828_
timestamp 1644511149
transform -1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0829_
timestamp 1644511149
transform -1 0 9844 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0830_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0831_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0832_
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0833_
timestamp 1644511149
transform 1 0 4876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0834_
timestamp 1644511149
transform -1 0 19596 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0835_
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0836_
timestamp 1644511149
transform 1 0 6440 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0837_
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0838_
timestamp 1644511149
transform 1 0 6992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0839_
timestamp 1644511149
transform 1 0 7912 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0840_
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0841_
timestamp 1644511149
transform -1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0842_
timestamp 1644511149
transform -1 0 19412 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0843_
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0845_
timestamp 1644511149
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0846_
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0847_
timestamp 1644511149
transform 1 0 19964 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0848_
timestamp 1644511149
transform -1 0 17664 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0849_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0850_
timestamp 1644511149
transform -1 0 18492 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0851_
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0852_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0853_
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0854_
timestamp 1644511149
transform 1 0 20424 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0855_
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0856_
timestamp 1644511149
transform 1 0 21712 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0857_
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0858_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0859_
timestamp 1644511149
transform -1 0 22080 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0860_
timestamp 1644511149
transform -1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1644511149
transform -1 0 24656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0862_
timestamp 1644511149
transform 1 0 24380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0863_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0864_
timestamp 1644511149
transform -1 0 26220 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0865_
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0866_
timestamp 1644511149
transform -1 0 25668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0867_
timestamp 1644511149
transform -1 0 25760 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0868_
timestamp 1644511149
transform -1 0 25576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0869_
timestamp 1644511149
transform -1 0 26036 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0870_
timestamp 1644511149
transform -1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform -1 0 26036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0872_
timestamp 1644511149
transform 1 0 22172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0873_
timestamp 1644511149
transform 1 0 21896 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0874_
timestamp 1644511149
transform 1 0 21804 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0875_
timestamp 1644511149
transform 1 0 22724 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0876_
timestamp 1644511149
transform -1 0 23460 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0877_
timestamp 1644511149
transform -1 0 13800 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0878_
timestamp 1644511149
transform 1 0 11040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0879_
timestamp 1644511149
transform -1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0880_
timestamp 1644511149
transform 1 0 12328 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0881_
timestamp 1644511149
transform -1 0 12420 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0882_
timestamp 1644511149
transform -1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0883_
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0884_
timestamp 1644511149
transform 1 0 3312 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0885_
timestamp 1644511149
transform 1 0 4600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0886_
timestamp 1644511149
transform 1 0 2760 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0887_
timestamp 1644511149
transform 1 0 4140 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0888_
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1644511149
transform 1 0 9108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0890_
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0891_
timestamp 1644511149
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0892_
timestamp 1644511149
transform 1 0 9016 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0893_
timestamp 1644511149
transform 1 0 8004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0894_
timestamp 1644511149
transform -1 0 11040 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0895_
timestamp 1644511149
transform -1 0 11316 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0896_
timestamp 1644511149
transform -1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0897_
timestamp 1644511149
transform 1 0 9568 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0898_
timestamp 1644511149
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0899_
timestamp 1644511149
transform 1 0 9384 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0900_
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0901_
timestamp 1644511149
transform 1 0 7912 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0902_
timestamp 1644511149
transform 1 0 9752 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0903_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0904_
timestamp 1644511149
transform -1 0 8464 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0905_
timestamp 1644511149
transform 1 0 9016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0906_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0907_
timestamp 1644511149
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0908_
timestamp 1644511149
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0909_
timestamp 1644511149
transform -1 0 15456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0910_
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0911_
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0912_
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0913_
timestamp 1644511149
transform 1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0914_
timestamp 1644511149
transform 1 0 14260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0915_
timestamp 1644511149
transform -1 0 19136 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0916_
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0917_
timestamp 1644511149
transform -1 0 18308 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0918_
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0919_
timestamp 1644511149
transform -1 0 17480 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0920_
timestamp 1644511149
transform -1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0921_
timestamp 1644511149
transform -1 0 27968 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0922_
timestamp 1644511149
transform 1 0 26404 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0923_
timestamp 1644511149
transform -1 0 26496 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0924_
timestamp 1644511149
transform 1 0 24748 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0925_
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0926_
timestamp 1644511149
transform 1 0 29072 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0927_
timestamp 1644511149
transform -1 0 29256 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0928_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1644511149
transform 1 0 36340 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1644511149
transform 1 0 35328 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1644511149
transform 1 0 36064 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1644511149
transform 1 0 34500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1644511149
transform 1 0 36156 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1644511149
transform 1 0 34868 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1644511149
transform 1 0 36524 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1644511149
transform -1 0 32936 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1644511149
transform 1 0 35512 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1644511149
transform 1 0 35328 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1644511149
transform -1 0 33580 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1644511149
transform -1 0 32476 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1644511149
transform -1 0 29624 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1644511149
transform 1 0 30820 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1644511149
transform 1 0 30912 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1644511149
transform 1 0 31188 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1644511149
transform 1 0 30360 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1644511149
transform 1 0 30912 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1644511149
transform -1 0 31004 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1644511149
transform 1 0 26404 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1644511149
transform -1 0 28336 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0962_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0963_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0964_
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0965_
timestamp 1644511149
transform 1 0 22264 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1644511149
transform 1 0 6992 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1644511149
transform -1 0 16192 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1644511149
transform -1 0 16652 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1644511149
transform -1 0 17204 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1644511149
transform 1 0 18768 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1644511149
transform 1 0 25392 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1644511149
transform 1 0 27232 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1644511149
transform 1 0 21528 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0984_
timestamp 1644511149
transform 1 0 23000 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1644511149
transform 1 0 2668 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1644511149
transform 1 0 2760 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1644511149
transform 1 0 6624 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1644511149
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1644511149
transform 1 0 7728 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1644511149
transform 1 0 7544 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1644511149
transform 1 0 6992 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0994_
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0995_
timestamp 1644511149
transform -1 0 15916 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0996_
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1644511149
transform 1 0 13984 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0999_
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1644511149
transform 1 0 27508 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1001_
timestamp 1644511149
transform 1 0 26036 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1002_
timestamp 1644511149
transform 1 0 24472 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _1004__181 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1005__182
timestamp 1644511149
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1006__183
timestamp 1644511149
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1007__184
timestamp 1644511149
transform -1 0 1656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1008__185
timestamp 1644511149
transform -1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1009__186
timestamp 1644511149
transform -1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1010__187
timestamp 1644511149
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1011__188
timestamp 1644511149
transform -1 0 1656 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1012__189
timestamp 1644511149
transform -1 0 1656 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1013__190
timestamp 1644511149
transform -1 0 1656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1014__191
timestamp 1644511149
transform -1 0 1656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1015__192
timestamp 1644511149
transform -1 0 1656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1016__193
timestamp 1644511149
transform -1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1017__194
timestamp 1644511149
transform -1 0 2944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21344 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform -1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform -1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform 1 0 31188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform -1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk
timestamp 1644511149
transform -1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk
timestamp 1644511149
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk
timestamp 1644511149
transform -1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk
timestamp 1644511149
transform -1 0 29992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk
timestamp 1644511149
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk
timestamp 1644511149
transform -1 0 28520 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk
timestamp 1644511149
transform 1 0 30728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform -1 0 34592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 37904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 37904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 37904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 37904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 37904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 37904 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 37168 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 36064 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 37904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 36340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform -1 0 36708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform -1 0 36708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 37904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 37904 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 37904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 37904 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1644511149
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform -1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform -1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform -1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform -1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1644511149
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform -1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform -1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform -1 0 2944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform -1 0 2392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform -1 0 2392 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1644511149
transform -1 0 3588 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform -1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform -1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform -1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1644511149
transform 1 0 1472 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1644511149
transform -1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1644511149
transform -1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform -1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input63
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input64
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input65
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input68
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input69
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input72 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input73
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input74
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input75
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1644511149
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input81
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input84
timestamp 1644511149
transform -1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 37812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 37812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 37812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 37812 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 37812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 37812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 37812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 37812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 37812 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 37812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 37812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 37812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 36432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 37076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 37076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 37812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 35972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 35972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 37812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 35972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform -1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform -1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform -1 0 23736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform -1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform -1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1644511149
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1644511149
transform -1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1644511149
transform -1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1644511149
transform -1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1644511149
transform -1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1644511149
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform -1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform -1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 19320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform -1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform -1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform -1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform -1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform -1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform -1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform -1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform -1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform 1 0 20056 0 1 36992
box -38 -48 406 592
<< labels >>
rlabel metal2 s 38934 0 38990 800 6 clk
port 0 nsew signal input
rlabel metal3 s 39200 280 40000 400 6 gpio0_input[0]
port 1 nsew signal input
rlabel metal3 s 39200 21224 40000 21344 6 gpio0_input[10]
port 2 nsew signal input
rlabel metal3 s 39200 23400 40000 23520 6 gpio0_input[11]
port 3 nsew signal input
rlabel metal3 s 39200 25440 40000 25560 6 gpio0_input[12]
port 4 nsew signal input
rlabel metal3 s 39200 27616 40000 27736 6 gpio0_input[13]
port 5 nsew signal input
rlabel metal3 s 39200 29656 40000 29776 6 gpio0_input[14]
port 6 nsew signal input
rlabel metal3 s 39200 31832 40000 31952 6 gpio0_input[15]
port 7 nsew signal input
rlabel metal3 s 39200 33872 40000 33992 6 gpio0_input[16]
port 8 nsew signal input
rlabel metal3 s 39200 36048 40000 36168 6 gpio0_input[17]
port 9 nsew signal input
rlabel metal3 s 39200 38088 40000 38208 6 gpio0_input[18]
port 10 nsew signal input
rlabel metal3 s 39200 2320 40000 2440 6 gpio0_input[1]
port 11 nsew signal input
rlabel metal3 s 39200 4360 40000 4480 6 gpio0_input[2]
port 12 nsew signal input
rlabel metal3 s 39200 6536 40000 6656 6 gpio0_input[3]
port 13 nsew signal input
rlabel metal3 s 39200 8576 40000 8696 6 gpio0_input[4]
port 14 nsew signal input
rlabel metal3 s 39200 10752 40000 10872 6 gpio0_input[5]
port 15 nsew signal input
rlabel metal3 s 39200 12792 40000 12912 6 gpio0_input[6]
port 16 nsew signal input
rlabel metal3 s 39200 14968 40000 15088 6 gpio0_input[7]
port 17 nsew signal input
rlabel metal3 s 39200 17008 40000 17128 6 gpio0_input[8]
port 18 nsew signal input
rlabel metal3 s 39200 19184 40000 19304 6 gpio0_input[9]
port 19 nsew signal input
rlabel metal3 s 39200 960 40000 1080 6 gpio0_oe[0]
port 20 nsew signal tristate
rlabel metal3 s 39200 21904 40000 22024 6 gpio0_oe[10]
port 21 nsew signal tristate
rlabel metal3 s 39200 24080 40000 24200 6 gpio0_oe[11]
port 22 nsew signal tristate
rlabel metal3 s 39200 26120 40000 26240 6 gpio0_oe[12]
port 23 nsew signal tristate
rlabel metal3 s 39200 28296 40000 28416 6 gpio0_oe[13]
port 24 nsew signal tristate
rlabel metal3 s 39200 30336 40000 30456 6 gpio0_oe[14]
port 25 nsew signal tristate
rlabel metal3 s 39200 32512 40000 32632 6 gpio0_oe[15]
port 26 nsew signal tristate
rlabel metal3 s 39200 34552 40000 34672 6 gpio0_oe[16]
port 27 nsew signal tristate
rlabel metal3 s 39200 36728 40000 36848 6 gpio0_oe[17]
port 28 nsew signal tristate
rlabel metal3 s 39200 38768 40000 38888 6 gpio0_oe[18]
port 29 nsew signal tristate
rlabel metal3 s 39200 3000 40000 3120 6 gpio0_oe[1]
port 30 nsew signal tristate
rlabel metal3 s 39200 5176 40000 5296 6 gpio0_oe[2]
port 31 nsew signal tristate
rlabel metal3 s 39200 7216 40000 7336 6 gpio0_oe[3]
port 32 nsew signal tristate
rlabel metal3 s 39200 9392 40000 9512 6 gpio0_oe[4]
port 33 nsew signal tristate
rlabel metal3 s 39200 11432 40000 11552 6 gpio0_oe[5]
port 34 nsew signal tristate
rlabel metal3 s 39200 13608 40000 13728 6 gpio0_oe[6]
port 35 nsew signal tristate
rlabel metal3 s 39200 15648 40000 15768 6 gpio0_oe[7]
port 36 nsew signal tristate
rlabel metal3 s 39200 17688 40000 17808 6 gpio0_oe[8]
port 37 nsew signal tristate
rlabel metal3 s 39200 19864 40000 19984 6 gpio0_oe[9]
port 38 nsew signal tristate
rlabel metal3 s 39200 1640 40000 1760 6 gpio0_output[0]
port 39 nsew signal tristate
rlabel metal3 s 39200 22720 40000 22840 6 gpio0_output[10]
port 40 nsew signal tristate
rlabel metal3 s 39200 24760 40000 24880 6 gpio0_output[11]
port 41 nsew signal tristate
rlabel metal3 s 39200 26936 40000 27056 6 gpio0_output[12]
port 42 nsew signal tristate
rlabel metal3 s 39200 28976 40000 29096 6 gpio0_output[13]
port 43 nsew signal tristate
rlabel metal3 s 39200 31016 40000 31136 6 gpio0_output[14]
port 44 nsew signal tristate
rlabel metal3 s 39200 33192 40000 33312 6 gpio0_output[15]
port 45 nsew signal tristate
rlabel metal3 s 39200 35232 40000 35352 6 gpio0_output[16]
port 46 nsew signal tristate
rlabel metal3 s 39200 37408 40000 37528 6 gpio0_output[17]
port 47 nsew signal tristate
rlabel metal3 s 39200 39448 40000 39568 6 gpio0_output[18]
port 48 nsew signal tristate
rlabel metal3 s 39200 3680 40000 3800 6 gpio0_output[1]
port 49 nsew signal tristate
rlabel metal3 s 39200 5856 40000 5976 6 gpio0_output[2]
port 50 nsew signal tristate
rlabel metal3 s 39200 7896 40000 8016 6 gpio0_output[3]
port 51 nsew signal tristate
rlabel metal3 s 39200 10072 40000 10192 6 gpio0_output[4]
port 52 nsew signal tristate
rlabel metal3 s 39200 12112 40000 12232 6 gpio0_output[5]
port 53 nsew signal tristate
rlabel metal3 s 39200 14288 40000 14408 6 gpio0_output[6]
port 54 nsew signal tristate
rlabel metal3 s 39200 16328 40000 16448 6 gpio0_output[7]
port 55 nsew signal tristate
rlabel metal3 s 39200 18504 40000 18624 6 gpio0_output[8]
port 56 nsew signal tristate
rlabel metal3 s 39200 20544 40000 20664 6 gpio0_output[9]
port 57 nsew signal tristate
rlabel metal2 s 294 0 350 800 6 gpio1_input[0]
port 58 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 gpio1_input[10]
port 59 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 gpio1_input[11]
port 60 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 gpio1_input[12]
port 61 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 gpio1_input[13]
port 62 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 gpio1_input[14]
port 63 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gpio1_input[15]
port 64 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 gpio1_input[16]
port 65 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 gpio1_input[17]
port 66 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 gpio1_input[18]
port 67 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 gpio1_input[1]
port 68 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 gpio1_input[2]
port 69 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 gpio1_input[3]
port 70 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpio1_input[4]
port 71 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 gpio1_input[5]
port 72 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 gpio1_input[6]
port 73 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 gpio1_input[7]
port 74 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 gpio1_input[8]
port 75 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 gpio1_input[9]
port 76 nsew signal input
rlabel metal2 s 938 0 994 800 6 gpio1_oe[0]
port 77 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 gpio1_oe[10]
port 78 nsew signal tristate
rlabel metal2 s 23294 0 23350 800 6 gpio1_oe[11]
port 79 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 gpio1_oe[12]
port 80 nsew signal tristate
rlabel metal2 s 27342 0 27398 800 6 gpio1_oe[13]
port 81 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 gpio1_oe[14]
port 82 nsew signal tristate
rlabel metal2 s 31482 0 31538 800 6 gpio1_oe[15]
port 83 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 gpio1_oe[16]
port 84 nsew signal tristate
rlabel metal2 s 35530 0 35586 800 6 gpio1_oe[17]
port 85 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 gpio1_oe[18]
port 86 nsew signal tristate
rlabel metal2 s 2962 0 3018 800 6 gpio1_oe[1]
port 87 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 gpio1_oe[2]
port 88 nsew signal tristate
rlabel metal2 s 7010 0 7066 800 6 gpio1_oe[3]
port 89 nsew signal tristate
rlabel metal2 s 9034 0 9090 800 6 gpio1_oe[4]
port 90 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 gpio1_oe[5]
port 91 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 gpio1_oe[6]
port 92 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 gpio1_oe[7]
port 93 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 gpio1_oe[8]
port 94 nsew signal tristate
rlabel metal2 s 19246 0 19302 800 6 gpio1_oe[9]
port 95 nsew signal tristate
rlabel metal2 s 1582 0 1638 800 6 gpio1_output[0]
port 96 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 gpio1_output[10]
port 97 nsew signal tristate
rlabel metal2 s 24030 0 24086 800 6 gpio1_output[11]
port 98 nsew signal tristate
rlabel metal2 s 26054 0 26110 800 6 gpio1_output[12]
port 99 nsew signal tristate
rlabel metal2 s 28078 0 28134 800 6 gpio1_output[13]
port 100 nsew signal tristate
rlabel metal2 s 30102 0 30158 800 6 gpio1_output[14]
port 101 nsew signal tristate
rlabel metal2 s 32126 0 32182 800 6 gpio1_output[15]
port 102 nsew signal tristate
rlabel metal2 s 34150 0 34206 800 6 gpio1_output[16]
port 103 nsew signal tristate
rlabel metal2 s 36174 0 36230 800 6 gpio1_output[17]
port 104 nsew signal tristate
rlabel metal2 s 38198 0 38254 800 6 gpio1_output[18]
port 105 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 gpio1_output[1]
port 106 nsew signal tristate
rlabel metal2 s 5630 0 5686 800 6 gpio1_output[2]
port 107 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 gpio1_output[3]
port 108 nsew signal tristate
rlabel metal2 s 9770 0 9826 800 6 gpio1_output[4]
port 109 nsew signal tristate
rlabel metal2 s 11794 0 11850 800 6 gpio1_output[5]
port 110 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 gpio1_output[6]
port 111 nsew signal tristate
rlabel metal2 s 15842 0 15898 800 6 gpio1_output[7]
port 112 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 gpio1_output[8]
port 113 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 gpio1_output[9]
port 114 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 peripheralBus_address[0]
port 115 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 peripheralBus_address[10]
port 116 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 peripheralBus_address[11]
port 117 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 peripheralBus_address[12]
port 118 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 peripheralBus_address[13]
port 119 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 peripheralBus_address[14]
port 120 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 peripheralBus_address[15]
port 121 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 peripheralBus_address[16]
port 122 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 peripheralBus_address[17]
port 123 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 peripheralBus_address[18]
port 124 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 peripheralBus_address[19]
port 125 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 peripheralBus_address[1]
port 126 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 peripheralBus_address[20]
port 127 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 peripheralBus_address[21]
port 128 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 peripheralBus_address[22]
port 129 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 peripheralBus_address[23]
port 130 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 peripheralBus_address[2]
port 131 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 peripheralBus_address[3]
port 132 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 peripheralBus_address[4]
port 133 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 peripheralBus_address[5]
port 134 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 peripheralBus_address[6]
port 135 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 peripheralBus_address[7]
port 136 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 peripheralBus_address[8]
port 137 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 peripheralBus_address[9]
port 138 nsew signal input
rlabel metal3 s 0 144 800 264 6 peripheralBus_busy
port 139 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 peripheralBus_dataIn[0]
port 140 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 peripheralBus_dataIn[10]
port 141 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 peripheralBus_dataIn[11]
port 142 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 peripheralBus_dataIn[12]
port 143 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 peripheralBus_dataIn[13]
port 144 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 peripheralBus_dataIn[14]
port 145 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 peripheralBus_dataIn[15]
port 146 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 peripheralBus_dataIn[16]
port 147 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 peripheralBus_dataIn[17]
port 148 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 peripheralBus_dataIn[18]
port 149 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 peripheralBus_dataIn[19]
port 150 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 peripheralBus_dataIn[1]
port 151 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 peripheralBus_dataIn[20]
port 152 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 peripheralBus_dataIn[21]
port 153 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 peripheralBus_dataIn[22]
port 154 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 peripheralBus_dataIn[23]
port 155 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 peripheralBus_dataIn[24]
port 156 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 peripheralBus_dataIn[25]
port 157 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 peripheralBus_dataIn[26]
port 158 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 peripheralBus_dataIn[27]
port 159 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 peripheralBus_dataIn[28]
port 160 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 peripheralBus_dataIn[29]
port 161 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 peripheralBus_dataIn[2]
port 162 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 peripheralBus_dataIn[30]
port 163 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 peripheralBus_dataIn[31]
port 164 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 peripheralBus_dataIn[3]
port 165 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 peripheralBus_dataIn[4]
port 166 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 peripheralBus_dataIn[5]
port 167 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 peripheralBus_dataIn[6]
port 168 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 peripheralBus_dataIn[7]
port 169 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 peripheralBus_dataIn[8]
port 170 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 peripheralBus_dataIn[9]
port 171 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 peripheralBus_dataOut[0]
port 172 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 peripheralBus_dataOut[10]
port 173 nsew signal tristate
rlabel metal3 s 0 16736 800 16856 6 peripheralBus_dataOut[11]
port 174 nsew signal tristate
rlabel metal3 s 0 18096 800 18216 6 peripheralBus_dataOut[12]
port 175 nsew signal tristate
rlabel metal3 s 0 19456 800 19576 6 peripheralBus_dataOut[13]
port 176 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 peripheralBus_dataOut[14]
port 177 nsew signal tristate
rlabel metal3 s 0 22040 800 22160 6 peripheralBus_dataOut[15]
port 178 nsew signal tristate
rlabel metal3 s 0 23400 800 23520 6 peripheralBus_dataOut[16]
port 179 nsew signal tristate
rlabel metal3 s 0 24624 800 24744 6 peripheralBus_dataOut[17]
port 180 nsew signal tristate
rlabel metal3 s 0 25984 800 26104 6 peripheralBus_dataOut[18]
port 181 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 peripheralBus_dataOut[19]
port 182 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 peripheralBus_dataOut[1]
port 183 nsew signal tristate
rlabel metal3 s 0 28704 800 28824 6 peripheralBus_dataOut[20]
port 184 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 peripheralBus_dataOut[21]
port 185 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 peripheralBus_dataOut[22]
port 186 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 peripheralBus_dataOut[23]
port 187 nsew signal tristate
rlabel metal3 s 0 33464 800 33584 6 peripheralBus_dataOut[24]
port 188 nsew signal tristate
rlabel metal3 s 0 34416 800 34536 6 peripheralBus_dataOut[25]
port 189 nsew signal tristate
rlabel metal3 s 0 35232 800 35352 6 peripheralBus_dataOut[26]
port 190 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 peripheralBus_dataOut[27]
port 191 nsew signal tristate
rlabel metal3 s 0 37000 800 37120 6 peripheralBus_dataOut[28]
port 192 nsew signal tristate
rlabel metal3 s 0 37816 800 37936 6 peripheralBus_dataOut[29]
port 193 nsew signal tristate
rlabel metal3 s 0 4904 800 5024 6 peripheralBus_dataOut[2]
port 194 nsew signal tristate
rlabel metal3 s 0 38768 800 38888 6 peripheralBus_dataOut[30]
port 195 nsew signal tristate
rlabel metal3 s 0 39584 800 39704 6 peripheralBus_dataOut[31]
port 196 nsew signal tristate
rlabel metal3 s 0 6264 800 6384 6 peripheralBus_dataOut[3]
port 197 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 peripheralBus_dataOut[4]
port 198 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 peripheralBus_dataOut[5]
port 199 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 peripheralBus_dataOut[6]
port 200 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 peripheralBus_dataOut[7]
port 201 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 peripheralBus_dataOut[8]
port 202 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 peripheralBus_dataOut[9]
port 203 nsew signal tristate
rlabel metal3 s 0 552 800 672 6 peripheralBus_oe
port 204 nsew signal input
rlabel metal3 s 0 960 800 1080 6 peripheralBus_we
port 205 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 requestOutput
port 206 nsew signal tristate
rlabel metal2 s 39578 0 39634 800 6 rst
port 207 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 208 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 208 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 209 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
