VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 950.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 946.000 4.050 950.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 946.000 82.710 950.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 946.000 90.530 950.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 946.000 98.350 950.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 946.000 106.630 950.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 946.000 114.450 950.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 946.000 122.270 950.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 946.000 130.090 950.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 946.000 137.910 950.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 946.000 145.730 950.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 946.000 154.010 950.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 946.000 11.870 950.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 946.000 161.830 950.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 946.000 169.650 950.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 946.000 177.470 950.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 946.000 185.290 950.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 946.000 193.110 950.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 946.000 200.930 950.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 946.000 209.210 950.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 946.000 217.030 950.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 946.000 224.850 950.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 946.000 232.670 950.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 946.000 19.690 950.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 946.000 240.490 950.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 946.000 248.310 950.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 946.000 256.590 950.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 946.000 264.410 950.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 946.000 272.230 950.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 946.000 280.050 950.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 946.000 287.870 950.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 946.000 295.690 950.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 946.000 27.510 950.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 946.000 35.330 950.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 946.000 43.150 950.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 946.000 50.970 950.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 946.000 59.250 950.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 946.000 67.070 950.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 946.000 74.890 950.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 946.000 303.970 950.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 946.000 382.630 950.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 946.000 390.450 950.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 946.000 398.270 950.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 946.000 406.550 950.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 946.000 414.370 950.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 946.000 422.190 950.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 946.000 430.010 950.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 946.000 437.830 950.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 946.000 445.650 950.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 946.000 453.930 950.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 946.000 311.790 950.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 946.000 461.750 950.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 946.000 469.570 950.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 946.000 477.390 950.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 946.000 485.210 950.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 946.000 493.030 950.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 946.000 500.850 950.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 946.000 509.130 950.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 946.000 516.950 950.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 946.000 524.770 950.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 946.000 532.590 950.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 946.000 319.610 950.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 946.000 540.410 950.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 946.000 548.230 950.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 946.000 556.510 950.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 946.000 564.330 950.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 946.000 572.150 950.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 946.000 579.970 950.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 946.000 587.790 950.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 946.000 595.610 950.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 946.000 327.430 950.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 946.000 335.250 950.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 946.000 343.070 950.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 946.000 350.890 950.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 946.000 359.170 950.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 946.000 366.990 950.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 946.000 374.810 950.000 ;
    END
  END io_out[9]
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 395.120 600.000 395.720 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 553.560 600.000 554.160 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 712.000 600.000 712.600 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 870.440 600.000 871.040 ;
    END
  END jtag_tms
  PIN peripheral_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END peripheral_irq[0]
  PIN peripheral_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END peripheral_irq[1]
  PIN peripheral_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END peripheral_irq[2]
  PIN peripheral_irq[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END peripheral_irq[3]
  PIN peripheral_irq[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END peripheral_irq[4]
  PIN peripheral_irq[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END peripheral_irq[5]
  PIN peripheral_irq[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END peripheral_irq[6]
  PIN peripheral_irq[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END peripheral_irq[7]
  PIN peripheral_irq[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END peripheral_irq[8]
  PIN peripheral_irq[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END peripheral_irq[9]
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 78.920 600.000 79.520 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 236.680 600.000 237.280 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 938.640 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 938.640 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.160 4.000 754.760 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.880 4.000 859.480 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.920 4.000 878.520 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.000 4.000 916.600 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.680 4.000 764.280 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 830.320 4.000 830.920 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 849.360 4.000 849.960 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 906.480 4.000 907.080 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 938.485 ;
      LAYER met1 ;
        RECT 4.210 7.180 595.630 939.040 ;
      LAYER met2 ;
        RECT 4.330 945.720 11.310 946.290 ;
        RECT 12.150 945.720 19.130 946.290 ;
        RECT 19.970 945.720 26.950 946.290 ;
        RECT 27.790 945.720 34.770 946.290 ;
        RECT 35.610 945.720 42.590 946.290 ;
        RECT 43.430 945.720 50.410 946.290 ;
        RECT 51.250 945.720 58.690 946.290 ;
        RECT 59.530 945.720 66.510 946.290 ;
        RECT 67.350 945.720 74.330 946.290 ;
        RECT 75.170 945.720 82.150 946.290 ;
        RECT 82.990 945.720 89.970 946.290 ;
        RECT 90.810 945.720 97.790 946.290 ;
        RECT 98.630 945.720 106.070 946.290 ;
        RECT 106.910 945.720 113.890 946.290 ;
        RECT 114.730 945.720 121.710 946.290 ;
        RECT 122.550 945.720 129.530 946.290 ;
        RECT 130.370 945.720 137.350 946.290 ;
        RECT 138.190 945.720 145.170 946.290 ;
        RECT 146.010 945.720 153.450 946.290 ;
        RECT 154.290 945.720 161.270 946.290 ;
        RECT 162.110 945.720 169.090 946.290 ;
        RECT 169.930 945.720 176.910 946.290 ;
        RECT 177.750 945.720 184.730 946.290 ;
        RECT 185.570 945.720 192.550 946.290 ;
        RECT 193.390 945.720 200.370 946.290 ;
        RECT 201.210 945.720 208.650 946.290 ;
        RECT 209.490 945.720 216.470 946.290 ;
        RECT 217.310 945.720 224.290 946.290 ;
        RECT 225.130 945.720 232.110 946.290 ;
        RECT 232.950 945.720 239.930 946.290 ;
        RECT 240.770 945.720 247.750 946.290 ;
        RECT 248.590 945.720 256.030 946.290 ;
        RECT 256.870 945.720 263.850 946.290 ;
        RECT 264.690 945.720 271.670 946.290 ;
        RECT 272.510 945.720 279.490 946.290 ;
        RECT 280.330 945.720 287.310 946.290 ;
        RECT 288.150 945.720 295.130 946.290 ;
        RECT 295.970 945.720 303.410 946.290 ;
        RECT 304.250 945.720 311.230 946.290 ;
        RECT 312.070 945.720 319.050 946.290 ;
        RECT 319.890 945.720 326.870 946.290 ;
        RECT 327.710 945.720 334.690 946.290 ;
        RECT 335.530 945.720 342.510 946.290 ;
        RECT 343.350 945.720 350.330 946.290 ;
        RECT 351.170 945.720 358.610 946.290 ;
        RECT 359.450 945.720 366.430 946.290 ;
        RECT 367.270 945.720 374.250 946.290 ;
        RECT 375.090 945.720 382.070 946.290 ;
        RECT 382.910 945.720 389.890 946.290 ;
        RECT 390.730 945.720 397.710 946.290 ;
        RECT 398.550 945.720 405.990 946.290 ;
        RECT 406.830 945.720 413.810 946.290 ;
        RECT 414.650 945.720 421.630 946.290 ;
        RECT 422.470 945.720 429.450 946.290 ;
        RECT 430.290 945.720 437.270 946.290 ;
        RECT 438.110 945.720 445.090 946.290 ;
        RECT 445.930 945.720 453.370 946.290 ;
        RECT 454.210 945.720 461.190 946.290 ;
        RECT 462.030 945.720 469.010 946.290 ;
        RECT 469.850 945.720 476.830 946.290 ;
        RECT 477.670 945.720 484.650 946.290 ;
        RECT 485.490 945.720 492.470 946.290 ;
        RECT 493.310 945.720 500.290 946.290 ;
        RECT 501.130 945.720 508.570 946.290 ;
        RECT 509.410 945.720 516.390 946.290 ;
        RECT 517.230 945.720 524.210 946.290 ;
        RECT 525.050 945.720 532.030 946.290 ;
        RECT 532.870 945.720 539.850 946.290 ;
        RECT 540.690 945.720 547.670 946.290 ;
        RECT 548.510 945.720 555.950 946.290 ;
        RECT 556.790 945.720 563.770 946.290 ;
        RECT 564.610 945.720 571.590 946.290 ;
        RECT 572.430 945.720 579.410 946.290 ;
        RECT 580.250 945.720 587.230 946.290 ;
        RECT 588.070 945.720 595.050 946.290 ;
        RECT 4.240 4.280 595.600 945.720 ;
        RECT 4.790 3.670 12.690 4.280 ;
        RECT 13.530 3.670 21.890 4.280 ;
        RECT 22.730 3.670 31.090 4.280 ;
        RECT 31.930 3.670 40.290 4.280 ;
        RECT 41.130 3.670 49.030 4.280 ;
        RECT 49.870 3.670 58.230 4.280 ;
        RECT 59.070 3.670 67.430 4.280 ;
        RECT 68.270 3.670 76.630 4.280 ;
        RECT 77.470 3.670 85.370 4.280 ;
        RECT 86.210 3.670 94.570 4.280 ;
        RECT 95.410 3.670 103.770 4.280 ;
        RECT 104.610 3.670 112.970 4.280 ;
        RECT 113.810 3.670 121.710 4.280 ;
        RECT 122.550 3.670 130.910 4.280 ;
        RECT 131.750 3.670 140.110 4.280 ;
        RECT 140.950 3.670 149.310 4.280 ;
        RECT 150.150 3.670 158.050 4.280 ;
        RECT 158.890 3.670 167.250 4.280 ;
        RECT 168.090 3.670 176.450 4.280 ;
        RECT 177.290 3.670 185.650 4.280 ;
        RECT 186.490 3.670 194.390 4.280 ;
        RECT 195.230 3.670 203.590 4.280 ;
        RECT 204.430 3.670 212.790 4.280 ;
        RECT 213.630 3.670 221.990 4.280 ;
        RECT 222.830 3.670 230.730 4.280 ;
        RECT 231.570 3.670 239.930 4.280 ;
        RECT 240.770 3.670 249.130 4.280 ;
        RECT 249.970 3.670 258.330 4.280 ;
        RECT 259.170 3.670 267.070 4.280 ;
        RECT 267.910 3.670 276.270 4.280 ;
        RECT 277.110 3.670 285.470 4.280 ;
        RECT 286.310 3.670 294.670 4.280 ;
        RECT 295.510 3.670 303.870 4.280 ;
        RECT 304.710 3.670 312.610 4.280 ;
        RECT 313.450 3.670 321.810 4.280 ;
        RECT 322.650 3.670 331.010 4.280 ;
        RECT 331.850 3.670 340.210 4.280 ;
        RECT 341.050 3.670 348.950 4.280 ;
        RECT 349.790 3.670 358.150 4.280 ;
        RECT 358.990 3.670 367.350 4.280 ;
        RECT 368.190 3.670 376.550 4.280 ;
        RECT 377.390 3.670 385.290 4.280 ;
        RECT 386.130 3.670 394.490 4.280 ;
        RECT 395.330 3.670 403.690 4.280 ;
        RECT 404.530 3.670 412.890 4.280 ;
        RECT 413.730 3.670 421.630 4.280 ;
        RECT 422.470 3.670 430.830 4.280 ;
        RECT 431.670 3.670 440.030 4.280 ;
        RECT 440.870 3.670 449.230 4.280 ;
        RECT 450.070 3.670 457.970 4.280 ;
        RECT 458.810 3.670 467.170 4.280 ;
        RECT 468.010 3.670 476.370 4.280 ;
        RECT 477.210 3.670 485.570 4.280 ;
        RECT 486.410 3.670 494.310 4.280 ;
        RECT 495.150 3.670 503.510 4.280 ;
        RECT 504.350 3.670 512.710 4.280 ;
        RECT 513.550 3.670 521.910 4.280 ;
        RECT 522.750 3.670 530.650 4.280 ;
        RECT 531.490 3.670 539.850 4.280 ;
        RECT 540.690 3.670 549.050 4.280 ;
        RECT 549.890 3.670 558.250 4.280 ;
        RECT 559.090 3.670 566.990 4.280 ;
        RECT 567.830 3.670 576.190 4.280 ;
        RECT 577.030 3.670 585.390 4.280 ;
        RECT 586.230 3.670 594.590 4.280 ;
        RECT 595.430 3.670 595.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 944.160 596.000 945.025 ;
        RECT 4.000 936.040 596.000 944.160 ;
        RECT 4.400 934.640 596.000 936.040 ;
        RECT 4.000 926.520 596.000 934.640 ;
        RECT 4.400 925.120 596.000 926.520 ;
        RECT 4.000 917.000 596.000 925.120 ;
        RECT 4.400 915.600 596.000 917.000 ;
        RECT 4.000 907.480 596.000 915.600 ;
        RECT 4.400 906.080 596.000 907.480 ;
        RECT 4.000 897.960 596.000 906.080 ;
        RECT 4.400 896.560 596.000 897.960 ;
        RECT 4.000 888.440 596.000 896.560 ;
        RECT 4.400 887.040 596.000 888.440 ;
        RECT 4.000 878.920 596.000 887.040 ;
        RECT 4.400 877.520 596.000 878.920 ;
        RECT 4.000 871.440 596.000 877.520 ;
        RECT 4.000 870.040 595.600 871.440 ;
        RECT 4.000 869.400 596.000 870.040 ;
        RECT 4.400 868.000 596.000 869.400 ;
        RECT 4.000 859.880 596.000 868.000 ;
        RECT 4.400 858.480 596.000 859.880 ;
        RECT 4.000 850.360 596.000 858.480 ;
        RECT 4.400 848.960 596.000 850.360 ;
        RECT 4.000 840.840 596.000 848.960 ;
        RECT 4.400 839.440 596.000 840.840 ;
        RECT 4.000 831.320 596.000 839.440 ;
        RECT 4.400 829.920 596.000 831.320 ;
        RECT 4.000 821.800 596.000 829.920 ;
        RECT 4.400 820.400 596.000 821.800 ;
        RECT 4.000 812.280 596.000 820.400 ;
        RECT 4.400 810.880 596.000 812.280 ;
        RECT 4.000 802.760 596.000 810.880 ;
        RECT 4.400 801.360 596.000 802.760 ;
        RECT 4.000 793.240 596.000 801.360 ;
        RECT 4.400 791.840 596.000 793.240 ;
        RECT 4.000 783.720 596.000 791.840 ;
        RECT 4.400 782.320 596.000 783.720 ;
        RECT 4.000 774.200 596.000 782.320 ;
        RECT 4.400 772.800 596.000 774.200 ;
        RECT 4.000 764.680 596.000 772.800 ;
        RECT 4.400 763.280 596.000 764.680 ;
        RECT 4.000 755.160 596.000 763.280 ;
        RECT 4.400 753.760 596.000 755.160 ;
        RECT 4.000 745.640 596.000 753.760 ;
        RECT 4.400 744.240 596.000 745.640 ;
        RECT 4.000 736.120 596.000 744.240 ;
        RECT 4.400 734.720 596.000 736.120 ;
        RECT 4.000 726.600 596.000 734.720 ;
        RECT 4.400 725.200 596.000 726.600 ;
        RECT 4.000 717.080 596.000 725.200 ;
        RECT 4.400 715.680 596.000 717.080 ;
        RECT 4.000 713.000 596.000 715.680 ;
        RECT 4.000 711.600 595.600 713.000 ;
        RECT 4.000 707.560 596.000 711.600 ;
        RECT 4.400 706.160 596.000 707.560 ;
        RECT 4.000 698.040 596.000 706.160 ;
        RECT 4.400 696.640 596.000 698.040 ;
        RECT 4.000 688.520 596.000 696.640 ;
        RECT 4.400 687.120 596.000 688.520 ;
        RECT 4.000 679.000 596.000 687.120 ;
        RECT 4.400 677.600 596.000 679.000 ;
        RECT 4.000 669.480 596.000 677.600 ;
        RECT 4.400 668.080 596.000 669.480 ;
        RECT 4.000 659.960 596.000 668.080 ;
        RECT 4.400 658.560 596.000 659.960 ;
        RECT 4.000 650.440 596.000 658.560 ;
        RECT 4.400 649.040 596.000 650.440 ;
        RECT 4.000 640.920 596.000 649.040 ;
        RECT 4.400 639.520 596.000 640.920 ;
        RECT 4.000 632.080 596.000 639.520 ;
        RECT 4.400 630.680 596.000 632.080 ;
        RECT 4.000 622.560 596.000 630.680 ;
        RECT 4.400 621.160 596.000 622.560 ;
        RECT 4.000 613.040 596.000 621.160 ;
        RECT 4.400 611.640 596.000 613.040 ;
        RECT 4.000 603.520 596.000 611.640 ;
        RECT 4.400 602.120 596.000 603.520 ;
        RECT 4.000 594.000 596.000 602.120 ;
        RECT 4.400 592.600 596.000 594.000 ;
        RECT 4.000 584.480 596.000 592.600 ;
        RECT 4.400 583.080 596.000 584.480 ;
        RECT 4.000 574.960 596.000 583.080 ;
        RECT 4.400 573.560 596.000 574.960 ;
        RECT 4.000 565.440 596.000 573.560 ;
        RECT 4.400 564.040 596.000 565.440 ;
        RECT 4.000 555.920 596.000 564.040 ;
        RECT 4.400 554.560 596.000 555.920 ;
        RECT 4.400 554.520 595.600 554.560 ;
        RECT 4.000 553.160 595.600 554.520 ;
        RECT 4.000 546.400 596.000 553.160 ;
        RECT 4.400 545.000 596.000 546.400 ;
        RECT 4.000 536.880 596.000 545.000 ;
        RECT 4.400 535.480 596.000 536.880 ;
        RECT 4.000 527.360 596.000 535.480 ;
        RECT 4.400 525.960 596.000 527.360 ;
        RECT 4.000 517.840 596.000 525.960 ;
        RECT 4.400 516.440 596.000 517.840 ;
        RECT 4.000 508.320 596.000 516.440 ;
        RECT 4.400 506.920 596.000 508.320 ;
        RECT 4.000 498.800 596.000 506.920 ;
        RECT 4.400 497.400 596.000 498.800 ;
        RECT 4.000 489.280 596.000 497.400 ;
        RECT 4.400 487.880 596.000 489.280 ;
        RECT 4.000 479.760 596.000 487.880 ;
        RECT 4.400 478.360 596.000 479.760 ;
        RECT 4.000 470.240 596.000 478.360 ;
        RECT 4.400 468.840 596.000 470.240 ;
        RECT 4.000 460.720 596.000 468.840 ;
        RECT 4.400 459.320 596.000 460.720 ;
        RECT 4.000 451.200 596.000 459.320 ;
        RECT 4.400 449.800 596.000 451.200 ;
        RECT 4.000 441.680 596.000 449.800 ;
        RECT 4.400 440.280 596.000 441.680 ;
        RECT 4.000 432.160 596.000 440.280 ;
        RECT 4.400 430.760 596.000 432.160 ;
        RECT 4.000 422.640 596.000 430.760 ;
        RECT 4.400 421.240 596.000 422.640 ;
        RECT 4.000 413.120 596.000 421.240 ;
        RECT 4.400 411.720 596.000 413.120 ;
        RECT 4.000 403.600 596.000 411.720 ;
        RECT 4.400 402.200 596.000 403.600 ;
        RECT 4.000 396.120 596.000 402.200 ;
        RECT 4.000 394.720 595.600 396.120 ;
        RECT 4.000 394.080 596.000 394.720 ;
        RECT 4.400 392.680 596.000 394.080 ;
        RECT 4.000 384.560 596.000 392.680 ;
        RECT 4.400 383.160 596.000 384.560 ;
        RECT 4.000 375.040 596.000 383.160 ;
        RECT 4.400 373.640 596.000 375.040 ;
        RECT 4.000 365.520 596.000 373.640 ;
        RECT 4.400 364.120 596.000 365.520 ;
        RECT 4.000 356.000 596.000 364.120 ;
        RECT 4.400 354.600 596.000 356.000 ;
        RECT 4.000 346.480 596.000 354.600 ;
        RECT 4.400 345.080 596.000 346.480 ;
        RECT 4.000 336.960 596.000 345.080 ;
        RECT 4.400 335.560 596.000 336.960 ;
        RECT 4.000 327.440 596.000 335.560 ;
        RECT 4.400 326.040 596.000 327.440 ;
        RECT 4.000 318.600 596.000 326.040 ;
        RECT 4.400 317.200 596.000 318.600 ;
        RECT 4.000 309.080 596.000 317.200 ;
        RECT 4.400 307.680 596.000 309.080 ;
        RECT 4.000 299.560 596.000 307.680 ;
        RECT 4.400 298.160 596.000 299.560 ;
        RECT 4.000 290.040 596.000 298.160 ;
        RECT 4.400 288.640 596.000 290.040 ;
        RECT 4.000 280.520 596.000 288.640 ;
        RECT 4.400 279.120 596.000 280.520 ;
        RECT 4.000 271.000 596.000 279.120 ;
        RECT 4.400 269.600 596.000 271.000 ;
        RECT 4.000 261.480 596.000 269.600 ;
        RECT 4.400 260.080 596.000 261.480 ;
        RECT 4.000 251.960 596.000 260.080 ;
        RECT 4.400 250.560 596.000 251.960 ;
        RECT 4.000 242.440 596.000 250.560 ;
        RECT 4.400 241.040 596.000 242.440 ;
        RECT 4.000 237.680 596.000 241.040 ;
        RECT 4.000 236.280 595.600 237.680 ;
        RECT 4.000 232.920 596.000 236.280 ;
        RECT 4.400 231.520 596.000 232.920 ;
        RECT 4.000 223.400 596.000 231.520 ;
        RECT 4.400 222.000 596.000 223.400 ;
        RECT 4.000 213.880 596.000 222.000 ;
        RECT 4.400 212.480 596.000 213.880 ;
        RECT 4.000 204.360 596.000 212.480 ;
        RECT 4.400 202.960 596.000 204.360 ;
        RECT 4.000 194.840 596.000 202.960 ;
        RECT 4.400 193.440 596.000 194.840 ;
        RECT 4.000 185.320 596.000 193.440 ;
        RECT 4.400 183.920 596.000 185.320 ;
        RECT 4.000 175.800 596.000 183.920 ;
        RECT 4.400 174.400 596.000 175.800 ;
        RECT 4.000 166.280 596.000 174.400 ;
        RECT 4.400 164.880 596.000 166.280 ;
        RECT 4.000 156.760 596.000 164.880 ;
        RECT 4.400 155.360 596.000 156.760 ;
        RECT 4.000 147.240 596.000 155.360 ;
        RECT 4.400 145.840 596.000 147.240 ;
        RECT 4.000 137.720 596.000 145.840 ;
        RECT 4.400 136.320 596.000 137.720 ;
        RECT 4.000 128.200 596.000 136.320 ;
        RECT 4.400 126.800 596.000 128.200 ;
        RECT 4.000 118.680 596.000 126.800 ;
        RECT 4.400 117.280 596.000 118.680 ;
        RECT 4.000 109.160 596.000 117.280 ;
        RECT 4.400 107.760 596.000 109.160 ;
        RECT 4.000 99.640 596.000 107.760 ;
        RECT 4.400 98.240 596.000 99.640 ;
        RECT 4.000 90.120 596.000 98.240 ;
        RECT 4.400 88.720 596.000 90.120 ;
        RECT 4.000 80.600 596.000 88.720 ;
        RECT 4.400 79.920 596.000 80.600 ;
        RECT 4.400 79.200 595.600 79.920 ;
        RECT 4.000 78.520 595.600 79.200 ;
        RECT 4.000 71.080 596.000 78.520 ;
        RECT 4.400 69.680 596.000 71.080 ;
        RECT 4.000 61.560 596.000 69.680 ;
        RECT 4.400 60.160 596.000 61.560 ;
        RECT 4.000 52.040 596.000 60.160 ;
        RECT 4.400 50.640 596.000 52.040 ;
        RECT 4.000 42.520 596.000 50.640 ;
        RECT 4.400 41.120 596.000 42.520 ;
        RECT 4.000 33.000 596.000 41.120 ;
        RECT 4.400 31.600 596.000 33.000 ;
        RECT 4.000 23.480 596.000 31.600 ;
        RECT 4.400 22.080 596.000 23.480 ;
        RECT 4.000 13.960 596.000 22.080 ;
        RECT 4.400 12.560 596.000 13.960 ;
        RECT 4.000 5.120 596.000 12.560 ;
        RECT 4.400 4.255 596.000 5.120 ;
      LAYER met4 ;
        RECT 8.575 13.095 20.640 933.465 ;
        RECT 23.040 13.095 97.440 933.465 ;
        RECT 99.840 13.095 174.240 933.465 ;
        RECT 176.640 13.095 251.040 933.465 ;
        RECT 253.440 13.095 327.840 933.465 ;
        RECT 330.240 13.095 404.640 933.465 ;
        RECT 407.040 13.095 481.440 933.465 ;
        RECT 483.840 13.095 558.240 933.465 ;
        RECT 560.640 13.095 580.225 933.465 ;
  END
END Peripherals
END LIBRARY

