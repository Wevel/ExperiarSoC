magic
tech sky130A
magscale 1 2
timestamp 1651272268
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 106 1708 39914 37868
<< metal2 >>
rect 110 39200 166 40000
rect 386 39200 442 40000
rect 754 39200 810 40000
rect 1122 39200 1178 40000
rect 1490 39200 1546 40000
rect 1858 39200 1914 40000
rect 2134 39200 2190 40000
rect 2502 39200 2558 40000
rect 2870 39200 2926 40000
rect 3238 39200 3294 40000
rect 3606 39200 3662 40000
rect 3882 39200 3938 40000
rect 4250 39200 4306 40000
rect 4618 39200 4674 40000
rect 4986 39200 5042 40000
rect 5354 39200 5410 40000
rect 5722 39200 5778 40000
rect 5998 39200 6054 40000
rect 6366 39200 6422 40000
rect 6734 39200 6790 40000
rect 7102 39200 7158 40000
rect 7470 39200 7526 40000
rect 7746 39200 7802 40000
rect 8114 39200 8170 40000
rect 8482 39200 8538 40000
rect 8850 39200 8906 40000
rect 9218 39200 9274 40000
rect 9586 39200 9642 40000
rect 9862 39200 9918 40000
rect 10230 39200 10286 40000
rect 10598 39200 10654 40000
rect 10966 39200 11022 40000
rect 11334 39200 11390 40000
rect 11610 39200 11666 40000
rect 11978 39200 12034 40000
rect 12346 39200 12402 40000
rect 12714 39200 12770 40000
rect 13082 39200 13138 40000
rect 13450 39200 13506 40000
rect 13726 39200 13782 40000
rect 14094 39200 14150 40000
rect 14462 39200 14518 40000
rect 14830 39200 14886 40000
rect 15198 39200 15254 40000
rect 15474 39200 15530 40000
rect 15842 39200 15898 40000
rect 16210 39200 16266 40000
rect 16578 39200 16634 40000
rect 16946 39200 17002 40000
rect 17222 39200 17278 40000
rect 17590 39200 17646 40000
rect 17958 39200 18014 40000
rect 18326 39200 18382 40000
rect 18694 39200 18750 40000
rect 19062 39200 19118 40000
rect 19338 39200 19394 40000
rect 19706 39200 19762 40000
rect 20074 39200 20130 40000
rect 20442 39200 20498 40000
rect 20810 39200 20866 40000
rect 21086 39200 21142 40000
rect 21454 39200 21510 40000
rect 21822 39200 21878 40000
rect 22190 39200 22246 40000
rect 22558 39200 22614 40000
rect 22926 39200 22982 40000
rect 23202 39200 23258 40000
rect 23570 39200 23626 40000
rect 23938 39200 23994 40000
rect 24306 39200 24362 40000
rect 24674 39200 24730 40000
rect 24950 39200 25006 40000
rect 25318 39200 25374 40000
rect 25686 39200 25742 40000
rect 26054 39200 26110 40000
rect 26422 39200 26478 40000
rect 26790 39200 26846 40000
rect 27066 39200 27122 40000
rect 27434 39200 27490 40000
rect 27802 39200 27858 40000
rect 28170 39200 28226 40000
rect 28538 39200 28594 40000
rect 28814 39200 28870 40000
rect 29182 39200 29238 40000
rect 29550 39200 29606 40000
rect 29918 39200 29974 40000
rect 30286 39200 30342 40000
rect 30562 39200 30618 40000
rect 30930 39200 30986 40000
rect 31298 39200 31354 40000
rect 31666 39200 31722 40000
rect 32034 39200 32090 40000
rect 32402 39200 32458 40000
rect 32678 39200 32734 40000
rect 33046 39200 33102 40000
rect 33414 39200 33470 40000
rect 33782 39200 33838 40000
rect 34150 39200 34206 40000
rect 34426 39200 34482 40000
rect 34794 39200 34850 40000
rect 35162 39200 35218 40000
rect 35530 39200 35586 40000
rect 35898 39200 35954 40000
rect 36266 39200 36322 40000
rect 36542 39200 36598 40000
rect 36910 39200 36966 40000
rect 37278 39200 37334 40000
rect 37646 39200 37702 40000
rect 38014 39200 38070 40000
rect 38290 39200 38346 40000
rect 38658 39200 38714 40000
rect 39026 39200 39082 40000
rect 39394 39200 39450 40000
rect 39762 39200 39818 40000
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
<< obsm2 >>
rect 222 39144 330 39250
rect 498 39144 698 39250
rect 866 39144 1066 39250
rect 1234 39144 1434 39250
rect 1602 39144 1802 39250
rect 1970 39144 2078 39250
rect 2246 39144 2446 39250
rect 2614 39144 2814 39250
rect 2982 39144 3182 39250
rect 3350 39144 3550 39250
rect 3718 39144 3826 39250
rect 3994 39144 4194 39250
rect 4362 39144 4562 39250
rect 4730 39144 4930 39250
rect 5098 39144 5298 39250
rect 5466 39144 5666 39250
rect 5834 39144 5942 39250
rect 6110 39144 6310 39250
rect 6478 39144 6678 39250
rect 6846 39144 7046 39250
rect 7214 39144 7414 39250
rect 7582 39144 7690 39250
rect 7858 39144 8058 39250
rect 8226 39144 8426 39250
rect 8594 39144 8794 39250
rect 8962 39144 9162 39250
rect 9330 39144 9530 39250
rect 9698 39144 9806 39250
rect 9974 39144 10174 39250
rect 10342 39144 10542 39250
rect 10710 39144 10910 39250
rect 11078 39144 11278 39250
rect 11446 39144 11554 39250
rect 11722 39144 11922 39250
rect 12090 39144 12290 39250
rect 12458 39144 12658 39250
rect 12826 39144 13026 39250
rect 13194 39144 13394 39250
rect 13562 39144 13670 39250
rect 13838 39144 14038 39250
rect 14206 39144 14406 39250
rect 14574 39144 14774 39250
rect 14942 39144 15142 39250
rect 15310 39144 15418 39250
rect 15586 39144 15786 39250
rect 15954 39144 16154 39250
rect 16322 39144 16522 39250
rect 16690 39144 16890 39250
rect 17058 39144 17166 39250
rect 17334 39144 17534 39250
rect 17702 39144 17902 39250
rect 18070 39144 18270 39250
rect 18438 39144 18638 39250
rect 18806 39144 19006 39250
rect 19174 39144 19282 39250
rect 19450 39144 19650 39250
rect 19818 39144 20018 39250
rect 20186 39144 20386 39250
rect 20554 39144 20754 39250
rect 20922 39144 21030 39250
rect 21198 39144 21398 39250
rect 21566 39144 21766 39250
rect 21934 39144 22134 39250
rect 22302 39144 22502 39250
rect 22670 39144 22870 39250
rect 23038 39144 23146 39250
rect 23314 39144 23514 39250
rect 23682 39144 23882 39250
rect 24050 39144 24250 39250
rect 24418 39144 24618 39250
rect 24786 39144 24894 39250
rect 25062 39144 25262 39250
rect 25430 39144 25630 39250
rect 25798 39144 25998 39250
rect 26166 39144 26366 39250
rect 26534 39144 26734 39250
rect 26902 39144 27010 39250
rect 27178 39144 27378 39250
rect 27546 39144 27746 39250
rect 27914 39144 28114 39250
rect 28282 39144 28482 39250
rect 28650 39144 28758 39250
rect 28926 39144 29126 39250
rect 29294 39144 29494 39250
rect 29662 39144 29862 39250
rect 30030 39144 30230 39250
rect 30398 39144 30506 39250
rect 30674 39144 30874 39250
rect 31042 39144 31242 39250
rect 31410 39144 31610 39250
rect 31778 39144 31978 39250
rect 32146 39144 32346 39250
rect 32514 39144 32622 39250
rect 32790 39144 32990 39250
rect 33158 39144 33358 39250
rect 33526 39144 33726 39250
rect 33894 39144 34094 39250
rect 34262 39144 34370 39250
rect 34538 39144 34738 39250
rect 34906 39144 35106 39250
rect 35274 39144 35474 39250
rect 35642 39144 35842 39250
rect 36010 39144 36210 39250
rect 36378 39144 36486 39250
rect 36654 39144 36854 39250
rect 37022 39144 37222 39250
rect 37390 39144 37590 39250
rect 37758 39144 37958 39250
rect 38126 39144 38234 39250
rect 38402 39144 38602 39250
rect 38770 39144 38970 39250
rect 39138 39144 39338 39250
rect 39506 39144 39706 39250
rect 39874 39144 39908 39250
rect 112 856 39908 39144
rect 222 800 238 856
rect 406 800 514 856
rect 682 800 790 856
rect 958 800 1066 856
rect 1234 800 1342 856
rect 1510 800 1618 856
rect 1786 800 1894 856
rect 2062 800 2170 856
rect 2338 800 2446 856
rect 2614 800 2722 856
rect 2890 800 2998 856
rect 3166 800 3274 856
rect 3442 800 3550 856
rect 3718 800 3826 856
rect 3994 800 4102 856
rect 4270 800 4378 856
rect 4546 800 4654 856
rect 4822 800 4930 856
rect 5098 800 5206 856
rect 5374 800 5482 856
rect 5650 800 5758 856
rect 5926 800 6034 856
rect 6202 800 6310 856
rect 6478 800 6586 856
rect 6754 800 6862 856
rect 7030 800 7138 856
rect 7306 800 7414 856
rect 7582 800 7690 856
rect 7858 800 7966 856
rect 8134 800 8242 856
rect 8410 800 8518 856
rect 8686 800 8794 856
rect 8962 800 9070 856
rect 9238 800 9346 856
rect 9514 800 9622 856
rect 9790 800 9898 856
rect 10066 800 10174 856
rect 10342 800 10450 856
rect 10618 800 10726 856
rect 10894 800 11002 856
rect 11170 800 11278 856
rect 11446 800 11554 856
rect 11722 800 11830 856
rect 11998 800 12106 856
rect 12274 800 12382 856
rect 12550 800 12658 856
rect 12826 800 12934 856
rect 13102 800 13210 856
rect 13378 800 13394 856
rect 13562 800 13670 856
rect 13838 800 13946 856
rect 14114 800 14222 856
rect 14390 800 14498 856
rect 14666 800 14774 856
rect 14942 800 15050 856
rect 15218 800 15326 856
rect 15494 800 15602 856
rect 15770 800 15878 856
rect 16046 800 16154 856
rect 16322 800 16430 856
rect 16598 800 16706 856
rect 16874 800 16982 856
rect 17150 800 17258 856
rect 17426 800 17534 856
rect 17702 800 17810 856
rect 17978 800 18086 856
rect 18254 800 18362 856
rect 18530 800 18638 856
rect 18806 800 18914 856
rect 19082 800 19190 856
rect 19358 800 19466 856
rect 19634 800 19742 856
rect 19910 800 20018 856
rect 20186 800 20294 856
rect 20462 800 20570 856
rect 20738 800 20846 856
rect 21014 800 21122 856
rect 21290 800 21398 856
rect 21566 800 21674 856
rect 21842 800 21950 856
rect 22118 800 22226 856
rect 22394 800 22502 856
rect 22670 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23330 856
rect 23498 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24158 856
rect 24326 800 24434 856
rect 24602 800 24710 856
rect 24878 800 24986 856
rect 25154 800 25262 856
rect 25430 800 25538 856
rect 25706 800 25814 856
rect 25982 800 26090 856
rect 26258 800 26366 856
rect 26534 800 26642 856
rect 26810 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27378 856
rect 27546 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28206 856
rect 28374 800 28482 856
rect 28650 800 28758 856
rect 28926 800 29034 856
rect 29202 800 29310 856
rect 29478 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30138 856
rect 30306 800 30414 856
rect 30582 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31242 856
rect 31410 800 31518 856
rect 31686 800 31794 856
rect 31962 800 32070 856
rect 32238 800 32346 856
rect 32514 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33174 856
rect 33342 800 33450 856
rect 33618 800 33726 856
rect 33894 800 34002 856
rect 34170 800 34278 856
rect 34446 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35106 856
rect 35274 800 35382 856
rect 35550 800 35658 856
rect 35826 800 35934 856
rect 36102 800 36210 856
rect 36378 800 36486 856
rect 36654 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37314 856
rect 37482 800 37590 856
rect 37758 800 37866 856
rect 38034 800 38142 856
rect 38310 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38970 856
rect 39138 800 39246 856
rect 39414 800 39522 856
rect 39690 800 39798 856
<< metal3 >>
rect 39200 39040 40000 39160
rect 39200 37408 40000 37528
rect 39200 35776 40000 35896
rect 39200 34144 40000 34264
rect 39200 32376 40000 32496
rect 39200 30744 40000 30864
rect 0 29928 800 30048
rect 39200 29112 40000 29232
rect 39200 27480 40000 27600
rect 39200 25712 40000 25832
rect 39200 24080 40000 24200
rect 39200 22448 40000 22568
rect 39200 20816 40000 20936
rect 39200 19048 40000 19168
rect 39200 17416 40000 17536
rect 39200 15784 40000 15904
rect 39200 14152 40000 14272
rect 39200 12384 40000 12504
rect 39200 10752 40000 10872
rect 0 9936 800 10056
rect 39200 9120 40000 9240
rect 39200 7488 40000 7608
rect 39200 5720 40000 5840
rect 39200 4088 40000 4208
rect 39200 2456 40000 2576
rect 39200 824 40000 944
<< obsm3 >>
rect 800 38960 39120 39133
rect 800 37608 39200 38960
rect 800 37328 39120 37608
rect 800 35976 39200 37328
rect 800 35696 39120 35976
rect 800 34344 39200 35696
rect 800 34064 39120 34344
rect 800 32576 39200 34064
rect 800 32296 39120 32576
rect 800 30944 39200 32296
rect 800 30664 39120 30944
rect 800 30128 39200 30664
rect 880 29848 39200 30128
rect 800 29312 39200 29848
rect 800 29032 39120 29312
rect 800 27680 39200 29032
rect 800 27400 39120 27680
rect 800 25912 39200 27400
rect 800 25632 39120 25912
rect 800 24280 39200 25632
rect 800 24000 39120 24280
rect 800 22648 39200 24000
rect 800 22368 39120 22648
rect 800 21016 39200 22368
rect 800 20736 39120 21016
rect 800 19248 39200 20736
rect 800 18968 39120 19248
rect 800 17616 39200 18968
rect 800 17336 39120 17616
rect 800 15984 39200 17336
rect 800 15704 39120 15984
rect 800 14352 39200 15704
rect 800 14072 39120 14352
rect 800 12584 39200 14072
rect 800 12304 39120 12584
rect 800 10952 39200 12304
rect 800 10672 39120 10952
rect 800 10136 39200 10672
rect 880 9856 39200 10136
rect 800 9320 39200 9856
rect 800 9040 39120 9320
rect 800 7688 39200 9040
rect 800 7408 39120 7688
rect 800 5920 39200 7408
rect 800 5640 39120 5920
rect 800 4288 39200 5640
rect 800 4008 39120 4288
rect 800 2656 39200 4008
rect 800 2376 39120 2656
rect 800 1024 39200 2376
rect 800 851 39120 1024
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 0 9936 800 10056 6 clk
port 1 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 gpio0_input[0]
port 2 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 gpio0_input[10]
port 3 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 gpio0_input[11]
port 4 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 gpio0_input[12]
port 5 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 gpio0_input[13]
port 6 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 gpio0_input[14]
port 7 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 gpio0_input[15]
port 8 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 gpio0_input[16]
port 9 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 gpio0_input[17]
port 10 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 gpio0_input[18]
port 11 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 gpio0_input[1]
port 12 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 gpio0_input[2]
port 13 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 gpio0_input[3]
port 14 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 gpio0_input[4]
port 15 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 gpio0_input[5]
port 16 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 gpio0_input[6]
port 17 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 gpio0_input[7]
port 18 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 gpio0_input[8]
port 19 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 gpio0_input[9]
port 20 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 gpio0_oe[0]
port 21 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 gpio0_oe[10]
port 22 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 gpio0_oe[11]
port 23 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 gpio0_oe[12]
port 24 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 gpio0_oe[13]
port 25 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 gpio0_oe[14]
port 26 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 gpio0_oe[15]
port 27 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 gpio0_oe[16]
port 28 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 gpio0_oe[17]
port 29 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 gpio0_oe[18]
port 30 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 gpio0_oe[1]
port 31 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 gpio0_oe[2]
port 32 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 gpio0_oe[3]
port 33 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 gpio0_oe[4]
port 34 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 gpio0_oe[5]
port 35 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 gpio0_oe[6]
port 36 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 gpio0_oe[7]
port 37 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 gpio0_oe[8]
port 38 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 gpio0_oe[9]
port 39 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 gpio0_output[0]
port 40 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 gpio0_output[10]
port 41 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 gpio0_output[11]
port 42 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 gpio0_output[12]
port 43 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 gpio0_output[13]
port 44 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 gpio0_output[14]
port 45 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 gpio0_output[15]
port 46 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 gpio0_output[16]
port 47 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 gpio0_output[17]
port 48 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 gpio0_output[18]
port 49 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 gpio0_output[1]
port 50 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 gpio0_output[2]
port 51 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 gpio0_output[3]
port 52 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 gpio0_output[4]
port 53 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 gpio0_output[5]
port 54 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 gpio0_output[6]
port 55 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gpio0_output[7]
port 56 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 gpio0_output[8]
port 57 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 gpio0_output[9]
port 58 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 gpio1_input[0]
port 59 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 gpio1_input[10]
port 60 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 gpio1_input[11]
port 61 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 gpio1_input[12]
port 62 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 gpio1_input[13]
port 63 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 gpio1_input[14]
port 64 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 gpio1_input[15]
port 65 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 gpio1_input[16]
port 66 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 gpio1_input[17]
port 67 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 gpio1_input[18]
port 68 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 gpio1_input[1]
port 69 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 gpio1_input[2]
port 70 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 gpio1_input[3]
port 71 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 gpio1_input[4]
port 72 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 gpio1_input[5]
port 73 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 gpio1_input[6]
port 74 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 gpio1_input[7]
port 75 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 gpio1_input[8]
port 76 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 gpio1_input[9]
port 77 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 gpio1_oe[0]
port 78 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 gpio1_oe[10]
port 79 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 gpio1_oe[11]
port 80 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 gpio1_oe[12]
port 81 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 gpio1_oe[13]
port 82 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 gpio1_oe[14]
port 83 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 gpio1_oe[15]
port 84 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 gpio1_oe[16]
port 85 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 gpio1_oe[17]
port 86 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 gpio1_oe[18]
port 87 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 gpio1_oe[1]
port 88 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 gpio1_oe[2]
port 89 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 gpio1_oe[3]
port 90 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 gpio1_oe[4]
port 91 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 gpio1_oe[5]
port 92 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 gpio1_oe[6]
port 93 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 gpio1_oe[7]
port 94 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 gpio1_oe[8]
port 95 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 gpio1_oe[9]
port 96 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 gpio1_output[0]
port 97 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 gpio1_output[10]
port 98 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 gpio1_output[11]
port 99 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 gpio1_output[12]
port 100 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 gpio1_output[13]
port 101 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 gpio1_output[14]
port 102 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 gpio1_output[15]
port 103 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 gpio1_output[16]
port 104 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 gpio1_output[17]
port 105 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 gpio1_output[18]
port 106 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 gpio1_output[1]
port 107 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 gpio1_output[2]
port 108 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 gpio1_output[3]
port 109 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 gpio1_output[4]
port 110 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 gpio1_output[5]
port 111 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 gpio1_output[6]
port 112 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 gpio1_output[7]
port 113 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 gpio1_output[8]
port 114 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 gpio1_output[9]
port 115 nsew signal input
rlabel metal2 s 110 39200 166 40000 6 io_in[0]
port 116 nsew signal input
rlabel metal2 s 10598 39200 10654 40000 6 io_in[10]
port 117 nsew signal input
rlabel metal2 s 11610 39200 11666 40000 6 io_in[11]
port 118 nsew signal input
rlabel metal2 s 12714 39200 12770 40000 6 io_in[12]
port 119 nsew signal input
rlabel metal2 s 13726 39200 13782 40000 6 io_in[13]
port 120 nsew signal input
rlabel metal2 s 14830 39200 14886 40000 6 io_in[14]
port 121 nsew signal input
rlabel metal2 s 15842 39200 15898 40000 6 io_in[15]
port 122 nsew signal input
rlabel metal2 s 16946 39200 17002 40000 6 io_in[16]
port 123 nsew signal input
rlabel metal2 s 17958 39200 18014 40000 6 io_in[17]
port 124 nsew signal input
rlabel metal2 s 19062 39200 19118 40000 6 io_in[18]
port 125 nsew signal input
rlabel metal2 s 20074 39200 20130 40000 6 io_in[19]
port 126 nsew signal input
rlabel metal2 s 1122 39200 1178 40000 6 io_in[1]
port 127 nsew signal input
rlabel metal2 s 21086 39200 21142 40000 6 io_in[20]
port 128 nsew signal input
rlabel metal2 s 22190 39200 22246 40000 6 io_in[21]
port 129 nsew signal input
rlabel metal2 s 23202 39200 23258 40000 6 io_in[22]
port 130 nsew signal input
rlabel metal2 s 24306 39200 24362 40000 6 io_in[23]
port 131 nsew signal input
rlabel metal2 s 25318 39200 25374 40000 6 io_in[24]
port 132 nsew signal input
rlabel metal2 s 26422 39200 26478 40000 6 io_in[25]
port 133 nsew signal input
rlabel metal2 s 27434 39200 27490 40000 6 io_in[26]
port 134 nsew signal input
rlabel metal2 s 28538 39200 28594 40000 6 io_in[27]
port 135 nsew signal input
rlabel metal2 s 29550 39200 29606 40000 6 io_in[28]
port 136 nsew signal input
rlabel metal2 s 30562 39200 30618 40000 6 io_in[29]
port 137 nsew signal input
rlabel metal2 s 2134 39200 2190 40000 6 io_in[2]
port 138 nsew signal input
rlabel metal2 s 31666 39200 31722 40000 6 io_in[30]
port 139 nsew signal input
rlabel metal2 s 32678 39200 32734 40000 6 io_in[31]
port 140 nsew signal input
rlabel metal2 s 33782 39200 33838 40000 6 io_in[32]
port 141 nsew signal input
rlabel metal2 s 34794 39200 34850 40000 6 io_in[33]
port 142 nsew signal input
rlabel metal2 s 35898 39200 35954 40000 6 io_in[34]
port 143 nsew signal input
rlabel metal2 s 36910 39200 36966 40000 6 io_in[35]
port 144 nsew signal input
rlabel metal2 s 38014 39200 38070 40000 6 io_in[36]
port 145 nsew signal input
rlabel metal2 s 39026 39200 39082 40000 6 io_in[37]
port 146 nsew signal input
rlabel metal2 s 3238 39200 3294 40000 6 io_in[3]
port 147 nsew signal input
rlabel metal2 s 4250 39200 4306 40000 6 io_in[4]
port 148 nsew signal input
rlabel metal2 s 5354 39200 5410 40000 6 io_in[5]
port 149 nsew signal input
rlabel metal2 s 6366 39200 6422 40000 6 io_in[6]
port 150 nsew signal input
rlabel metal2 s 7470 39200 7526 40000 6 io_in[7]
port 151 nsew signal input
rlabel metal2 s 8482 39200 8538 40000 6 io_in[8]
port 152 nsew signal input
rlabel metal2 s 9586 39200 9642 40000 6 io_in[9]
port 153 nsew signal input
rlabel metal2 s 386 39200 442 40000 6 io_oeb[0]
port 154 nsew signal output
rlabel metal2 s 10966 39200 11022 40000 6 io_oeb[10]
port 155 nsew signal output
rlabel metal2 s 11978 39200 12034 40000 6 io_oeb[11]
port 156 nsew signal output
rlabel metal2 s 13082 39200 13138 40000 6 io_oeb[12]
port 157 nsew signal output
rlabel metal2 s 14094 39200 14150 40000 6 io_oeb[13]
port 158 nsew signal output
rlabel metal2 s 15198 39200 15254 40000 6 io_oeb[14]
port 159 nsew signal output
rlabel metal2 s 16210 39200 16266 40000 6 io_oeb[15]
port 160 nsew signal output
rlabel metal2 s 17222 39200 17278 40000 6 io_oeb[16]
port 161 nsew signal output
rlabel metal2 s 18326 39200 18382 40000 6 io_oeb[17]
port 162 nsew signal output
rlabel metal2 s 19338 39200 19394 40000 6 io_oeb[18]
port 163 nsew signal output
rlabel metal2 s 20442 39200 20498 40000 6 io_oeb[19]
port 164 nsew signal output
rlabel metal2 s 1490 39200 1546 40000 6 io_oeb[1]
port 165 nsew signal output
rlabel metal2 s 21454 39200 21510 40000 6 io_oeb[20]
port 166 nsew signal output
rlabel metal2 s 22558 39200 22614 40000 6 io_oeb[21]
port 167 nsew signal output
rlabel metal2 s 23570 39200 23626 40000 6 io_oeb[22]
port 168 nsew signal output
rlabel metal2 s 24674 39200 24730 40000 6 io_oeb[23]
port 169 nsew signal output
rlabel metal2 s 25686 39200 25742 40000 6 io_oeb[24]
port 170 nsew signal output
rlabel metal2 s 26790 39200 26846 40000 6 io_oeb[25]
port 171 nsew signal output
rlabel metal2 s 27802 39200 27858 40000 6 io_oeb[26]
port 172 nsew signal output
rlabel metal2 s 28814 39200 28870 40000 6 io_oeb[27]
port 173 nsew signal output
rlabel metal2 s 29918 39200 29974 40000 6 io_oeb[28]
port 174 nsew signal output
rlabel metal2 s 30930 39200 30986 40000 6 io_oeb[29]
port 175 nsew signal output
rlabel metal2 s 2502 39200 2558 40000 6 io_oeb[2]
port 176 nsew signal output
rlabel metal2 s 32034 39200 32090 40000 6 io_oeb[30]
port 177 nsew signal output
rlabel metal2 s 33046 39200 33102 40000 6 io_oeb[31]
port 178 nsew signal output
rlabel metal2 s 34150 39200 34206 40000 6 io_oeb[32]
port 179 nsew signal output
rlabel metal2 s 35162 39200 35218 40000 6 io_oeb[33]
port 180 nsew signal output
rlabel metal2 s 36266 39200 36322 40000 6 io_oeb[34]
port 181 nsew signal output
rlabel metal2 s 37278 39200 37334 40000 6 io_oeb[35]
port 182 nsew signal output
rlabel metal2 s 38290 39200 38346 40000 6 io_oeb[36]
port 183 nsew signal output
rlabel metal2 s 39394 39200 39450 40000 6 io_oeb[37]
port 184 nsew signal output
rlabel metal2 s 3606 39200 3662 40000 6 io_oeb[3]
port 185 nsew signal output
rlabel metal2 s 4618 39200 4674 40000 6 io_oeb[4]
port 186 nsew signal output
rlabel metal2 s 5722 39200 5778 40000 6 io_oeb[5]
port 187 nsew signal output
rlabel metal2 s 6734 39200 6790 40000 6 io_oeb[6]
port 188 nsew signal output
rlabel metal2 s 7746 39200 7802 40000 6 io_oeb[7]
port 189 nsew signal output
rlabel metal2 s 8850 39200 8906 40000 6 io_oeb[8]
port 190 nsew signal output
rlabel metal2 s 9862 39200 9918 40000 6 io_oeb[9]
port 191 nsew signal output
rlabel metal2 s 754 39200 810 40000 6 io_out[0]
port 192 nsew signal output
rlabel metal2 s 11334 39200 11390 40000 6 io_out[10]
port 193 nsew signal output
rlabel metal2 s 12346 39200 12402 40000 6 io_out[11]
port 194 nsew signal output
rlabel metal2 s 13450 39200 13506 40000 6 io_out[12]
port 195 nsew signal output
rlabel metal2 s 14462 39200 14518 40000 6 io_out[13]
port 196 nsew signal output
rlabel metal2 s 15474 39200 15530 40000 6 io_out[14]
port 197 nsew signal output
rlabel metal2 s 16578 39200 16634 40000 6 io_out[15]
port 198 nsew signal output
rlabel metal2 s 17590 39200 17646 40000 6 io_out[16]
port 199 nsew signal output
rlabel metal2 s 18694 39200 18750 40000 6 io_out[17]
port 200 nsew signal output
rlabel metal2 s 19706 39200 19762 40000 6 io_out[18]
port 201 nsew signal output
rlabel metal2 s 20810 39200 20866 40000 6 io_out[19]
port 202 nsew signal output
rlabel metal2 s 1858 39200 1914 40000 6 io_out[1]
port 203 nsew signal output
rlabel metal2 s 21822 39200 21878 40000 6 io_out[20]
port 204 nsew signal output
rlabel metal2 s 22926 39200 22982 40000 6 io_out[21]
port 205 nsew signal output
rlabel metal2 s 23938 39200 23994 40000 6 io_out[22]
port 206 nsew signal output
rlabel metal2 s 24950 39200 25006 40000 6 io_out[23]
port 207 nsew signal output
rlabel metal2 s 26054 39200 26110 40000 6 io_out[24]
port 208 nsew signal output
rlabel metal2 s 27066 39200 27122 40000 6 io_out[25]
port 209 nsew signal output
rlabel metal2 s 28170 39200 28226 40000 6 io_out[26]
port 210 nsew signal output
rlabel metal2 s 29182 39200 29238 40000 6 io_out[27]
port 211 nsew signal output
rlabel metal2 s 30286 39200 30342 40000 6 io_out[28]
port 212 nsew signal output
rlabel metal2 s 31298 39200 31354 40000 6 io_out[29]
port 213 nsew signal output
rlabel metal2 s 2870 39200 2926 40000 6 io_out[2]
port 214 nsew signal output
rlabel metal2 s 32402 39200 32458 40000 6 io_out[30]
port 215 nsew signal output
rlabel metal2 s 33414 39200 33470 40000 6 io_out[31]
port 216 nsew signal output
rlabel metal2 s 34426 39200 34482 40000 6 io_out[32]
port 217 nsew signal output
rlabel metal2 s 35530 39200 35586 40000 6 io_out[33]
port 218 nsew signal output
rlabel metal2 s 36542 39200 36598 40000 6 io_out[34]
port 219 nsew signal output
rlabel metal2 s 37646 39200 37702 40000 6 io_out[35]
port 220 nsew signal output
rlabel metal2 s 38658 39200 38714 40000 6 io_out[36]
port 221 nsew signal output
rlabel metal2 s 39762 39200 39818 40000 6 io_out[37]
port 222 nsew signal output
rlabel metal2 s 3882 39200 3938 40000 6 io_out[3]
port 223 nsew signal output
rlabel metal2 s 4986 39200 5042 40000 6 io_out[4]
port 224 nsew signal output
rlabel metal2 s 5998 39200 6054 40000 6 io_out[5]
port 225 nsew signal output
rlabel metal2 s 7102 39200 7158 40000 6 io_out[6]
port 226 nsew signal output
rlabel metal2 s 8114 39200 8170 40000 6 io_out[7]
port 227 nsew signal output
rlabel metal2 s 9218 39200 9274 40000 6 io_out[8]
port 228 nsew signal output
rlabel metal2 s 10230 39200 10286 40000 6 io_out[9]
port 229 nsew signal output
rlabel metal3 s 39200 37408 40000 37528 6 la_blink[0]
port 230 nsew signal output
rlabel metal3 s 39200 39040 40000 39160 6 la_blink[1]
port 231 nsew signal output
rlabel metal2 s 110 0 166 800 6 pwm_en[0]
port 232 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 pwm_en[10]
port 233 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 pwm_en[11]
port 234 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 pwm_en[12]
port 235 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 pwm_en[13]
port 236 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 pwm_en[14]
port 237 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 pwm_en[15]
port 238 nsew signal input
rlabel metal2 s 570 0 626 800 6 pwm_en[1]
port 239 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 pwm_en[2]
port 240 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 pwm_en[3]
port 241 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 pwm_en[4]
port 242 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 pwm_en[5]
port 243 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 pwm_en[6]
port 244 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 pwm_en[7]
port 245 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 pwm_en[8]
port 246 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 pwm_en[9]
port 247 nsew signal input
rlabel metal2 s 294 0 350 800 6 pwm_out[0]
port 248 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 pwm_out[10]
port 249 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 pwm_out[11]
port 250 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 pwm_out[12]
port 251 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 pwm_out[13]
port 252 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 pwm_out[14]
port 253 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 pwm_out[15]
port 254 nsew signal input
rlabel metal2 s 846 0 902 800 6 pwm_out[1]
port 255 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 pwm_out[2]
port 256 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 pwm_out[3]
port 257 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 pwm_out[4]
port 258 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 pwm_out[5]
port 259 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 pwm_out[6]
port 260 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 pwm_out[7]
port 261 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 pwm_out[8]
port 262 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 pwm_out[9]
port 263 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 rst
port 264 nsew signal input
rlabel metal3 s 39200 20816 40000 20936 6 spi_clk[0]
port 265 nsew signal input
rlabel metal3 s 39200 29112 40000 29232 6 spi_clk[1]
port 266 nsew signal input
rlabel metal3 s 39200 22448 40000 22568 6 spi_cs[0]
port 267 nsew signal input
rlabel metal3 s 39200 30744 40000 30864 6 spi_cs[1]
port 268 nsew signal input
rlabel metal3 s 39200 24080 40000 24200 6 spi_en[0]
port 269 nsew signal input
rlabel metal3 s 39200 32376 40000 32496 6 spi_en[1]
port 270 nsew signal input
rlabel metal3 s 39200 25712 40000 25832 6 spi_miso[0]
port 271 nsew signal output
rlabel metal3 s 39200 34144 40000 34264 6 spi_miso[1]
port 272 nsew signal output
rlabel metal3 s 39200 27480 40000 27600 6 spi_mosi[0]
port 273 nsew signal input
rlabel metal3 s 39200 35776 40000 35896 6 spi_mosi[1]
port 274 nsew signal input
rlabel metal3 s 39200 824 40000 944 6 uart_en[0]
port 275 nsew signal input
rlabel metal3 s 39200 5720 40000 5840 6 uart_en[1]
port 276 nsew signal input
rlabel metal3 s 39200 10752 40000 10872 6 uart_en[2]
port 277 nsew signal input
rlabel metal3 s 39200 15784 40000 15904 6 uart_en[3]
port 278 nsew signal input
rlabel metal3 s 39200 2456 40000 2576 6 uart_rx[0]
port 279 nsew signal output
rlabel metal3 s 39200 7488 40000 7608 6 uart_rx[1]
port 280 nsew signal output
rlabel metal3 s 39200 12384 40000 12504 6 uart_rx[2]
port 281 nsew signal output
rlabel metal3 s 39200 17416 40000 17536 6 uart_rx[3]
port 282 nsew signal output
rlabel metal3 s 39200 4088 40000 4208 6 uart_tx[0]
port 283 nsew signal input
rlabel metal3 s 39200 9120 40000 9240 6 uart_tx[1]
port 284 nsew signal input
rlabel metal3 s 39200 14152 40000 14272 6 uart_tx[2]
port 285 nsew signal input
rlabel metal3 s 39200 19048 40000 19168 6 uart_tx[3]
port 286 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 287 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 287 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 288 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2019436
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_IOMultiplexer/runs/Peripheral_IOMultiplexer/results/finishing/IOMultiplexer.magic.gds
string GDS_START 216428
<< end >>

