magic
tech sky130A
magscale 1 2
timestamp 1651272265
<< viali >>
rect 2145 37417 2179 37451
rect 4261 37417 4295 37451
rect 7113 37417 7147 37451
rect 12265 37417 12299 37451
rect 9689 37349 9723 37383
rect 13185 37349 13219 37383
rect 15945 37349 15979 37383
rect 18429 37349 18463 37383
rect 2973 37281 3007 37315
rect 4905 37281 4939 37315
rect 15485 37281 15519 37315
rect 17049 37281 17083 37315
rect 22201 37281 22235 37315
rect 23673 37281 23707 37315
rect 30665 37281 30699 37315
rect 32505 37281 32539 37315
rect 33977 37281 34011 37315
rect 38025 37281 38059 37315
rect 1869 37213 1903 37247
rect 2789 37213 2823 37247
rect 5089 37213 5123 37247
rect 5825 37213 5859 37247
rect 6837 37213 6871 37247
rect 7665 37213 7699 37247
rect 9413 37213 9447 37247
rect 10241 37213 10275 37247
rect 11989 37213 12023 37247
rect 14565 37213 14599 37247
rect 15301 37213 15335 37247
rect 17233 37213 17267 37247
rect 18153 37213 18187 37247
rect 19257 37213 19291 37247
rect 20177 37213 20211 37247
rect 20913 37213 20947 37247
rect 22385 37213 22419 37247
rect 22937 37213 22971 37247
rect 24409 37213 24443 37247
rect 25421 37213 25455 37247
rect 26157 37213 26191 37247
rect 26985 37213 27019 37247
rect 27905 37213 27939 37247
rect 28825 37213 28859 37247
rect 29561 37213 29595 37247
rect 30849 37213 30883 37247
rect 31585 37213 31619 37247
rect 32689 37213 32723 37247
rect 33517 37213 33551 37247
rect 34989 37213 35023 37247
rect 35725 37213 35759 37247
rect 36461 37213 36495 37247
rect 37289 37213 37323 37247
rect 4353 37145 4387 37179
rect 12909 37145 12943 37179
rect 5641 37077 5675 37111
rect 7849 37077 7883 37111
rect 10425 37077 10459 37111
rect 14657 37077 14691 37111
rect 19441 37077 19475 37111
rect 20361 37077 20395 37111
rect 21097 37077 21131 37111
rect 23121 37077 23155 37111
rect 24593 37077 24627 37111
rect 25605 37077 25639 37111
rect 26341 37077 26375 37111
rect 27169 37077 27203 37111
rect 28089 37077 28123 37111
rect 28733 37077 28767 37111
rect 29745 37077 29779 37111
rect 31401 37077 31435 37111
rect 33333 37077 33367 37111
rect 34805 37077 34839 37111
rect 35541 37077 35575 37111
rect 36277 37077 36311 37111
rect 37473 37077 37507 37111
rect 3433 36873 3467 36907
rect 4077 36873 4111 36907
rect 4813 36873 4847 36907
rect 5641 36873 5675 36907
rect 7297 36873 7331 36907
rect 8769 36873 8803 36907
rect 9413 36873 9447 36907
rect 10885 36873 10919 36907
rect 12173 36873 12207 36907
rect 13645 36873 13679 36907
rect 14473 36873 14507 36907
rect 15761 36873 15795 36907
rect 17877 36873 17911 36907
rect 18613 36873 18647 36907
rect 19533 36873 19567 36907
rect 20269 36873 20303 36907
rect 21097 36873 21131 36907
rect 22017 36873 22051 36907
rect 22753 36873 22787 36907
rect 24225 36873 24259 36907
rect 24961 36873 24995 36907
rect 25697 36873 25731 36907
rect 27905 36873 27939 36907
rect 28549 36873 28583 36907
rect 29469 36873 29503 36907
rect 30205 36873 30239 36907
rect 31217 36873 31251 36907
rect 32321 36873 32355 36907
rect 33333 36873 33367 36907
rect 34437 36873 34471 36907
rect 35449 36873 35483 36907
rect 36553 36873 36587 36907
rect 1869 36805 1903 36839
rect 10057 36805 10091 36839
rect 12909 36805 12943 36839
rect 15025 36805 15059 36839
rect 17141 36805 17175 36839
rect 37289 36805 37323 36839
rect 37933 36805 37967 36839
rect 2789 36737 2823 36771
rect 3249 36737 3283 36771
rect 4261 36737 4295 36771
rect 4997 36737 5031 36771
rect 5457 36737 5491 36771
rect 6469 36737 6503 36771
rect 7113 36737 7147 36771
rect 8125 36737 8159 36771
rect 8585 36737 8619 36771
rect 9597 36737 9631 36771
rect 10701 36737 10735 36771
rect 12357 36737 12391 36771
rect 13829 36737 13863 36771
rect 14289 36737 14323 36771
rect 15945 36737 15979 36771
rect 18061 36737 18095 36771
rect 18797 36737 18831 36771
rect 19717 36737 19751 36771
rect 20453 36737 20487 36771
rect 20913 36737 20947 36771
rect 21833 36737 21867 36771
rect 22569 36737 22603 36771
rect 23581 36737 23615 36771
rect 24041 36737 24075 36771
rect 24777 36737 24811 36771
rect 25513 36737 25547 36771
rect 26433 36737 26467 36771
rect 26985 36737 27019 36771
rect 27721 36737 27755 36771
rect 28733 36737 28767 36771
rect 29285 36737 29319 36771
rect 30021 36737 30055 36771
rect 31033 36737 31067 36771
rect 32137 36737 32171 36771
rect 33149 36737 33183 36771
rect 34253 36737 34287 36771
rect 35265 36737 35299 36771
rect 36369 36737 36403 36771
rect 11529 36669 11563 36703
rect 2053 36601 2087 36635
rect 6653 36601 6687 36635
rect 7941 36601 7975 36635
rect 13093 36601 13127 36635
rect 17325 36601 17359 36635
rect 27169 36601 27203 36635
rect 38117 36601 38151 36635
rect 2605 36533 2639 36567
rect 23397 36533 23431 36567
rect 26249 36533 26283 36567
rect 1501 36329 1535 36363
rect 2237 36329 2271 36363
rect 3065 36329 3099 36363
rect 4077 36329 4111 36363
rect 5365 36329 5399 36363
rect 6193 36329 6227 36363
rect 7297 36329 7331 36363
rect 7941 36329 7975 36363
rect 9045 36329 9079 36363
rect 10057 36329 10091 36363
rect 10793 36329 10827 36363
rect 11529 36329 11563 36363
rect 12541 36329 12575 36363
rect 14289 36329 14323 36363
rect 15209 36329 15243 36363
rect 15945 36329 15979 36363
rect 16773 36329 16807 36363
rect 17785 36329 17819 36363
rect 19349 36329 19383 36363
rect 20177 36329 20211 36363
rect 20821 36329 20855 36363
rect 21741 36329 21775 36363
rect 24501 36329 24535 36363
rect 25329 36329 25363 36363
rect 26617 36329 26651 36363
rect 27261 36329 27295 36363
rect 28641 36329 28675 36363
rect 29561 36329 29595 36363
rect 31861 36329 31895 36363
rect 34897 36329 34931 36363
rect 35449 36329 35483 36363
rect 13553 36261 13587 36295
rect 18429 36261 18463 36295
rect 22753 36261 22787 36295
rect 23673 36261 23707 36295
rect 25973 36261 26007 36295
rect 28181 36261 28215 36295
rect 32413 36261 32447 36295
rect 30941 36193 30975 36227
rect 36553 36193 36587 36227
rect 37565 36193 37599 36227
rect 1685 36125 1719 36159
rect 2421 36125 2455 36159
rect 3249 36125 3283 36159
rect 4261 36125 4295 36159
rect 5549 36125 5583 36159
rect 6377 36125 6411 36159
rect 7481 36125 7515 36159
rect 8125 36125 8159 36159
rect 9229 36125 9263 36159
rect 10241 36125 10275 36159
rect 10977 36125 11011 36159
rect 11713 36125 11747 36159
rect 12725 36125 12759 36159
rect 13369 36125 13403 36159
rect 14105 36125 14139 36159
rect 15025 36125 15059 36159
rect 16129 36125 16163 36159
rect 16957 36125 16991 36159
rect 17969 36125 18003 36159
rect 19533 36125 19567 36159
rect 19993 36125 20027 36159
rect 20637 36125 20671 36159
rect 21925 36125 21959 36159
rect 24685 36125 24719 36159
rect 26433 36125 26467 36159
rect 27077 36125 27111 36159
rect 27997 36125 28031 36159
rect 28825 36125 28859 36159
rect 30205 36125 30239 36159
rect 31677 36125 31711 36159
rect 34713 36125 34747 36159
rect 36829 36125 36863 36159
rect 37289 36125 37323 36159
rect 4905 36057 4939 36091
rect 22385 36057 22419 36091
rect 23305 36057 23339 36091
rect 30389 36057 30423 36091
rect 31125 36057 31159 36091
rect 32597 36057 32631 36091
rect 33517 36057 33551 36091
rect 34069 36057 34103 36091
rect 22845 35989 22879 36023
rect 23765 35989 23799 36023
rect 33425 35989 33459 36023
rect 1501 35785 1535 35819
rect 2697 35785 2731 35819
rect 3341 35785 3375 35819
rect 4537 35785 4571 35819
rect 5089 35785 5123 35819
rect 6653 35785 6687 35819
rect 8585 35785 8619 35819
rect 9781 35785 9815 35819
rect 10793 35785 10827 35819
rect 12265 35785 12299 35819
rect 14197 35785 14231 35819
rect 14841 35785 14875 35819
rect 15669 35785 15703 35819
rect 16681 35785 16715 35819
rect 19717 35785 19751 35819
rect 22477 35785 22511 35819
rect 23213 35785 23247 35819
rect 23765 35785 23799 35819
rect 24317 35785 24351 35819
rect 26433 35785 26467 35819
rect 30481 35785 30515 35819
rect 31217 35785 31251 35819
rect 34253 35785 34287 35819
rect 35817 35785 35851 35819
rect 37289 35785 37323 35819
rect 29929 35717 29963 35751
rect 1685 35649 1719 35683
rect 2881 35649 2915 35683
rect 3525 35649 3559 35683
rect 3985 35649 4019 35683
rect 6469 35649 6503 35683
rect 8769 35649 8803 35683
rect 9965 35649 9999 35683
rect 10977 35649 11011 35683
rect 11529 35649 11563 35683
rect 12449 35649 12483 35683
rect 14381 35649 14415 35683
rect 15025 35649 15059 35683
rect 15853 35649 15887 35683
rect 16865 35649 16899 35683
rect 17509 35649 17543 35683
rect 19533 35649 19567 35683
rect 23029 35649 23063 35683
rect 26249 35649 26283 35683
rect 27537 35649 27571 35683
rect 28365 35649 28399 35683
rect 28825 35649 28859 35683
rect 30665 35649 30699 35683
rect 32781 35649 32815 35683
rect 33609 35649 33643 35683
rect 34069 35649 34103 35683
rect 35173 35649 35207 35683
rect 35633 35649 35667 35683
rect 36461 35649 36495 35683
rect 38025 35649 38059 35683
rect 2237 35581 2271 35615
rect 18981 35581 19015 35615
rect 11713 35513 11747 35547
rect 13001 35513 13035 35547
rect 17325 35513 17359 35547
rect 27721 35513 27755 35547
rect 33425 35513 33459 35547
rect 34989 35513 35023 35547
rect 36645 35513 36679 35547
rect 37841 35513 37875 35547
rect 5733 35445 5767 35479
rect 7205 35445 7239 35479
rect 8125 35445 8159 35479
rect 13461 35445 13495 35479
rect 17969 35445 18003 35479
rect 20177 35445 20211 35479
rect 20729 35445 20763 35479
rect 22017 35445 22051 35479
rect 24869 35445 24903 35479
rect 25421 35445 25455 35479
rect 26985 35445 27019 35479
rect 28181 35445 28215 35479
rect 32689 35445 32723 35479
rect 1593 35241 1627 35275
rect 2145 35241 2179 35275
rect 6193 35241 6227 35275
rect 6745 35241 6779 35275
rect 7849 35241 7883 35275
rect 9965 35241 9999 35275
rect 10425 35241 10459 35275
rect 12173 35241 12207 35275
rect 12725 35241 12759 35275
rect 17509 35241 17543 35275
rect 18061 35241 18095 35275
rect 18613 35241 18647 35275
rect 19349 35241 19383 35275
rect 20085 35241 20119 35275
rect 29561 35241 29595 35275
rect 33517 35241 33551 35275
rect 35357 35241 35391 35275
rect 38025 35241 38059 35275
rect 2697 35173 2731 35207
rect 15301 35173 15335 35207
rect 20545 35173 20579 35207
rect 26341 35173 26375 35207
rect 34713 35173 34747 35207
rect 13369 35105 13403 35139
rect 30113 35105 30147 35139
rect 2881 35037 2915 35071
rect 10609 35037 10643 35071
rect 15117 35037 15151 35071
rect 15761 35037 15795 35071
rect 16405 35037 16439 35071
rect 31401 35037 31435 35071
rect 35541 35037 35575 35071
rect 36001 35037 36035 35071
rect 37841 35037 37875 35071
rect 11161 34969 11195 35003
rect 25973 34969 26007 35003
rect 30021 34969 30055 35003
rect 36268 34969 36302 35003
rect 3893 34901 3927 34935
rect 4445 34901 4479 34935
rect 4905 34901 4939 34935
rect 5549 34901 5583 34935
rect 7297 34901 7331 34935
rect 9045 34901 9079 34935
rect 11621 34901 11655 34935
rect 14473 34901 14507 34935
rect 15945 34901 15979 34935
rect 16957 34901 16991 34935
rect 21097 34901 21131 34935
rect 22845 34901 22879 34935
rect 26433 34901 26467 34935
rect 29009 34901 29043 34935
rect 29929 34901 29963 34935
rect 30849 34901 30883 34935
rect 31953 34901 31987 34935
rect 32965 34901 32999 34935
rect 34069 34901 34103 34935
rect 37381 34901 37415 34935
rect 2605 34697 2639 34731
rect 12081 34697 12115 34731
rect 12909 34697 12943 34731
rect 15669 34697 15703 34731
rect 16957 34697 16991 34731
rect 23305 34697 23339 34731
rect 24225 34697 24259 34731
rect 36553 34697 36587 34731
rect 37381 34697 37415 34731
rect 6377 34629 6411 34663
rect 34805 34629 34839 34663
rect 3617 34561 3651 34595
rect 4445 34561 4479 34595
rect 4712 34561 4746 34595
rect 9229 34561 9263 34595
rect 13921 34561 13955 34595
rect 14565 34561 14599 34595
rect 15117 34561 15151 34595
rect 18328 34561 18362 34595
rect 22845 34561 22879 34595
rect 23765 34561 23799 34595
rect 36737 34561 36771 34595
rect 37841 34561 37875 34595
rect 3065 34493 3099 34527
rect 9781 34493 9815 34527
rect 10793 34493 10827 34527
rect 11529 34493 11563 34527
rect 17601 34493 17635 34527
rect 18061 34493 18095 34527
rect 19993 34493 20027 34527
rect 20453 34493 20487 34527
rect 32965 34493 32999 34527
rect 33701 34493 33735 34527
rect 35265 34493 35299 34527
rect 23121 34425 23155 34459
rect 24041 34425 24075 34459
rect 38025 34425 38059 34459
rect 5825 34357 5859 34391
rect 19441 34357 19475 34391
rect 22293 34357 22327 34391
rect 36001 34357 36035 34391
rect 18061 34153 18095 34187
rect 31309 34153 31343 34187
rect 36369 34153 36403 34187
rect 37197 34153 37231 34187
rect 37933 34153 37967 34187
rect 35909 34085 35943 34119
rect 35265 34017 35299 34051
rect 9413 33949 9447 33983
rect 31493 33949 31527 33983
rect 34713 33949 34747 33983
rect 36553 33949 36587 33983
rect 37013 33949 37047 33983
rect 37749 33949 37783 33983
rect 9680 33881 9714 33915
rect 10793 33813 10827 33847
rect 11345 33813 11379 33847
rect 16037 33813 16071 33847
rect 17141 33813 17175 33847
rect 23581 33813 23615 33847
rect 33885 33813 33919 33847
rect 5273 33609 5307 33643
rect 10149 33609 10183 33643
rect 11621 33609 11655 33643
rect 18429 33609 18463 33643
rect 29377 33609 29411 33643
rect 36645 33609 36679 33643
rect 37381 33609 37415 33643
rect 38025 33609 38059 33643
rect 5457 33473 5491 33507
rect 10333 33473 10367 33507
rect 10609 33473 10643 33507
rect 11529 33473 11563 33507
rect 11805 33473 11839 33507
rect 18613 33473 18647 33507
rect 27537 33473 27571 33507
rect 29193 33473 29227 33507
rect 37841 33473 37875 33507
rect 5733 33405 5767 33439
rect 10517 33405 10551 33439
rect 18889 33405 18923 33439
rect 27813 33405 27847 33439
rect 11805 33337 11839 33371
rect 12357 33337 12391 33371
rect 5641 33269 5675 33303
rect 18797 33269 18831 33303
rect 35265 33269 35299 33303
rect 36185 33269 36219 33303
rect 19533 33065 19567 33099
rect 28457 32997 28491 33031
rect 36737 32929 36771 32963
rect 19257 32861 19291 32895
rect 19533 32861 19567 32895
rect 19993 32861 20027 32895
rect 28273 32861 28307 32895
rect 37841 32861 37875 32895
rect 38117 32861 38151 32895
rect 19349 32725 19383 32759
rect 36277 32725 36311 32759
rect 26157 32521 26191 32555
rect 32137 32521 32171 32555
rect 38117 32453 38151 32487
rect 6745 32385 6779 32419
rect 6929 32385 6963 32419
rect 13645 32385 13679 32419
rect 14105 32385 14139 32419
rect 14372 32385 14406 32419
rect 25789 32385 25823 32419
rect 25973 32385 26007 32419
rect 32505 32385 32539 32419
rect 32597 32385 32631 32419
rect 32781 32317 32815 32351
rect 6929 32249 6963 32283
rect 7481 32181 7515 32215
rect 15485 32181 15519 32215
rect 25329 32181 25363 32215
rect 31493 32181 31527 32215
rect 37565 32181 37599 32215
rect 26525 31977 26559 32011
rect 28365 31977 28399 32011
rect 27445 31841 27479 31875
rect 25605 31773 25639 31807
rect 26157 31773 26191 31807
rect 26341 31773 26375 31807
rect 27997 31773 28031 31807
rect 28181 31773 28215 31807
rect 34897 31433 34931 31467
rect 37933 31433 37967 31467
rect 34713 31297 34747 31331
rect 36470 31297 36504 31331
rect 36737 31297 36771 31331
rect 37473 31297 37507 31331
rect 38117 31297 38151 31331
rect 35357 31093 35391 31127
rect 27077 30889 27111 30923
rect 33057 30889 33091 30923
rect 35265 30889 35299 30923
rect 32873 30821 32907 30855
rect 27629 30753 27663 30787
rect 1869 30685 1903 30719
rect 3801 30685 3835 30719
rect 4813 30685 4847 30719
rect 4997 30685 5031 30719
rect 23673 30685 23707 30719
rect 2136 30617 2170 30651
rect 23406 30617 23440 30651
rect 24501 30617 24535 30651
rect 32597 30617 32631 30651
rect 3249 30549 3283 30583
rect 4905 30549 4939 30583
rect 5549 30549 5583 30583
rect 22293 30549 22327 30583
rect 26617 30549 26651 30583
rect 27445 30549 27479 30583
rect 27537 30549 27571 30583
rect 4997 30345 5031 30379
rect 12909 30345 12943 30379
rect 22753 30345 22787 30379
rect 32321 30345 32355 30379
rect 32781 30345 32815 30379
rect 3617 30277 3651 30311
rect 5165 30277 5199 30311
rect 5365 30277 5399 30311
rect 6377 30277 6411 30311
rect 6745 30277 6779 30311
rect 8033 30277 8067 30311
rect 11529 30277 11563 30311
rect 13001 30277 13035 30311
rect 14381 30277 14415 30311
rect 15485 30277 15519 30311
rect 19149 30277 19183 30311
rect 19349 30277 19383 30311
rect 20085 30277 20119 30311
rect 20177 30277 20211 30311
rect 11759 30243 11793 30277
rect 1869 30209 1903 30243
rect 3801 30209 3835 30243
rect 6561 30209 6595 30243
rect 6653 30209 6687 30243
rect 6929 30209 6963 30243
rect 7849 30209 7883 30243
rect 12817 30209 12851 30243
rect 14565 30209 14599 30243
rect 15393 30209 15427 30243
rect 15577 30209 15611 30243
rect 17233 30209 17267 30243
rect 18245 30209 18279 30243
rect 18337 30209 18371 30243
rect 18521 30209 18555 30243
rect 19993 30209 20027 30243
rect 22569 30209 22603 30243
rect 32229 30209 32263 30243
rect 4077 30141 4111 30175
rect 14749 30141 14783 30175
rect 14841 30141 14875 30175
rect 17509 30141 17543 30175
rect 19809 30141 19843 30175
rect 22293 30141 22327 30175
rect 32137 30141 32171 30175
rect 32505 30141 32539 30175
rect 32597 30141 32631 30175
rect 2145 30073 2179 30107
rect 12633 30073 12667 30107
rect 18981 30073 19015 30107
rect 22385 30073 22419 30107
rect 3985 30005 4019 30039
rect 5181 30005 5215 30039
rect 11713 30005 11747 30039
rect 11897 30005 11931 30039
rect 13185 30005 13219 30039
rect 16129 30005 16163 30039
rect 18521 30005 18555 30039
rect 19165 30005 19199 30039
rect 20361 30005 20395 30039
rect 31493 30005 31527 30039
rect 1593 29801 1627 29835
rect 32689 29801 32723 29835
rect 37933 29801 37967 29835
rect 11345 29733 11379 29767
rect 32505 29665 32539 29699
rect 11069 29597 11103 29631
rect 11161 29597 11195 29631
rect 25421 29597 25455 29631
rect 32229 29597 32263 29631
rect 32321 29597 32355 29631
rect 32413 29597 32447 29631
rect 37473 29597 37507 29631
rect 38117 29597 38151 29631
rect 9873 29529 9907 29563
rect 10057 29529 10091 29563
rect 11345 29529 11379 29563
rect 25237 29529 25271 29563
rect 10517 29257 10551 29291
rect 11529 29257 11563 29291
rect 22937 29257 22971 29291
rect 8944 29189 8978 29223
rect 23489 29189 23523 29223
rect 11529 29121 11563 29155
rect 11621 29121 11655 29155
rect 22845 29121 22879 29155
rect 23029 29121 23063 29155
rect 31125 29121 31159 29155
rect 8677 29053 8711 29087
rect 11805 29053 11839 29087
rect 12265 29053 12299 29087
rect 10057 28985 10091 29019
rect 31309 28985 31343 29019
rect 6193 28713 6227 28747
rect 6929 28713 6963 28747
rect 18337 28645 18371 28679
rect 6745 28509 6779 28543
rect 18429 28509 18463 28543
rect 18153 28441 18187 28475
rect 30665 28441 30699 28475
rect 30849 28441 30883 28475
rect 17601 28373 17635 28407
rect 18429 28373 18463 28407
rect 26525 28373 26559 28407
rect 29101 28169 29135 28203
rect 32229 28101 32263 28135
rect 26157 28033 26191 28067
rect 26249 28033 26283 28067
rect 26433 28033 26467 28067
rect 27169 28033 27203 28067
rect 27436 28033 27470 28067
rect 32137 28033 32171 28067
rect 32413 28033 32447 28067
rect 37473 28033 37507 28067
rect 38117 28033 38151 28067
rect 28549 27897 28583 27931
rect 26433 27829 26467 27863
rect 32413 27829 32447 27863
rect 37933 27829 37967 27863
rect 27353 27625 27387 27659
rect 4813 27557 4847 27591
rect 6009 27557 6043 27591
rect 18705 27557 18739 27591
rect 37565 27557 37599 27591
rect 26985 27489 27019 27523
rect 31769 27489 31803 27523
rect 31953 27489 31987 27523
rect 35725 27489 35759 27523
rect 36185 27489 36219 27523
rect 4537 27421 4571 27455
rect 4629 27421 4663 27455
rect 5273 27421 5307 27455
rect 5457 27421 5491 27455
rect 17325 27421 17359 27455
rect 17592 27421 17626 27455
rect 26893 27421 26927 27455
rect 27169 27421 27203 27455
rect 31493 27421 31527 27455
rect 31585 27421 31619 27455
rect 31677 27421 31711 27455
rect 32413 27421 32447 27455
rect 32597 27421 32631 27455
rect 32505 27353 32539 27387
rect 36430 27353 36464 27387
rect 5365 27285 5399 27319
rect 16773 27285 16807 27319
rect 30849 27285 30883 27319
rect 34345 27081 34379 27115
rect 33885 27013 33919 27047
rect 15025 26945 15059 26979
rect 35458 26945 35492 26979
rect 35725 26945 35759 26979
rect 15209 26741 15243 26775
rect 15853 26741 15887 26775
rect 4169 26469 4203 26503
rect 3985 26333 4019 26367
rect 4261 26333 4295 26367
rect 3801 26197 3835 26231
rect 3709 25993 3743 26027
rect 27077 25993 27111 26027
rect 30849 25993 30883 26027
rect 4169 25925 4203 25959
rect 8401 25925 8435 25959
rect 23765 25925 23799 25959
rect 30205 25925 30239 25959
rect 30757 25925 30791 25959
rect 2329 25857 2363 25891
rect 2596 25857 2630 25891
rect 21833 25857 21867 25891
rect 22100 25857 22134 25891
rect 26433 25857 26467 25891
rect 27261 25857 27295 25891
rect 13921 25721 13955 25755
rect 38117 25721 38151 25755
rect 23213 25653 23247 25687
rect 9137 25449 9171 25483
rect 13093 25449 13127 25483
rect 22017 25449 22051 25483
rect 22385 25449 22419 25483
rect 31033 25449 31067 25483
rect 22937 25381 22971 25415
rect 6929 25313 6963 25347
rect 15485 25313 15519 25347
rect 31585 25313 31619 25347
rect 9873 25245 9907 25279
rect 10149 25245 10183 25279
rect 10333 25245 10367 25279
rect 22201 25245 22235 25279
rect 22477 25245 22511 25279
rect 23121 25245 23155 25279
rect 23213 25245 23247 25279
rect 31493 25245 31527 25279
rect 7196 25177 7230 25211
rect 15218 25177 15252 25211
rect 22937 25177 22971 25211
rect 23673 25177 23707 25211
rect 28825 25177 28859 25211
rect 29009 25177 29043 25211
rect 8309 25109 8343 25143
rect 9689 25109 9723 25143
rect 14105 25109 14139 25143
rect 28181 25109 28215 25143
rect 31401 25109 31435 25143
rect 32229 25109 32263 25143
rect 7941 24905 7975 24939
rect 13001 24905 13035 24939
rect 12633 24837 12667 24871
rect 12725 24837 12759 24871
rect 8125 24769 8159 24803
rect 9321 24769 9355 24803
rect 9505 24769 9539 24803
rect 10149 24769 10183 24803
rect 10333 24769 10367 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 12541 24769 12575 24803
rect 12909 24769 12943 24803
rect 13001 24769 13035 24803
rect 13645 24769 13679 24803
rect 9689 24701 9723 24735
rect 10977 24701 11011 24735
rect 13553 24701 13587 24735
rect 11621 24633 11655 24667
rect 20913 24361 20947 24395
rect 25697 24361 25731 24395
rect 29561 24293 29595 24327
rect 12817 24225 12851 24259
rect 12633 24157 12667 24191
rect 25053 24157 25087 24191
rect 25237 24157 25271 24191
rect 30389 24157 30423 24191
rect 30573 24157 30607 24191
rect 19625 24089 19659 24123
rect 29745 24089 29779 24123
rect 29929 24089 29963 24123
rect 30757 24089 30791 24123
rect 31217 24089 31251 24123
rect 37841 24089 37875 24123
rect 38025 24089 38059 24123
rect 12449 24021 12483 24055
rect 25145 24021 25179 24055
rect 37381 24021 37415 24055
rect 37749 23817 37783 23851
rect 31217 23749 31251 23783
rect 31401 23749 31435 23783
rect 17592 23681 17626 23715
rect 31585 23681 31619 23715
rect 37657 23681 37691 23715
rect 17325 23613 17359 23647
rect 37841 23613 37875 23647
rect 18705 23545 18739 23579
rect 37289 23545 37323 23579
rect 16773 23477 16807 23511
rect 19441 23477 19475 23511
rect 30021 23477 30055 23511
rect 32137 23477 32171 23511
rect 17233 23273 17267 23307
rect 18061 23273 18095 23307
rect 21005 23205 21039 23239
rect 17785 23137 17819 23171
rect 32505 23137 32539 23171
rect 17969 23069 18003 23103
rect 18061 23069 18095 23103
rect 21281 23069 21315 23103
rect 25789 23069 25823 23103
rect 27629 23069 27663 23103
rect 32229 23069 32263 23103
rect 38025 23069 38059 23103
rect 21005 23001 21039 23035
rect 26056 23001 26090 23035
rect 21189 22933 21223 22967
rect 27169 22933 27203 22967
rect 37565 22933 37599 22967
rect 25973 22729 26007 22763
rect 33241 22729 33275 22763
rect 33701 22729 33735 22763
rect 37749 22729 37783 22763
rect 35081 22661 35115 22695
rect 35633 22661 35667 22695
rect 22017 22593 22051 22627
rect 22109 22593 22143 22627
rect 26157 22593 26191 22627
rect 33609 22593 33643 22627
rect 37841 22593 37875 22627
rect 26433 22525 26467 22559
rect 33793 22525 33827 22559
rect 35909 22457 35943 22491
rect 21833 22389 21867 22423
rect 26341 22389 26375 22423
rect 32781 22389 32815 22423
rect 36093 22389 36127 22423
rect 20821 22049 20855 22083
rect 21189 22049 21223 22083
rect 31217 22049 31251 22083
rect 4629 21981 4663 22015
rect 21005 21981 21039 22015
rect 37473 21981 37507 22015
rect 38117 21981 38151 22015
rect 4896 21913 4930 21947
rect 30941 21913 30975 21947
rect 6009 21845 6043 21879
rect 6561 21845 6595 21879
rect 30021 21845 30055 21879
rect 30573 21845 30607 21879
rect 31033 21845 31067 21879
rect 37933 21845 37967 21879
rect 2053 21505 2087 21539
rect 2320 21505 2354 21539
rect 23397 21505 23431 21539
rect 23581 21505 23615 21539
rect 3433 21301 3467 21335
rect 3985 21301 4019 21335
rect 6377 21097 6411 21131
rect 6561 20961 6595 20995
rect 6653 20961 6687 20995
rect 7297 20961 7331 20995
rect 37013 20961 37047 20995
rect 6745 20893 6779 20927
rect 10977 20893 11011 20927
rect 37289 20893 37323 20927
rect 11222 20825 11256 20859
rect 10425 20757 10459 20791
rect 12357 20757 12391 20791
rect 6561 20553 6595 20587
rect 6745 20553 6779 20587
rect 10149 20553 10183 20587
rect 37933 20553 37967 20587
rect 6929 20485 6963 20519
rect 28273 20485 28307 20519
rect 28457 20485 28491 20519
rect 6837 20417 6871 20451
rect 10425 20417 10459 20451
rect 11529 20417 11563 20451
rect 15209 20417 15243 20451
rect 15945 20417 15979 20451
rect 37473 20417 37507 20451
rect 38117 20417 38151 20451
rect 7113 20349 7147 20383
rect 10333 20349 10367 20383
rect 10517 20349 10551 20383
rect 15393 20281 15427 20315
rect 6837 20009 6871 20043
rect 18153 20009 18187 20043
rect 26709 20009 26743 20043
rect 4169 19941 4203 19975
rect 13093 19941 13127 19975
rect 17325 19941 17359 19975
rect 23029 19941 23063 19975
rect 27261 19941 27295 19975
rect 7205 19873 7239 19907
rect 7297 19873 7331 19907
rect 18245 19873 18279 19907
rect 30389 19873 30423 19907
rect 4353 19805 4387 19839
rect 7021 19805 7055 19839
rect 7113 19805 7147 19839
rect 10149 19805 10183 19839
rect 12725 19805 12759 19839
rect 15945 19805 15979 19839
rect 17969 19805 18003 19839
rect 22477 19805 22511 19839
rect 23029 19805 23063 19839
rect 23305 19805 23339 19839
rect 26893 19805 26927 19839
rect 30113 19805 30147 19839
rect 30849 19805 30883 19839
rect 31033 19805 31067 19839
rect 31493 19805 31527 19839
rect 9965 19737 9999 19771
rect 12909 19737 12943 19771
rect 16212 19737 16246 19771
rect 17785 19737 17819 19771
rect 27077 19737 27111 19771
rect 12541 19669 12575 19703
rect 12817 19669 12851 19703
rect 15485 19669 15519 19703
rect 23213 19669 23247 19703
rect 26985 19669 27019 19703
rect 30941 19669 30975 19703
rect 12265 19465 12299 19499
rect 19993 19465 20027 19499
rect 26249 19465 26283 19499
rect 30205 19465 30239 19499
rect 33425 19465 33459 19499
rect 34345 19465 34379 19499
rect 36277 19465 36311 19499
rect 19901 19397 19935 19431
rect 27137 19397 27171 19431
rect 27353 19397 27387 19431
rect 37473 19397 37507 19431
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 19625 19329 19659 19363
rect 19809 19329 19843 19363
rect 26157 19329 26191 19363
rect 26433 19329 26467 19363
rect 31318 19329 31352 19363
rect 31585 19329 31619 19363
rect 34161 19329 34195 19363
rect 34437 19329 34471 19363
rect 34897 19329 34931 19363
rect 35153 19329 35187 19363
rect 37657 19329 37691 19363
rect 12541 19261 12575 19295
rect 12633 19261 12667 19295
rect 29653 19261 29687 19295
rect 33977 19261 34011 19295
rect 37289 19261 37323 19295
rect 20177 19193 20211 19227
rect 26433 19125 26467 19159
rect 26985 19125 27019 19159
rect 27169 19125 27203 19159
rect 19809 18921 19843 18955
rect 23121 18921 23155 18955
rect 34713 18921 34747 18955
rect 26341 18853 26375 18887
rect 25789 18785 25823 18819
rect 26525 18785 26559 18819
rect 23029 18717 23063 18751
rect 23305 18717 23339 18751
rect 26249 18717 26283 18751
rect 37473 18717 37507 18751
rect 38117 18717 38151 18751
rect 19793 18649 19827 18683
rect 19993 18649 20027 18683
rect 19625 18581 19659 18615
rect 23489 18581 23523 18615
rect 26249 18581 26283 18615
rect 37933 18581 37967 18615
rect 2973 18377 3007 18411
rect 17785 18377 17819 18411
rect 3157 18241 3191 18275
rect 17693 18241 17727 18275
rect 17877 18241 17911 18275
rect 3433 18173 3467 18207
rect 3341 18037 3375 18071
rect 3249 17833 3283 17867
rect 8309 17833 8343 17867
rect 9781 17833 9815 17867
rect 22385 17833 22419 17867
rect 4169 17697 4203 17731
rect 3065 17629 3099 17663
rect 3249 17629 3283 17663
rect 3985 17629 4019 17663
rect 8217 17629 8251 17663
rect 8953 17629 8987 17663
rect 23498 17629 23532 17663
rect 23765 17629 23799 17663
rect 38117 17629 38151 17663
rect 3801 17493 3835 17527
rect 9137 17493 9171 17527
rect 24501 17493 24535 17527
rect 8493 17289 8527 17323
rect 13001 17289 13035 17323
rect 7665 17153 7699 17187
rect 7849 17153 7883 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 13185 17153 13219 17187
rect 33885 17153 33919 17187
rect 7573 17085 7607 17119
rect 7757 17085 7791 17119
rect 13369 17085 13403 17119
rect 34161 17085 34195 17119
rect 7389 16949 7423 16983
rect 12265 16949 12299 16983
rect 7021 16745 7055 16779
rect 12449 16745 12483 16779
rect 31677 16609 31711 16643
rect 12265 16541 12299 16575
rect 12541 16541 12575 16575
rect 17699 16541 17733 16575
rect 17877 16541 17911 16575
rect 31401 16541 31435 16575
rect 7205 16473 7239 16507
rect 6837 16405 6871 16439
rect 7005 16405 7039 16439
rect 12081 16405 12115 16439
rect 17785 16405 17819 16439
rect 37473 16405 37507 16439
rect 29929 16201 29963 16235
rect 30665 16201 30699 16235
rect 33977 16201 34011 16235
rect 34437 16201 34471 16235
rect 37749 16133 37783 16167
rect 37933 16133 37967 16167
rect 4261 16065 4295 16099
rect 4445 16065 4479 16099
rect 18705 16065 18739 16099
rect 18889 16065 18923 16099
rect 18981 16065 19015 16099
rect 29837 16065 29871 16099
rect 30573 16065 30607 16099
rect 34345 16065 34379 16099
rect 34621 15997 34655 16031
rect 4445 15861 4479 15895
rect 18521 15861 18555 15895
rect 33425 15861 33459 15895
rect 4169 15657 4203 15691
rect 12449 15657 12483 15691
rect 20637 15657 20671 15691
rect 27721 15657 27755 15691
rect 30665 15657 30699 15691
rect 32505 15657 32539 15691
rect 34805 15657 34839 15691
rect 37933 15657 37967 15691
rect 27169 15589 27203 15623
rect 31677 15589 31711 15623
rect 18705 15521 18739 15555
rect 19257 15521 19291 15555
rect 25789 15521 25823 15555
rect 31953 15521 31987 15555
rect 3985 15453 4019 15487
rect 4261 15453 4295 15487
rect 10609 15453 10643 15487
rect 11069 15453 11103 15487
rect 19513 15453 19547 15487
rect 29745 15453 29779 15487
rect 30297 15453 30331 15487
rect 30481 15453 30515 15487
rect 34897 15453 34931 15487
rect 35357 15453 35391 15487
rect 36553 15453 36587 15487
rect 37197 15453 37231 15487
rect 38025 15453 38059 15487
rect 11336 15385 11370 15419
rect 26056 15385 26090 15419
rect 37013 15385 37047 15419
rect 3801 15317 3835 15351
rect 31493 15317 31527 15351
rect 7297 15113 7331 15147
rect 17141 15113 17175 15147
rect 23213 15113 23247 15147
rect 28273 15113 28307 15147
rect 29653 15113 29687 15147
rect 36645 15113 36679 15147
rect 37473 15113 37507 15147
rect 38025 15113 38059 15147
rect 22385 15045 22419 15079
rect 28733 15045 28767 15079
rect 29193 15045 29227 15079
rect 7481 14977 7515 15011
rect 17233 14977 17267 15011
rect 22569 14977 22603 15011
rect 36001 14977 36035 15011
rect 36553 14977 36587 15011
rect 37289 14977 37323 15011
rect 7665 14909 7699 14943
rect 28365 14841 28399 14875
rect 29469 14841 29503 14875
rect 14657 14773 14691 14807
rect 23765 14773 23799 14807
rect 27721 14773 27755 14807
rect 14289 14569 14323 14603
rect 15117 14569 15151 14603
rect 24409 14569 24443 14603
rect 29561 14569 29595 14603
rect 23857 14501 23891 14535
rect 15761 14433 15795 14467
rect 23121 14433 23155 14467
rect 7297 14365 7331 14399
rect 7573 14365 7607 14399
rect 7757 14365 7791 14399
rect 15025 14365 15059 14399
rect 22845 14365 22879 14399
rect 23673 14365 23707 14399
rect 36829 14365 36863 14399
rect 37289 14365 37323 14399
rect 37565 14365 37599 14399
rect 14841 14297 14875 14331
rect 7113 14229 7147 14263
rect 4077 14025 4111 14059
rect 31401 14025 31435 14059
rect 4537 13957 4571 13991
rect 14197 13957 14231 13991
rect 17049 13957 17083 13991
rect 24317 13957 24351 13991
rect 24501 13957 24535 13991
rect 25697 13957 25731 13991
rect 26249 13957 26283 13991
rect 31493 13957 31527 13991
rect 37933 13957 37967 13991
rect 2697 13889 2731 13923
rect 2964 13889 2998 13923
rect 14013 13889 14047 13923
rect 17233 13889 17267 13923
rect 23489 13889 23523 13923
rect 23765 13889 23799 13923
rect 25513 13889 25547 13923
rect 37749 13889 37783 13923
rect 14657 13821 14691 13855
rect 15117 13821 15151 13855
rect 14933 13753 14967 13787
rect 22845 13481 22879 13515
rect 24409 13481 24443 13515
rect 23489 13345 23523 13379
rect 23305 13277 23339 13311
rect 37473 13209 37507 13243
rect 14473 13141 14507 13175
rect 22293 13141 22327 13175
rect 23213 13141 23247 13175
rect 8309 12937 8343 12971
rect 25789 12937 25823 12971
rect 8769 12869 8803 12903
rect 13277 12869 13311 12903
rect 6929 12801 6963 12835
rect 7196 12801 7230 12835
rect 13093 12801 13127 12835
rect 25973 12801 26007 12835
rect 32137 12801 32171 12835
rect 33425 12801 33459 12835
rect 34069 12801 34103 12835
rect 32413 12733 32447 12767
rect 19809 12597 19843 12631
rect 23765 12597 23799 12631
rect 33609 12597 33643 12631
rect 38117 12597 38151 12631
rect 10241 12393 10275 12427
rect 19533 12393 19567 12427
rect 31125 12393 31159 12427
rect 4445 12325 4479 12359
rect 20637 12325 20671 12359
rect 21925 12325 21959 12359
rect 9505 12189 9539 12223
rect 4261 12121 4295 12155
rect 18613 12121 18647 12155
rect 19257 12121 19291 12155
rect 19441 12121 19475 12155
rect 20913 12121 20947 12155
rect 31401 12121 31435 12155
rect 9689 12053 9723 12087
rect 20453 12053 20487 12087
rect 21465 12053 21499 12087
rect 27997 12053 28031 12087
rect 2881 11849 2915 11883
rect 10333 11849 10367 11883
rect 17693 11849 17727 11883
rect 19073 11849 19107 11883
rect 30205 11849 30239 11883
rect 31125 11849 31159 11883
rect 3709 11781 3743 11815
rect 18153 11781 18187 11815
rect 18613 11781 18647 11815
rect 19533 11781 19567 11815
rect 22477 11781 22511 11815
rect 27629 11781 27663 11815
rect 28089 11781 28123 11815
rect 30665 11781 30699 11815
rect 31585 11781 31619 11815
rect 2789 11713 2823 11747
rect 3525 11713 3559 11747
rect 10149 11713 10183 11747
rect 22293 11713 22327 11747
rect 12081 11645 12115 11679
rect 12449 11577 12483 11611
rect 17785 11577 17819 11611
rect 18889 11577 18923 11611
rect 27261 11577 27295 11611
rect 28365 11577 28399 11611
rect 30389 11577 30423 11611
rect 31217 11577 31251 11611
rect 12541 11509 12575 11543
rect 13093 11509 13127 11543
rect 27169 11509 27203 11543
rect 28549 11509 28583 11543
rect 2053 11305 2087 11339
rect 12725 11305 12759 11339
rect 18337 11305 18371 11339
rect 26985 11305 27019 11339
rect 37933 11305 37967 11339
rect 28273 11237 28307 11271
rect 33333 11237 33367 11271
rect 27997 11169 28031 11203
rect 28457 11169 28491 11203
rect 2697 11101 2731 11135
rect 12817 11101 12851 11135
rect 37381 11101 37415 11135
rect 38117 11101 38151 11135
rect 2881 11033 2915 11067
rect 13001 11033 13035 11067
rect 22109 11033 22143 11067
rect 33149 11033 33183 11067
rect 27813 10761 27847 10795
rect 36001 10761 36035 10795
rect 37473 10761 37507 10795
rect 5089 10693 5123 10727
rect 4905 10625 4939 10659
rect 12173 10625 12207 10659
rect 36553 10625 36587 10659
rect 37289 10625 37323 10659
rect 12357 10421 12391 10455
rect 17509 10421 17543 10455
rect 36737 10421 36771 10455
rect 2881 10217 2915 10251
rect 15393 10217 15427 10251
rect 17693 10217 17727 10251
rect 6193 10149 6227 10183
rect 14841 10149 14875 10183
rect 17049 10149 17083 10183
rect 28457 10013 28491 10047
rect 2789 9945 2823 9979
rect 6009 9945 6043 9979
rect 14473 9945 14507 9979
rect 16221 9945 16255 9979
rect 16681 9945 16715 9979
rect 17785 9945 17819 9979
rect 17969 9945 18003 9979
rect 18521 9945 18555 9979
rect 14933 9877 14967 9911
rect 17141 9877 17175 9911
rect 28641 9877 28675 9911
rect 9781 9605 9815 9639
rect 14105 9605 14139 9639
rect 14289 9605 14323 9639
rect 17325 9605 17359 9639
rect 24409 9605 24443 9639
rect 13461 9537 13495 9571
rect 14473 9537 14507 9571
rect 24777 9537 24811 9571
rect 29009 9537 29043 9571
rect 30021 9537 30055 9571
rect 37749 9537 37783 9571
rect 24317 9469 24351 9503
rect 29193 9401 29227 9435
rect 13645 9333 13679 9367
rect 25329 9333 25363 9367
rect 30205 9333 30239 9367
rect 37841 9333 37875 9367
rect 3801 9129 3835 9163
rect 4997 9129 5031 9163
rect 5917 9129 5951 9163
rect 34805 9129 34839 9163
rect 2881 9061 2915 9095
rect 5733 9061 5767 9095
rect 9597 9061 9631 9095
rect 10517 9061 10551 9095
rect 21005 9061 21039 9095
rect 21557 9061 21591 9095
rect 25605 8993 25639 9027
rect 24501 8925 24535 8959
rect 25881 8925 25915 8959
rect 35909 8925 35943 8959
rect 36553 8925 36587 8959
rect 37473 8925 37507 8959
rect 38117 8925 38151 8959
rect 2513 8857 2547 8891
rect 5457 8857 5491 8891
rect 9229 8857 9263 8891
rect 10149 8857 10183 8891
rect 10333 8857 10367 8891
rect 20085 8857 20119 8891
rect 20637 8857 20671 8891
rect 24961 8857 24995 8891
rect 26065 8857 26099 8891
rect 35081 8857 35115 8891
rect 35357 8857 35391 8891
rect 2973 8789 3007 8823
rect 9689 8789 9723 8823
rect 21097 8789 21131 8823
rect 24685 8789 24719 8823
rect 26617 8789 26651 8823
rect 35265 8789 35299 8823
rect 36093 8789 36127 8823
rect 37933 8789 37967 8823
rect 2697 8585 2731 8619
rect 4169 8585 4203 8619
rect 23489 8585 23523 8619
rect 24869 8585 24903 8619
rect 25421 8585 25455 8619
rect 38117 8585 38151 8619
rect 4077 8517 4111 8551
rect 6377 8517 6411 8551
rect 6745 8517 6779 8551
rect 7297 8517 7331 8551
rect 12541 8517 12575 8551
rect 20913 8517 20947 8551
rect 32321 8517 32355 8551
rect 33241 8517 33275 8551
rect 33425 8517 33459 8551
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 6561 8449 6595 8483
rect 9781 8449 9815 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 20729 8449 20763 8483
rect 32689 8449 32723 8483
rect 33609 8449 33643 8483
rect 11529 8381 11563 8415
rect 24409 8381 24443 8415
rect 32229 8381 32263 8415
rect 35725 8381 35759 8415
rect 9965 8313 9999 8347
rect 11897 8313 11931 8347
rect 20085 8313 20119 8347
rect 24041 8313 24075 8347
rect 36277 8313 36311 8347
rect 37473 8313 37507 8347
rect 11989 8245 12023 8279
rect 23949 8245 23983 8279
rect 30113 8041 30147 8075
rect 37197 8041 37231 8075
rect 11805 7973 11839 8007
rect 32045 7905 32079 7939
rect 11621 7837 11655 7871
rect 24869 7837 24903 7871
rect 32413 7837 32447 7871
rect 35081 7837 35115 7871
rect 38117 7837 38151 7871
rect 11437 7769 11471 7803
rect 30021 7769 30055 7803
rect 31953 7769 31987 7803
rect 37105 7769 37139 7803
rect 3249 7701 3283 7735
rect 20453 7701 20487 7735
rect 25053 7701 25087 7735
rect 35541 7701 35575 7735
rect 36553 7701 36587 7735
rect 14749 7497 14783 7531
rect 26341 7497 26375 7531
rect 28641 7497 28675 7531
rect 7481 7429 7515 7463
rect 7849 7429 7883 7463
rect 8401 7429 8435 7463
rect 28089 7429 28123 7463
rect 37841 7429 37875 7463
rect 7665 7361 7699 7395
rect 11529 7361 11563 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 15577 7361 15611 7395
rect 26985 7361 27019 7395
rect 34069 7361 34103 7395
rect 6561 7293 6595 7327
rect 7021 7293 7055 7327
rect 14289 7293 14323 7327
rect 20361 7293 20395 7327
rect 27905 7293 27939 7327
rect 35633 7293 35667 7327
rect 6837 7225 6871 7259
rect 14565 7225 14599 7259
rect 20637 7225 20671 7259
rect 37657 7225 37691 7259
rect 11713 7157 11747 7191
rect 16129 7157 16163 7191
rect 20821 7157 20855 7191
rect 27169 7157 27203 7191
rect 34621 7157 34655 7191
rect 36093 7157 36127 7191
rect 36737 7157 36771 7191
rect 14841 6953 14875 6987
rect 16865 6885 16899 6919
rect 31769 6885 31803 6919
rect 7113 6817 7147 6851
rect 16037 6817 16071 6851
rect 20361 6817 20395 6851
rect 25053 6817 25087 6851
rect 31217 6817 31251 6851
rect 32137 6817 32171 6851
rect 19533 6749 19567 6783
rect 21005 6749 21039 6783
rect 27629 6749 27663 6783
rect 28273 6749 28307 6783
rect 35265 6749 35299 6783
rect 36645 6749 36679 6783
rect 37197 6749 37231 6783
rect 37841 6749 37875 6783
rect 16589 6681 16623 6715
rect 19993 6681 20027 6715
rect 20177 6681 20211 6715
rect 24869 6681 24903 6715
rect 5273 6613 5307 6647
rect 17049 6613 17083 6647
rect 19349 6613 19383 6647
rect 27813 6613 27847 6647
rect 29929 6613 29963 6647
rect 30573 6613 30607 6647
rect 31677 6613 31711 6647
rect 32597 6613 32631 6647
rect 33241 6613 33275 6647
rect 33793 6613 33827 6647
rect 34713 6613 34747 6647
rect 36093 6613 36127 6647
rect 37381 6613 37415 6647
rect 38025 6613 38059 6647
rect 3801 6409 3835 6443
rect 36737 6409 36771 6443
rect 4353 6341 4387 6375
rect 15577 6341 15611 6375
rect 16681 6341 16715 6375
rect 37841 6341 37875 6375
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 35265 6273 35299 6307
rect 36093 6273 36127 6307
rect 36553 6273 36587 6307
rect 3341 6205 3375 6239
rect 34805 6205 34839 6239
rect 3709 6137 3743 6171
rect 31493 6137 31527 6171
rect 35449 6137 35483 6171
rect 1501 6069 1535 6103
rect 2513 6069 2547 6103
rect 4813 6069 4847 6103
rect 5457 6069 5491 6103
rect 15025 6069 15059 6103
rect 17601 6069 17635 6103
rect 29653 6069 29687 6103
rect 30481 6069 30515 6103
rect 30941 6069 30975 6103
rect 32137 6069 32171 6103
rect 32873 6069 32907 6103
rect 33609 6069 33643 6103
rect 34161 6069 34195 6103
rect 35909 6069 35943 6103
rect 37749 6069 37783 6103
rect 3801 5865 3835 5899
rect 16221 5865 16255 5899
rect 18521 5865 18555 5899
rect 25145 5865 25179 5899
rect 26893 5865 26927 5899
rect 30021 5865 30055 5899
rect 30665 5865 30699 5899
rect 31309 5865 31343 5899
rect 33333 5865 33367 5899
rect 33977 5865 34011 5899
rect 34897 5865 34931 5899
rect 37933 5865 37967 5899
rect 36461 5797 36495 5831
rect 12541 5729 12575 5763
rect 4169 5661 4203 5695
rect 4721 5661 4755 5695
rect 25697 5661 25731 5695
rect 26341 5661 26375 5695
rect 30113 5661 30147 5695
rect 33517 5661 33551 5695
rect 34713 5661 34747 5695
rect 35449 5661 35483 5695
rect 36645 5661 36679 5695
rect 37105 5661 37139 5695
rect 2513 5593 2547 5627
rect 3985 5593 4019 5627
rect 12633 5593 12667 5627
rect 38025 5593 38059 5627
rect 1409 5525 1443 5559
rect 1961 5525 1995 5559
rect 3249 5525 3283 5559
rect 5181 5525 5215 5559
rect 5733 5525 5767 5559
rect 6377 5525 6411 5559
rect 6929 5525 6963 5559
rect 8033 5525 8067 5559
rect 9413 5525 9447 5559
rect 11069 5525 11103 5559
rect 12725 5525 12759 5559
rect 13093 5525 13127 5559
rect 14105 5525 14139 5559
rect 14657 5525 14691 5559
rect 15669 5525 15703 5559
rect 20361 5525 20395 5559
rect 21189 5525 21223 5559
rect 22109 5525 22143 5559
rect 24593 5525 24627 5559
rect 25881 5525 25915 5559
rect 29009 5525 29043 5559
rect 31953 5525 31987 5559
rect 32873 5525 32907 5559
rect 35633 5525 35667 5559
rect 37289 5525 37323 5559
rect 26341 5321 26375 5355
rect 29285 5321 29319 5355
rect 30021 5321 30055 5355
rect 32137 5321 32171 5355
rect 33057 5321 33091 5355
rect 33885 5321 33919 5355
rect 34897 5321 34931 5355
rect 37381 5321 37415 5355
rect 34805 5253 34839 5287
rect 35449 5253 35483 5287
rect 29837 5185 29871 5219
rect 31401 5185 31435 5219
rect 32321 5185 32355 5219
rect 33241 5185 33275 5219
rect 34069 5185 34103 5219
rect 35633 5185 35667 5219
rect 36461 5185 36495 5219
rect 38117 5185 38151 5219
rect 30481 5117 30515 5151
rect 4537 5049 4571 5083
rect 37933 5049 37967 5083
rect 1501 4981 1535 5015
rect 1961 4981 1995 5015
rect 2605 4981 2639 5015
rect 3157 4981 3191 5015
rect 3801 4981 3835 5015
rect 4997 4981 5031 5015
rect 5733 4981 5767 5015
rect 6469 4981 6503 5015
rect 7205 4981 7239 5015
rect 7941 4981 7975 5015
rect 8493 4981 8527 5015
rect 9045 4981 9079 5015
rect 9597 4981 9631 5015
rect 10149 4981 10183 5015
rect 10701 4981 10735 5015
rect 11713 4981 11747 5015
rect 12265 4981 12299 5015
rect 12817 4981 12851 5015
rect 13369 4981 13403 5015
rect 14013 4981 14047 5015
rect 14841 4981 14875 5015
rect 15761 4981 15795 5015
rect 16681 4981 16715 5015
rect 17233 4981 17267 5015
rect 18337 4981 18371 5015
rect 18981 4981 19015 5015
rect 19441 4981 19475 5015
rect 20453 4981 20487 5015
rect 21097 4981 21131 5015
rect 21833 4981 21867 5015
rect 22477 4981 22511 5015
rect 22937 4981 22971 5015
rect 23765 4981 23799 5015
rect 24317 4981 24351 5015
rect 25053 4981 25087 5015
rect 25789 4981 25823 5015
rect 27537 4981 27571 5015
rect 27997 4981 28031 5015
rect 28733 4981 28767 5015
rect 31585 4981 31619 5015
rect 36645 4981 36679 5015
rect 6101 4777 6135 4811
rect 8309 4777 8343 4811
rect 14105 4777 14139 4811
rect 25145 4777 25179 4811
rect 27445 4777 27479 4811
rect 30573 4777 30607 4811
rect 32321 4777 32355 4811
rect 33425 4777 33459 4811
rect 35265 4777 35299 4811
rect 1593 4709 1627 4743
rect 3893 4709 3927 4743
rect 9597 4709 9631 4743
rect 37197 4709 37231 4743
rect 25973 4641 26007 4675
rect 1409 4573 1443 4607
rect 2053 4573 2087 4607
rect 2697 4573 2731 4607
rect 5365 4573 5399 4607
rect 7113 4573 7147 4607
rect 9045 4573 9079 4607
rect 11345 4573 11379 4607
rect 13001 4573 13035 4607
rect 14289 4573 14323 4607
rect 15761 4573 15795 4607
rect 16589 4573 16623 4607
rect 20085 4573 20119 4607
rect 20913 4573 20947 4607
rect 21557 4573 21591 4607
rect 22201 4573 22235 4607
rect 25329 4573 25363 4607
rect 26433 4573 26467 4607
rect 26617 4573 26651 4607
rect 26709 4573 26743 4607
rect 30389 4573 30423 4607
rect 31033 4573 31067 4607
rect 32137 4573 32171 4607
rect 33241 4573 33275 4607
rect 33977 4573 34011 4607
rect 36093 4573 36127 4607
rect 38117 4573 38151 4607
rect 8217 4505 8251 4539
rect 9321 4505 9355 4539
rect 12265 4505 12299 4539
rect 27997 4505 28031 4539
rect 35173 4505 35207 4539
rect 37381 4505 37415 4539
rect 2237 4437 2271 4471
rect 2881 4437 2915 4471
rect 4353 4437 4387 4471
rect 5549 4437 5583 4471
rect 6653 4437 6687 4471
rect 7297 4437 7331 4471
rect 9137 4437 9171 4471
rect 10149 4437 10183 4471
rect 11161 4437 11195 4471
rect 12817 4437 12851 4471
rect 13461 4437 13495 4471
rect 14933 4437 14967 4471
rect 15577 4437 15611 4471
rect 16405 4437 16439 4471
rect 17049 4437 17083 4471
rect 17601 4437 17635 4471
rect 18153 4437 18187 4471
rect 19625 4437 19659 4471
rect 20269 4437 20303 4471
rect 21097 4437 21131 4471
rect 21741 4437 21775 4471
rect 22385 4437 22419 4471
rect 22937 4437 22971 4471
rect 23857 4437 23891 4471
rect 24685 4437 24719 4471
rect 28549 4437 28583 4471
rect 29561 4437 29595 4471
rect 31217 4437 31251 4471
rect 34161 4437 34195 4471
rect 36277 4437 36311 4471
rect 2789 4233 2823 4267
rect 4445 4233 4479 4267
rect 19257 4233 19291 4267
rect 20545 4233 20579 4267
rect 20913 4233 20947 4267
rect 24501 4233 24535 4267
rect 7481 4165 7515 4199
rect 10149 4165 10183 4199
rect 36553 4165 36587 4199
rect 1409 4097 1443 4131
rect 2881 4097 2915 4131
rect 3617 4097 3651 4131
rect 4261 4097 4295 4131
rect 4905 4097 4939 4131
rect 5549 4097 5583 4131
rect 6469 4097 6503 4131
rect 8677 4097 8711 4131
rect 11897 4097 11931 4131
rect 12541 4097 12575 4131
rect 13001 4097 13035 4131
rect 13737 4097 13771 4131
rect 14749 4097 14783 4131
rect 15485 4097 15519 4131
rect 17417 4097 17451 4131
rect 19349 4097 19383 4131
rect 22385 4097 22419 4131
rect 23213 4097 23247 4131
rect 24041 4097 24075 4131
rect 25237 4097 25271 4131
rect 27169 4097 27203 4131
rect 27813 4097 27847 4131
rect 28641 4097 28675 4131
rect 30297 4097 30331 4131
rect 30481 4097 30515 4131
rect 31033 4097 31067 4131
rect 32137 4097 32171 4131
rect 32873 4097 32907 4131
rect 33977 4097 34011 4131
rect 35265 4097 35299 4131
rect 36369 4097 36403 4131
rect 37289 4097 37323 4131
rect 38117 4097 38151 4131
rect 3065 4029 3099 4063
rect 8953 4029 8987 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 19073 4029 19107 4063
rect 20269 4029 20303 4063
rect 20453 4029 20487 4063
rect 25697 4029 25731 4063
rect 26157 4029 26191 4063
rect 29837 4029 29871 4063
rect 2421 3961 2455 3995
rect 3801 3961 3835 3995
rect 5089 3961 5123 3995
rect 5733 3961 5767 3995
rect 7665 3961 7699 3995
rect 12357 3961 12391 3995
rect 13921 3961 13955 3995
rect 17969 3961 18003 3995
rect 19717 3961 19751 3995
rect 25053 3961 25087 3995
rect 26065 3961 26099 3995
rect 27629 3961 27663 3995
rect 29469 3961 29503 3995
rect 34161 3961 34195 3995
rect 37473 3961 37507 3995
rect 1593 3893 1627 3927
rect 6653 3893 6687 3927
rect 8125 3893 8159 3927
rect 10609 3893 10643 3927
rect 11713 3893 11747 3927
rect 13185 3893 13219 3927
rect 14565 3893 14599 3927
rect 15301 3893 15335 3927
rect 16129 3893 16163 3927
rect 17233 3893 17267 3927
rect 18429 3893 18463 3927
rect 22201 3893 22235 3927
rect 23029 3893 23063 3927
rect 23857 3893 23891 3927
rect 26985 3893 27019 3927
rect 28825 3893 28859 3927
rect 29377 3893 29411 3927
rect 31217 3893 31251 3927
rect 32321 3893 32355 3927
rect 33057 3893 33091 3927
rect 34713 3893 34747 3927
rect 35449 3893 35483 3927
rect 4997 3689 5031 3723
rect 6193 3689 6227 3723
rect 11529 3689 11563 3723
rect 13185 3689 13219 3723
rect 14105 3689 14139 3723
rect 16497 3689 16531 3723
rect 19349 3689 19383 3723
rect 19993 3689 20027 3723
rect 20729 3689 20763 3723
rect 21373 3689 21407 3723
rect 25605 3689 25639 3723
rect 29009 3689 29043 3723
rect 31493 3689 31527 3723
rect 7757 3621 7791 3655
rect 8401 3621 8435 3655
rect 22569 3621 22603 3655
rect 24777 3621 24811 3655
rect 36185 3621 36219 3655
rect 2053 3553 2087 3587
rect 5549 3553 5583 3587
rect 6745 3553 6779 3587
rect 9505 3553 9539 3587
rect 12541 3553 12575 3587
rect 12725 3553 12759 3587
rect 14657 3553 14691 3587
rect 15853 3553 15887 3587
rect 17601 3553 17635 3587
rect 22017 3553 22051 3587
rect 23121 3553 23155 3587
rect 30021 3553 30055 3587
rect 37841 3553 37875 3587
rect 1777 3485 1811 3519
rect 3249 3485 3283 3519
rect 3801 3485 3835 3519
rect 8217 3485 8251 3519
rect 9781 3485 9815 3519
rect 11253 3485 11287 3519
rect 14473 3485 14507 3519
rect 16129 3485 16163 3519
rect 17325 3485 17359 3519
rect 18429 3485 18463 3519
rect 19533 3485 19567 3519
rect 20545 3485 20579 3519
rect 21189 3485 21223 3519
rect 22201 3485 22235 3519
rect 23397 3485 23431 3519
rect 24593 3485 24627 3519
rect 25237 3485 25271 3519
rect 26525 3485 26559 3519
rect 26985 3485 27019 3519
rect 27813 3485 27847 3519
rect 28641 3485 28675 3519
rect 30297 3485 30331 3519
rect 32045 3485 32079 3519
rect 32781 3485 32815 3519
rect 33885 3485 33919 3519
rect 35265 3485 35299 3519
rect 38117 3485 38151 3519
rect 6653 3417 6687 3451
rect 7573 3417 7607 3451
rect 8953 3417 8987 3451
rect 10977 3417 11011 3451
rect 14565 3417 14599 3451
rect 22109 3417 22143 3451
rect 23305 3417 23339 3451
rect 25421 3417 25455 3451
rect 28825 3417 28859 3451
rect 31401 3417 31435 3451
rect 35081 3417 35115 3451
rect 36369 3417 36403 3451
rect 3065 3349 3099 3383
rect 3985 3349 4019 3383
rect 4537 3349 4571 3383
rect 5365 3349 5399 3383
rect 5457 3349 5491 3383
rect 6561 3349 6595 3383
rect 11069 3349 11103 3383
rect 12817 3349 12851 3383
rect 16037 3349 16071 3383
rect 16957 3349 16991 3383
rect 17417 3349 17451 3383
rect 18245 3349 18279 3383
rect 23765 3349 23799 3383
rect 26341 3349 26375 3383
rect 27169 3349 27203 3383
rect 27997 3349 28031 3383
rect 32229 3349 32263 3383
rect 32965 3349 32999 3383
rect 34069 3349 34103 3383
rect 2973 3145 3007 3179
rect 3433 3145 3467 3179
rect 4813 3145 4847 3179
rect 5825 3145 5859 3179
rect 9597 3145 9631 3179
rect 12449 3145 12483 3179
rect 13737 3145 13771 3179
rect 14565 3145 14599 3179
rect 15393 3145 15427 3179
rect 15945 3145 15979 3179
rect 16865 3145 16899 3179
rect 18613 3145 18647 3179
rect 20085 3145 20119 3179
rect 3985 3077 4019 3111
rect 4721 3077 4755 3111
rect 6837 3077 6871 3111
rect 7021 3077 7055 3111
rect 17969 3077 18003 3111
rect 24041 3077 24075 3111
rect 24225 3077 24259 3111
rect 24777 3077 24811 3111
rect 24961 3077 24995 3111
rect 27721 3077 27755 3111
rect 28365 3077 28399 3111
rect 29745 3077 29779 3111
rect 35725 3077 35759 3111
rect 1409 3009 1443 3043
rect 3065 3009 3099 3043
rect 5641 3009 5675 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 9413 3009 9447 3043
rect 10057 3009 10091 3043
rect 10333 3009 10367 3043
rect 11529 3009 11563 3043
rect 12265 3009 12299 3043
rect 13001 3009 13035 3043
rect 13921 3009 13955 3043
rect 14381 3009 14415 3043
rect 15209 3009 15243 3043
rect 16129 3009 16163 3043
rect 16681 3009 16715 3043
rect 17785 3009 17819 3043
rect 18429 3009 18463 3043
rect 19441 3009 19475 3043
rect 19901 3009 19935 3043
rect 21005 3009 21039 3043
rect 22109 3009 22143 3043
rect 22661 3009 22695 3043
rect 25421 3009 25455 3043
rect 26157 3009 26191 3043
rect 29009 3009 29043 3043
rect 29561 3009 29595 3043
rect 30573 3009 30607 3043
rect 30849 3009 30883 3043
rect 32505 3009 32539 3043
rect 32781 3009 32815 3043
rect 33793 3009 33827 3043
rect 34897 3009 34931 3043
rect 35081 3009 35115 3043
rect 36461 3009 36495 3043
rect 37289 3009 37323 3043
rect 37565 3009 37599 3043
rect 1685 2941 1719 2975
rect 2881 2941 2915 2975
rect 22937 2941 22971 2975
rect 4169 2873 4203 2907
rect 13185 2873 13219 2907
rect 26341 2873 26375 2907
rect 27537 2873 27571 2907
rect 28825 2873 28859 2907
rect 36645 2873 36679 2907
rect 7573 2805 7607 2839
rect 11713 2805 11747 2839
rect 19257 2805 19291 2839
rect 20821 2805 20855 2839
rect 21925 2805 21959 2839
rect 25605 2805 25639 2839
rect 26985 2805 27019 2839
rect 33977 2805 34011 2839
rect 35633 2805 35667 2839
rect 6607 2601 6641 2635
rect 10701 2601 10735 2635
rect 13369 2601 13403 2635
rect 15117 2601 15151 2635
rect 16865 2601 16899 2635
rect 17601 2601 17635 2635
rect 28825 2601 28859 2635
rect 34897 2601 34931 2635
rect 4077 2533 4111 2567
rect 12817 2533 12851 2567
rect 15945 2533 15979 2567
rect 18521 2533 18555 2567
rect 20545 2533 20579 2567
rect 26157 2533 26191 2567
rect 27353 2533 27387 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 4537 2465 4571 2499
rect 4813 2465 4847 2499
rect 9229 2465 9263 2499
rect 21925 2465 21959 2499
rect 22385 2465 22419 2499
rect 22661 2465 22695 2499
rect 29745 2465 29779 2499
rect 30021 2465 30055 2499
rect 32505 2465 32539 2499
rect 35909 2465 35943 2499
rect 37289 2465 37323 2499
rect 37565 2465 37599 2499
rect 2789 2397 2823 2431
rect 6377 2397 6411 2431
rect 7757 2397 7791 2431
rect 9505 2397 9539 2431
rect 10609 2397 10643 2431
rect 11989 2397 12023 2431
rect 12633 2397 12667 2431
rect 14105 2397 14139 2431
rect 14933 2397 14967 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 19901 2397 19935 2431
rect 20361 2397 20395 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 24685 2397 24719 2431
rect 26341 2397 26375 2431
rect 28273 2397 28307 2431
rect 29009 2397 29043 2431
rect 31217 2397 31251 2431
rect 32229 2397 32263 2431
rect 34069 2397 34103 2431
rect 34713 2397 34747 2431
rect 36185 2397 36219 2431
rect 3893 2329 3927 2363
rect 7941 2329 7975 2363
rect 18337 2329 18371 2363
rect 19717 2329 19751 2363
rect 21281 2329 21315 2363
rect 27537 2329 27571 2363
rect 2881 2261 2915 2295
rect 12081 2261 12115 2295
rect 14289 2261 14323 2295
rect 23857 2261 23891 2295
rect 28181 2261 28215 2295
rect 31125 2261 31159 2295
rect 33977 2261 34011 2295
<< metal1 >>
rect 2222 37816 2228 37868
rect 2280 37856 2286 37868
rect 23658 37856 23664 37868
rect 2280 37828 23664 37856
rect 2280 37816 2286 37828
rect 23658 37816 23664 37828
rect 23716 37816 23722 37868
rect 7282 37748 7288 37800
rect 7340 37788 7346 37800
rect 26694 37788 26700 37800
rect 7340 37760 26700 37788
rect 7340 37748 7346 37760
rect 26694 37748 26700 37760
rect 26752 37748 26758 37800
rect 12250 37680 12256 37732
rect 12308 37720 12314 37732
rect 31478 37720 31484 37732
rect 12308 37692 31484 37720
rect 12308 37680 12314 37692
rect 31478 37680 31484 37692
rect 31536 37680 31542 37732
rect 13170 37612 13176 37664
rect 13228 37652 13234 37664
rect 31570 37652 31576 37664
rect 13228 37624 31576 37652
rect 13228 37612 13234 37624
rect 31570 37612 31576 37624
rect 31628 37612 31634 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 2133 37451 2191 37457
rect 2133 37417 2145 37451
rect 2179 37448 2191 37451
rect 2222 37448 2228 37460
rect 2179 37420 2228 37448
rect 2179 37417 2191 37420
rect 2133 37411 2191 37417
rect 2222 37408 2228 37420
rect 2280 37408 2286 37460
rect 4249 37451 4307 37457
rect 4249 37417 4261 37451
rect 4295 37448 4307 37451
rect 4890 37448 4896 37460
rect 4295 37420 4896 37448
rect 4295 37417 4307 37420
rect 4249 37411 4307 37417
rect 4890 37408 4896 37420
rect 4948 37408 4954 37460
rect 7101 37451 7159 37457
rect 7101 37417 7113 37451
rect 7147 37448 7159 37451
rect 7282 37448 7288 37460
rect 7147 37420 7288 37448
rect 7147 37417 7159 37420
rect 7101 37411 7159 37417
rect 7282 37408 7288 37420
rect 7340 37408 7346 37460
rect 12250 37448 12256 37460
rect 12211 37420 12256 37448
rect 12250 37408 12256 37420
rect 12308 37408 12314 37460
rect 29086 37448 29092 37460
rect 12406 37420 29092 37448
rect 9677 37383 9735 37389
rect 9677 37349 9689 37383
rect 9723 37380 9735 37383
rect 12406 37380 12434 37420
rect 29086 37408 29092 37420
rect 29144 37408 29150 37460
rect 13170 37380 13176 37392
rect 9723 37352 12434 37380
rect 13131 37352 13176 37380
rect 9723 37349 9735 37352
rect 9677 37343 9735 37349
rect 13170 37340 13176 37352
rect 13228 37340 13234 37392
rect 15933 37383 15991 37389
rect 15933 37380 15945 37383
rect 14568 37352 15945 37380
rect 2961 37315 3019 37321
rect 2961 37281 2973 37315
rect 3007 37312 3019 37315
rect 3694 37312 3700 37324
rect 3007 37284 3700 37312
rect 3007 37281 3019 37284
rect 2961 37275 3019 37281
rect 3694 37272 3700 37284
rect 3752 37272 3758 37324
rect 4893 37315 4951 37321
rect 4893 37281 4905 37315
rect 4939 37312 4951 37315
rect 5258 37312 5264 37324
rect 4939 37284 5264 37312
rect 4939 37281 4951 37284
rect 4893 37275 4951 37281
rect 5258 37272 5264 37284
rect 5316 37272 5322 37324
rect 1118 37204 1124 37256
rect 1176 37244 1182 37256
rect 1857 37247 1915 37253
rect 1857 37244 1869 37247
rect 1176 37216 1869 37244
rect 1176 37204 1182 37216
rect 1857 37213 1869 37216
rect 1903 37244 1915 37247
rect 1946 37244 1952 37256
rect 1903 37216 1952 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 1946 37204 1952 37216
rect 2004 37204 2010 37256
rect 2130 37204 2136 37256
rect 2188 37244 2194 37256
rect 2590 37244 2596 37256
rect 2188 37216 2596 37244
rect 2188 37204 2194 37216
rect 2590 37204 2596 37216
rect 2648 37244 2654 37256
rect 2777 37247 2835 37253
rect 2777 37244 2789 37247
rect 2648 37216 2789 37244
rect 2648 37204 2654 37216
rect 2777 37213 2789 37216
rect 2823 37213 2835 37247
rect 2777 37207 2835 37213
rect 4154 37204 4160 37256
rect 4212 37244 4218 37256
rect 5074 37244 5080 37256
rect 4212 37216 5080 37244
rect 4212 37204 4218 37216
rect 5074 37204 5080 37216
rect 5132 37204 5138 37256
rect 5718 37204 5724 37256
rect 5776 37244 5782 37256
rect 5813 37247 5871 37253
rect 5813 37244 5825 37247
rect 5776 37216 5825 37244
rect 5776 37204 5782 37216
rect 5813 37213 5825 37216
rect 5859 37213 5871 37247
rect 5813 37207 5871 37213
rect 6362 37204 6368 37256
rect 6420 37244 6426 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6420 37216 6837 37244
rect 6420 37204 6426 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 6825 37207 6883 37213
rect 7466 37204 7472 37256
rect 7524 37244 7530 37256
rect 7653 37247 7711 37253
rect 7653 37244 7665 37247
rect 7524 37216 7665 37244
rect 7524 37204 7530 37216
rect 7653 37213 7665 37216
rect 7699 37213 7711 37247
rect 7653 37207 7711 37213
rect 8478 37204 8484 37256
rect 8536 37244 8542 37256
rect 9398 37244 9404 37256
rect 8536 37216 9404 37244
rect 8536 37204 8542 37216
rect 9398 37204 9404 37216
rect 9456 37204 9462 37256
rect 10134 37204 10140 37256
rect 10192 37244 10198 37256
rect 10229 37247 10287 37253
rect 10229 37244 10241 37247
rect 10192 37216 10241 37244
rect 10192 37204 10198 37216
rect 10229 37213 10241 37216
rect 10275 37213 10287 37247
rect 10229 37207 10287 37213
rect 10594 37204 10600 37256
rect 10652 37244 10658 37256
rect 11977 37247 12035 37253
rect 11977 37244 11989 37247
rect 10652 37216 11989 37244
rect 10652 37204 10658 37216
rect 11977 37213 11989 37216
rect 12023 37244 12035 37247
rect 12158 37244 12164 37256
rect 12023 37216 12164 37244
rect 12023 37213 12035 37216
rect 11977 37207 12035 37213
rect 12158 37204 12164 37216
rect 12216 37204 12222 37256
rect 13814 37204 13820 37256
rect 13872 37244 13878 37256
rect 14568 37253 14596 37352
rect 15933 37349 15945 37352
rect 15979 37349 15991 37383
rect 15933 37343 15991 37349
rect 18417 37383 18475 37389
rect 18417 37349 18429 37383
rect 18463 37380 18475 37383
rect 35986 37380 35992 37392
rect 18463 37352 35992 37380
rect 18463 37349 18475 37352
rect 18417 37343 18475 37349
rect 35986 37340 35992 37352
rect 36044 37340 36050 37392
rect 15473 37315 15531 37321
rect 15473 37281 15485 37315
rect 15519 37312 15531 37315
rect 15838 37312 15844 37324
rect 15519 37284 15844 37312
rect 15519 37281 15531 37284
rect 15473 37275 15531 37281
rect 15838 37272 15844 37284
rect 15896 37272 15902 37324
rect 17037 37315 17095 37321
rect 17037 37281 17049 37315
rect 17083 37312 17095 37315
rect 17402 37312 17408 37324
rect 17083 37284 17408 37312
rect 17083 37281 17095 37284
rect 17037 37275 17095 37281
rect 17402 37272 17408 37284
rect 17460 37272 17466 37324
rect 21910 37272 21916 37324
rect 21968 37312 21974 37324
rect 22189 37315 22247 37321
rect 22189 37312 22201 37315
rect 21968 37284 22201 37312
rect 21968 37272 21974 37284
rect 22189 37281 22201 37284
rect 22235 37281 22247 37315
rect 23661 37315 23719 37321
rect 23661 37312 23673 37315
rect 22189 37275 22247 37281
rect 22388 37284 23673 37312
rect 14553 37247 14611 37253
rect 14553 37244 14565 37247
rect 13872 37216 14565 37244
rect 13872 37204 13878 37216
rect 14553 37213 14565 37216
rect 14599 37213 14611 37247
rect 14553 37207 14611 37213
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15102 37244 15108 37256
rect 14884 37216 15108 37244
rect 14884 37204 14890 37216
rect 15102 37204 15108 37216
rect 15160 37244 15166 37256
rect 15289 37247 15347 37253
rect 15289 37244 15301 37247
rect 15160 37216 15301 37244
rect 15160 37204 15166 37216
rect 15289 37213 15301 37216
rect 15335 37213 15347 37247
rect 15289 37207 15347 37213
rect 15930 37204 15936 37256
rect 15988 37244 15994 37256
rect 17221 37247 17279 37253
rect 17221 37244 17233 37247
rect 15988 37216 17233 37244
rect 15988 37204 15994 37216
rect 17221 37213 17233 37216
rect 17267 37244 17279 37247
rect 17494 37244 17500 37256
rect 17267 37216 17500 37244
rect 17267 37213 17279 37216
rect 17221 37207 17279 37213
rect 17494 37204 17500 37216
rect 17552 37204 17558 37256
rect 17954 37204 17960 37256
rect 18012 37244 18018 37256
rect 18141 37247 18199 37253
rect 18141 37244 18153 37247
rect 18012 37216 18153 37244
rect 18012 37204 18018 37216
rect 18141 37213 18153 37216
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 19058 37204 19064 37256
rect 19116 37244 19122 37256
rect 19245 37247 19303 37253
rect 19245 37244 19257 37247
rect 19116 37216 19257 37244
rect 19116 37204 19122 37216
rect 19245 37213 19257 37216
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 20070 37204 20076 37256
rect 20128 37244 20134 37256
rect 20165 37247 20223 37253
rect 20165 37244 20177 37247
rect 20128 37216 20177 37244
rect 20128 37204 20134 37216
rect 20165 37213 20177 37216
rect 20211 37213 20223 37247
rect 20898 37244 20904 37256
rect 20859 37216 20904 37244
rect 20165 37207 20223 37213
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 21082 37204 21088 37256
rect 21140 37244 21146 37256
rect 22388 37253 22416 37284
rect 23661 37281 23673 37284
rect 23707 37281 23719 37315
rect 30650 37312 30656 37324
rect 30611 37284 30656 37312
rect 23661 37275 23719 37281
rect 30650 37272 30656 37284
rect 30708 37272 30714 37324
rect 32490 37312 32496 37324
rect 32451 37284 32496 37312
rect 32490 37272 32496 37284
rect 32548 37272 32554 37324
rect 33965 37315 34023 37321
rect 33965 37312 33977 37315
rect 32692 37284 33977 37312
rect 22373 37247 22431 37253
rect 22373 37244 22385 37247
rect 21140 37216 22385 37244
rect 21140 37204 21146 37216
rect 22373 37213 22385 37216
rect 22419 37213 22431 37247
rect 22373 37207 22431 37213
rect 22925 37247 22983 37253
rect 22925 37213 22937 37247
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 3234 37136 3240 37188
rect 3292 37176 3298 37188
rect 4062 37176 4068 37188
rect 3292 37148 4068 37176
rect 3292 37136 3298 37148
rect 4062 37136 4068 37148
rect 4120 37176 4126 37188
rect 4341 37179 4399 37185
rect 4341 37176 4353 37179
rect 4120 37148 4353 37176
rect 4120 37136 4126 37148
rect 4341 37145 4353 37148
rect 4387 37145 4399 37179
rect 4341 37139 4399 37145
rect 11606 37136 11612 37188
rect 11664 37176 11670 37188
rect 12897 37179 12955 37185
rect 12897 37176 12909 37179
rect 11664 37148 12909 37176
rect 11664 37136 11670 37148
rect 12897 37145 12909 37148
rect 12943 37176 12955 37179
rect 13170 37176 13176 37188
rect 12943 37148 13176 37176
rect 12943 37145 12955 37148
rect 12897 37139 12955 37145
rect 13170 37136 13176 37148
rect 13228 37136 13234 37188
rect 18046 37136 18052 37188
rect 18104 37176 18110 37188
rect 18104 37148 22094 37176
rect 18104 37136 18110 37148
rect 3050 37068 3056 37120
rect 3108 37108 3114 37120
rect 5629 37111 5687 37117
rect 5629 37108 5641 37111
rect 3108 37080 5641 37108
rect 3108 37068 3114 37080
rect 5629 37077 5641 37080
rect 5675 37077 5687 37111
rect 7834 37108 7840 37120
rect 7795 37080 7840 37108
rect 5629 37071 5687 37077
rect 7834 37068 7840 37080
rect 7892 37068 7898 37120
rect 10410 37108 10416 37120
rect 10371 37080 10416 37108
rect 10410 37068 10416 37080
rect 10468 37068 10474 37120
rect 13998 37068 14004 37120
rect 14056 37108 14062 37120
rect 14645 37111 14703 37117
rect 14645 37108 14657 37111
rect 14056 37080 14657 37108
rect 14056 37068 14062 37080
rect 14645 37077 14657 37080
rect 14691 37077 14703 37111
rect 19426 37108 19432 37120
rect 19387 37080 19432 37108
rect 14645 37071 14703 37077
rect 19426 37068 19432 37080
rect 19484 37068 19490 37120
rect 20346 37108 20352 37120
rect 20307 37080 20352 37108
rect 20346 37068 20352 37080
rect 20404 37068 20410 37120
rect 20438 37068 20444 37120
rect 20496 37108 20502 37120
rect 21085 37111 21143 37117
rect 21085 37108 21097 37111
rect 20496 37080 21097 37108
rect 20496 37068 20502 37080
rect 21085 37077 21097 37080
rect 21131 37077 21143 37111
rect 22066 37108 22094 37148
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 22940 37176 22968 37207
rect 24302 37204 24308 37256
rect 24360 37244 24366 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 24360 37216 24409 37244
rect 24360 37204 24366 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 25314 37204 25320 37256
rect 25372 37244 25378 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25372 37216 25421 37244
rect 25372 37204 25378 37216
rect 25409 37213 25421 37216
rect 25455 37213 25467 37247
rect 25409 37207 25467 37213
rect 25498 37204 25504 37256
rect 25556 37244 25562 37256
rect 26145 37247 26203 37253
rect 26145 37244 26157 37247
rect 25556 37216 26157 37244
rect 25556 37204 25562 37216
rect 26145 37213 26157 37216
rect 26191 37213 26203 37247
rect 26970 37244 26976 37256
rect 26931 37216 26976 37244
rect 26145 37207 26203 37213
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27893 37247 27951 37253
rect 27893 37213 27905 37247
rect 27939 37213 27951 37247
rect 27893 37207 27951 37213
rect 24118 37176 24124 37188
rect 22244 37148 22968 37176
rect 23032 37148 24124 37176
rect 22244 37136 22250 37148
rect 23032 37108 23060 37148
rect 24118 37136 24124 37148
rect 24176 37136 24182 37188
rect 26602 37136 26608 37188
rect 26660 37176 26666 37188
rect 27908 37176 27936 37207
rect 28534 37204 28540 37256
rect 28592 37244 28598 37256
rect 28810 37244 28816 37256
rect 28592 37216 28816 37244
rect 28592 37204 28598 37216
rect 28810 37204 28816 37216
rect 28868 37204 28874 37256
rect 29546 37244 29552 37256
rect 29507 37216 29552 37244
rect 29546 37204 29552 37216
rect 29604 37204 29610 37256
rect 30558 37204 30564 37256
rect 30616 37244 30622 37256
rect 30837 37247 30895 37253
rect 30837 37244 30849 37247
rect 30616 37216 30849 37244
rect 30616 37204 30622 37216
rect 30837 37213 30849 37216
rect 30883 37213 30895 37247
rect 30837 37207 30895 37213
rect 31202 37204 31208 37256
rect 31260 37244 31266 37256
rect 31573 37247 31631 37253
rect 31573 37244 31585 37247
rect 31260 37216 31585 37244
rect 31260 37204 31266 37216
rect 31573 37213 31585 37216
rect 31619 37213 31631 37247
rect 31573 37207 31631 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32692 37253 32720 37284
rect 33965 37281 33977 37284
rect 34011 37281 34023 37315
rect 38013 37315 38071 37321
rect 38013 37312 38025 37315
rect 33965 37275 34023 37281
rect 34716 37284 34928 37312
rect 32677 37247 32735 37253
rect 32677 37244 32689 37247
rect 31812 37216 32689 37244
rect 31812 37204 31818 37216
rect 32677 37213 32689 37216
rect 32723 37213 32735 37247
rect 32677 37207 32735 37213
rect 32766 37204 32772 37256
rect 32824 37244 32830 37256
rect 33502 37244 33508 37256
rect 32824 37216 33508 37244
rect 32824 37204 32830 37216
rect 33502 37204 33508 37216
rect 33560 37204 33566 37256
rect 33778 37204 33784 37256
rect 33836 37244 33842 37256
rect 34716 37244 34744 37284
rect 33836 37216 34744 37244
rect 34900 37244 34928 37284
rect 36464 37284 38025 37312
rect 34977 37247 35035 37253
rect 34977 37244 34989 37247
rect 34900 37216 34989 37244
rect 33836 37204 33842 37216
rect 34977 37213 34989 37216
rect 35023 37244 35035 37247
rect 35434 37244 35440 37256
rect 35023 37216 35440 37244
rect 35023 37213 35035 37216
rect 34977 37207 35035 37213
rect 35434 37204 35440 37216
rect 35492 37204 35498 37256
rect 35710 37244 35716 37256
rect 35671 37216 35716 37244
rect 35710 37204 35716 37216
rect 35768 37204 35774 37256
rect 35894 37204 35900 37256
rect 35952 37244 35958 37256
rect 36464 37253 36492 37284
rect 38013 37281 38025 37284
rect 38059 37281 38071 37315
rect 38013 37275 38071 37281
rect 36449 37247 36507 37253
rect 36449 37244 36461 37247
rect 35952 37216 36461 37244
rect 35952 37204 35958 37216
rect 36449 37213 36461 37216
rect 36495 37213 36507 37247
rect 37274 37244 37280 37256
rect 37235 37216 37280 37244
rect 36449 37207 36507 37213
rect 37274 37204 37280 37216
rect 37332 37204 37338 37256
rect 26660 37148 27936 37176
rect 26660 37136 26666 37148
rect 28442 37136 28448 37188
rect 28500 37176 28506 37188
rect 34330 37176 34336 37188
rect 28500 37148 31432 37176
rect 28500 37136 28506 37148
rect 22066 37080 23060 37108
rect 23109 37111 23167 37117
rect 21085 37071 21143 37077
rect 23109 37077 23121 37111
rect 23155 37108 23167 37111
rect 23290 37108 23296 37120
rect 23155 37080 23296 37108
rect 23155 37077 23167 37080
rect 23109 37071 23167 37077
rect 23290 37068 23296 37080
rect 23348 37068 23354 37120
rect 24578 37108 24584 37120
rect 24539 37080 24584 37108
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 25590 37108 25596 37120
rect 25551 37080 25596 37108
rect 25590 37068 25596 37080
rect 25648 37068 25654 37120
rect 25682 37068 25688 37120
rect 25740 37108 25746 37120
rect 26329 37111 26387 37117
rect 26329 37108 26341 37111
rect 25740 37080 26341 37108
rect 25740 37068 25746 37080
rect 26329 37077 26341 37080
rect 26375 37077 26387 37111
rect 26329 37071 26387 37077
rect 26786 37068 26792 37120
rect 26844 37108 26850 37120
rect 27157 37111 27215 37117
rect 27157 37108 27169 37111
rect 26844 37080 27169 37108
rect 26844 37068 26850 37080
rect 27157 37077 27169 37080
rect 27203 37077 27215 37111
rect 27157 37071 27215 37077
rect 27798 37068 27804 37120
rect 27856 37108 27862 37120
rect 28077 37111 28135 37117
rect 28077 37108 28089 37111
rect 27856 37080 28089 37108
rect 27856 37068 27862 37080
rect 28077 37077 28089 37080
rect 28123 37077 28135 37111
rect 28718 37108 28724 37120
rect 28679 37080 28724 37108
rect 28077 37071 28135 37077
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 29730 37108 29736 37120
rect 29691 37080 29736 37108
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 31202 37108 31208 37120
rect 29880 37080 31208 37108
rect 29880 37068 29886 37080
rect 31202 37068 31208 37080
rect 31260 37068 31266 37120
rect 31404 37117 31432 37148
rect 33336 37148 34336 37176
rect 33336 37117 33364 37148
rect 34330 37136 34336 37148
rect 34388 37136 34394 37188
rect 38378 37176 38384 37188
rect 37476 37148 38384 37176
rect 31389 37111 31447 37117
rect 31389 37077 31401 37111
rect 31435 37077 31447 37111
rect 31389 37071 31447 37077
rect 33321 37111 33379 37117
rect 33321 37077 33333 37111
rect 33367 37077 33379 37111
rect 34790 37108 34796 37120
rect 34751 37080 34796 37108
rect 33321 37071 33379 37077
rect 34790 37068 34796 37080
rect 34848 37068 34854 37120
rect 35526 37108 35532 37120
rect 35487 37080 35532 37108
rect 35526 37068 35532 37080
rect 35584 37068 35590 37120
rect 36262 37108 36268 37120
rect 36223 37080 36268 37108
rect 36262 37068 36268 37080
rect 36320 37068 36326 37120
rect 37476 37117 37504 37148
rect 38378 37136 38384 37148
rect 38436 37136 38442 37188
rect 37461 37111 37519 37117
rect 37461 37077 37473 37111
rect 37507 37077 37519 37111
rect 37461 37071 37519 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 2498 36864 2504 36916
rect 2556 36904 2562 36916
rect 3421 36907 3479 36913
rect 3421 36904 3433 36907
rect 2556 36876 3433 36904
rect 2556 36864 2562 36876
rect 3421 36873 3433 36876
rect 3467 36873 3479 36907
rect 3421 36867 3479 36873
rect 3602 36864 3608 36916
rect 3660 36904 3666 36916
rect 4065 36907 4123 36913
rect 4065 36904 4077 36907
rect 3660 36876 4077 36904
rect 3660 36864 3666 36876
rect 4065 36873 4077 36876
rect 4111 36873 4123 36907
rect 4065 36867 4123 36873
rect 4614 36864 4620 36916
rect 4672 36904 4678 36916
rect 4801 36907 4859 36913
rect 4801 36904 4813 36907
rect 4672 36876 4813 36904
rect 4672 36864 4678 36876
rect 4801 36873 4813 36876
rect 4847 36873 4859 36907
rect 4801 36867 4859 36873
rect 4982 36864 4988 36916
rect 5040 36904 5046 36916
rect 5629 36907 5687 36913
rect 5629 36904 5641 36907
rect 5040 36876 5641 36904
rect 5040 36864 5046 36876
rect 5629 36873 5641 36876
rect 5675 36873 5687 36907
rect 5629 36867 5687 36873
rect 5810 36864 5816 36916
rect 5868 36904 5874 36916
rect 7285 36907 7343 36913
rect 7285 36904 7297 36907
rect 5868 36876 7297 36904
rect 5868 36864 5874 36876
rect 7285 36873 7297 36876
rect 7331 36873 7343 36907
rect 7285 36867 7343 36873
rect 7742 36864 7748 36916
rect 7800 36904 7806 36916
rect 8757 36907 8815 36913
rect 8757 36904 8769 36907
rect 7800 36876 8769 36904
rect 7800 36864 7806 36876
rect 8757 36873 8769 36876
rect 8803 36873 8815 36907
rect 8757 36867 8815 36873
rect 8846 36864 8852 36916
rect 8904 36904 8910 36916
rect 9401 36907 9459 36913
rect 9401 36904 9413 36907
rect 8904 36876 9413 36904
rect 8904 36864 8910 36876
rect 9401 36873 9413 36876
rect 9447 36873 9459 36907
rect 9401 36867 9459 36873
rect 10873 36907 10931 36913
rect 10873 36873 10885 36907
rect 10919 36904 10931 36907
rect 10962 36904 10968 36916
rect 10919 36876 10968 36904
rect 10919 36873 10931 36876
rect 10873 36867 10931 36873
rect 10962 36864 10968 36876
rect 11020 36864 11026 36916
rect 11974 36864 11980 36916
rect 12032 36904 12038 36916
rect 12161 36907 12219 36913
rect 12161 36904 12173 36907
rect 12032 36876 12173 36904
rect 12032 36864 12038 36876
rect 12161 36873 12173 36876
rect 12207 36873 12219 36907
rect 12161 36867 12219 36873
rect 13078 36864 13084 36916
rect 13136 36904 13142 36916
rect 13633 36907 13691 36913
rect 13633 36904 13645 36907
rect 13136 36876 13645 36904
rect 13136 36864 13142 36876
rect 13633 36873 13645 36876
rect 13679 36873 13691 36907
rect 13633 36867 13691 36873
rect 14090 36864 14096 36916
rect 14148 36904 14154 36916
rect 14461 36907 14519 36913
rect 14461 36904 14473 36907
rect 14148 36876 14473 36904
rect 14148 36864 14154 36876
rect 14461 36873 14473 36876
rect 14507 36873 14519 36907
rect 14461 36867 14519 36873
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 15749 36907 15807 36913
rect 15749 36904 15761 36907
rect 15252 36876 15761 36904
rect 15252 36864 15258 36876
rect 15749 36873 15761 36876
rect 15795 36873 15807 36907
rect 15749 36867 15807 36873
rect 17218 36864 17224 36916
rect 17276 36904 17282 36916
rect 17865 36907 17923 36913
rect 17865 36904 17877 36907
rect 17276 36876 17877 36904
rect 17276 36864 17282 36876
rect 17865 36873 17877 36876
rect 17911 36873 17923 36907
rect 17865 36867 17923 36873
rect 18322 36864 18328 36916
rect 18380 36904 18386 36916
rect 18601 36907 18659 36913
rect 18601 36904 18613 36907
rect 18380 36876 18613 36904
rect 18380 36864 18386 36876
rect 18601 36873 18613 36876
rect 18647 36873 18659 36907
rect 18601 36867 18659 36873
rect 19334 36864 19340 36916
rect 19392 36904 19398 36916
rect 19521 36907 19579 36913
rect 19521 36904 19533 36907
rect 19392 36876 19533 36904
rect 19392 36864 19398 36876
rect 19521 36873 19533 36876
rect 19567 36873 19579 36907
rect 19521 36867 19579 36873
rect 19978 36864 19984 36916
rect 20036 36904 20042 36916
rect 20257 36907 20315 36913
rect 20257 36904 20269 36907
rect 20036 36876 20269 36904
rect 20036 36864 20042 36876
rect 20257 36873 20269 36876
rect 20303 36873 20315 36907
rect 20257 36867 20315 36873
rect 20806 36864 20812 36916
rect 20864 36904 20870 36916
rect 21085 36907 21143 36913
rect 21085 36904 21097 36907
rect 20864 36876 21097 36904
rect 20864 36864 20870 36876
rect 21085 36873 21097 36876
rect 21131 36873 21143 36907
rect 21085 36867 21143 36873
rect 21450 36864 21456 36916
rect 21508 36904 21514 36916
rect 22005 36907 22063 36913
rect 22005 36904 22017 36907
rect 21508 36876 22017 36904
rect 21508 36864 21514 36876
rect 22005 36873 22017 36876
rect 22051 36873 22063 36907
rect 22005 36867 22063 36873
rect 22554 36864 22560 36916
rect 22612 36904 22618 36916
rect 22741 36907 22799 36913
rect 22741 36904 22753 36907
rect 22612 36876 22753 36904
rect 22612 36864 22618 36876
rect 22741 36873 22753 36876
rect 22787 36873 22799 36907
rect 22741 36867 22799 36873
rect 23566 36864 23572 36916
rect 23624 36904 23630 36916
rect 24213 36907 24271 36913
rect 24213 36904 24225 36907
rect 23624 36876 24225 36904
rect 23624 36864 23630 36876
rect 24213 36873 24225 36876
rect 24259 36873 24271 36907
rect 24213 36867 24271 36873
rect 24854 36864 24860 36916
rect 24912 36904 24918 36916
rect 24949 36907 25007 36913
rect 24949 36904 24961 36907
rect 24912 36876 24961 36904
rect 24912 36864 24918 36876
rect 24949 36873 24961 36876
rect 24995 36873 25007 36907
rect 24949 36867 25007 36873
rect 25038 36864 25044 36916
rect 25096 36904 25102 36916
rect 25685 36907 25743 36913
rect 25685 36904 25697 36907
rect 25096 36876 25697 36904
rect 25096 36864 25102 36876
rect 25685 36873 25697 36876
rect 25731 36873 25743 36907
rect 25685 36867 25743 36873
rect 27062 36864 27068 36916
rect 27120 36904 27126 36916
rect 27893 36907 27951 36913
rect 27893 36904 27905 36907
rect 27120 36876 27905 36904
rect 27120 36864 27126 36876
rect 27893 36873 27905 36876
rect 27939 36873 27951 36907
rect 27893 36867 27951 36873
rect 28166 36864 28172 36916
rect 28224 36904 28230 36916
rect 28537 36907 28595 36913
rect 28537 36904 28549 36907
rect 28224 36876 28549 36904
rect 28224 36864 28230 36876
rect 28537 36873 28549 36876
rect 28583 36873 28595 36907
rect 28537 36867 28595 36873
rect 29178 36864 29184 36916
rect 29236 36904 29242 36916
rect 29457 36907 29515 36913
rect 29457 36904 29469 36907
rect 29236 36876 29469 36904
rect 29236 36864 29242 36876
rect 29457 36873 29469 36876
rect 29503 36873 29515 36907
rect 29457 36867 29515 36873
rect 29914 36864 29920 36916
rect 29972 36904 29978 36916
rect 30193 36907 30251 36913
rect 30193 36904 30205 36907
rect 29972 36876 30205 36904
rect 29972 36864 29978 36876
rect 30193 36873 30205 36876
rect 30239 36873 30251 36907
rect 30193 36867 30251 36873
rect 30926 36864 30932 36916
rect 30984 36904 30990 36916
rect 31205 36907 31263 36913
rect 31205 36904 31217 36907
rect 30984 36876 31217 36904
rect 30984 36864 30990 36876
rect 31205 36873 31217 36876
rect 31251 36873 31263 36907
rect 31205 36867 31263 36873
rect 32030 36864 32036 36916
rect 32088 36904 32094 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 32088 36876 32321 36904
rect 32088 36864 32094 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 33134 36864 33140 36916
rect 33192 36904 33198 36916
rect 33321 36907 33379 36913
rect 33321 36904 33333 36907
rect 33192 36876 33333 36904
rect 33192 36864 33198 36876
rect 33321 36873 33333 36876
rect 33367 36873 33379 36907
rect 33321 36867 33379 36873
rect 34146 36864 34152 36916
rect 34204 36904 34210 36916
rect 34425 36907 34483 36913
rect 34425 36904 34437 36907
rect 34204 36876 34437 36904
rect 34204 36864 34210 36876
rect 34425 36873 34437 36876
rect 34471 36873 34483 36907
rect 34425 36867 34483 36873
rect 35342 36864 35348 36916
rect 35400 36904 35406 36916
rect 35437 36907 35495 36913
rect 35437 36904 35449 36907
rect 35400 36876 35449 36904
rect 35400 36864 35406 36876
rect 35437 36873 35449 36876
rect 35483 36873 35495 36907
rect 35437 36867 35495 36873
rect 36354 36864 36360 36916
rect 36412 36904 36418 36916
rect 36541 36907 36599 36913
rect 36541 36904 36553 36907
rect 36412 36876 36553 36904
rect 36412 36864 36418 36876
rect 36541 36873 36553 36876
rect 36587 36873 36599 36907
rect 36541 36867 36599 36873
rect 106 36796 112 36848
rect 164 36836 170 36848
rect 1578 36836 1584 36848
rect 164 36808 1584 36836
rect 164 36796 170 36808
rect 1578 36796 1584 36808
rect 1636 36836 1642 36848
rect 1857 36839 1915 36845
rect 1857 36836 1869 36839
rect 1636 36808 1869 36836
rect 1636 36796 1642 36808
rect 1857 36805 1869 36808
rect 1903 36805 1915 36839
rect 3050 36836 3056 36848
rect 1857 36799 1915 36805
rect 2792 36808 3056 36836
rect 2792 36777 2820 36808
rect 3050 36796 3056 36808
rect 3108 36796 3114 36848
rect 7466 36796 7472 36848
rect 7524 36836 7530 36848
rect 10045 36839 10103 36845
rect 10045 36836 10057 36839
rect 7524 36808 10057 36836
rect 7524 36796 7530 36808
rect 10045 36805 10057 36808
rect 10091 36805 10103 36839
rect 10045 36799 10103 36805
rect 12710 36796 12716 36848
rect 12768 36836 12774 36848
rect 12897 36839 12955 36845
rect 12897 36836 12909 36839
rect 12768 36808 12909 36836
rect 12768 36796 12774 36808
rect 12897 36805 12909 36808
rect 12943 36805 12955 36839
rect 12897 36799 12955 36805
rect 13170 36796 13176 36848
rect 13228 36836 13234 36848
rect 15013 36839 15071 36845
rect 15013 36836 15025 36839
rect 13228 36808 15025 36836
rect 13228 36796 13234 36808
rect 15013 36805 15025 36808
rect 15059 36805 15071 36839
rect 15013 36799 15071 36805
rect 16942 36796 16948 36848
rect 17000 36836 17006 36848
rect 17129 36839 17187 36845
rect 17129 36836 17141 36839
rect 17000 36808 17141 36836
rect 17000 36796 17006 36808
rect 17129 36805 17141 36808
rect 17175 36805 17187 36839
rect 17129 36799 17187 36805
rect 17236 36808 24072 36836
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36737 2835 36771
rect 2777 36731 2835 36737
rect 2958 36728 2964 36780
rect 3016 36768 3022 36780
rect 3237 36771 3295 36777
rect 3237 36768 3249 36771
rect 3016 36740 3249 36768
rect 3016 36728 3022 36740
rect 3237 36737 3249 36740
rect 3283 36737 3295 36771
rect 3237 36731 3295 36737
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36768 4307 36771
rect 4614 36768 4620 36780
rect 4295 36740 4620 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 4985 36771 5043 36777
rect 4985 36737 4997 36771
rect 5031 36768 5043 36771
rect 5350 36768 5356 36780
rect 5031 36740 5356 36768
rect 5031 36737 5043 36740
rect 4985 36731 5043 36737
rect 5350 36728 5356 36740
rect 5408 36728 5414 36780
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 5534 36768 5540 36780
rect 5491 36740 5540 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 5534 36728 5540 36740
rect 5592 36728 5598 36780
rect 5626 36728 5632 36780
rect 5684 36768 5690 36780
rect 6178 36768 6184 36780
rect 5684 36740 6184 36768
rect 5684 36728 5690 36740
rect 6178 36728 6184 36740
rect 6236 36768 6242 36780
rect 6457 36771 6515 36777
rect 6457 36768 6469 36771
rect 6236 36740 6469 36768
rect 6236 36728 6242 36740
rect 6457 36737 6469 36740
rect 6503 36737 6515 36771
rect 7098 36768 7104 36780
rect 7059 36740 7104 36768
rect 6457 36731 6515 36737
rect 7098 36728 7104 36740
rect 7156 36728 7162 36780
rect 7926 36728 7932 36780
rect 7984 36768 7990 36780
rect 8113 36771 8171 36777
rect 8113 36768 8125 36771
rect 7984 36740 8125 36768
rect 7984 36728 7990 36740
rect 8113 36737 8125 36740
rect 8159 36737 8171 36771
rect 8570 36768 8576 36780
rect 8531 36740 8576 36768
rect 8113 36731 8171 36737
rect 8570 36728 8576 36740
rect 8628 36728 8634 36780
rect 9585 36771 9643 36777
rect 9585 36737 9597 36771
rect 9631 36768 9643 36771
rect 9674 36768 9680 36780
rect 9631 36740 9680 36768
rect 9631 36737 9643 36740
rect 9585 36731 9643 36737
rect 9674 36728 9680 36740
rect 9732 36728 9738 36780
rect 10686 36768 10692 36780
rect 10647 36740 10692 36768
rect 10686 36728 10692 36740
rect 10744 36728 10750 36780
rect 12345 36771 12403 36777
rect 12345 36737 12357 36771
rect 12391 36768 12403 36771
rect 12526 36768 12532 36780
rect 12391 36740 12532 36768
rect 12391 36737 12403 36740
rect 12345 36731 12403 36737
rect 12526 36728 12532 36740
rect 12584 36728 12590 36780
rect 13817 36771 13875 36777
rect 13817 36737 13829 36771
rect 13863 36737 13875 36771
rect 14274 36768 14280 36780
rect 14235 36740 14280 36768
rect 13817 36731 13875 36737
rect 9398 36660 9404 36712
rect 9456 36700 9462 36712
rect 11517 36703 11575 36709
rect 11517 36700 11529 36703
rect 9456 36672 11529 36700
rect 9456 36660 9462 36672
rect 11517 36669 11529 36672
rect 11563 36669 11575 36703
rect 13832 36700 13860 36731
rect 14274 36728 14280 36740
rect 14332 36728 14338 36780
rect 15930 36768 15936 36780
rect 15891 36740 15936 36768
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 14826 36700 14832 36712
rect 13832 36672 14832 36700
rect 11517 36663 11575 36669
rect 14826 36660 14832 36672
rect 14884 36660 14890 36712
rect 14918 36660 14924 36712
rect 14976 36700 14982 36712
rect 17236 36700 17264 36808
rect 18049 36771 18107 36777
rect 18049 36737 18061 36771
rect 18095 36737 18107 36771
rect 18782 36768 18788 36780
rect 18743 36740 18788 36768
rect 18049 36731 18107 36737
rect 14976 36672 17264 36700
rect 14976 36660 14982 36672
rect 2038 36632 2044 36644
rect 1999 36604 2044 36632
rect 2038 36592 2044 36604
rect 2096 36592 2102 36644
rect 6638 36632 6644 36644
rect 6599 36604 6644 36632
rect 6638 36592 6644 36604
rect 6696 36592 6702 36644
rect 6914 36592 6920 36644
rect 6972 36632 6978 36644
rect 7929 36635 7987 36641
rect 7929 36632 7941 36635
rect 6972 36604 7941 36632
rect 6972 36592 6978 36604
rect 7929 36601 7941 36604
rect 7975 36601 7987 36635
rect 7929 36595 7987 36601
rect 13081 36635 13139 36641
rect 13081 36601 13093 36635
rect 13127 36632 13139 36635
rect 13262 36632 13268 36644
rect 13127 36604 13268 36632
rect 13127 36601 13139 36604
rect 13081 36595 13139 36601
rect 13262 36592 13268 36604
rect 13320 36592 13326 36644
rect 17310 36632 17316 36644
rect 17271 36604 17316 36632
rect 17310 36592 17316 36604
rect 17368 36592 17374 36644
rect 18064 36632 18092 36731
rect 18782 36728 18788 36740
rect 18840 36728 18846 36780
rect 19705 36771 19763 36777
rect 19705 36737 19717 36771
rect 19751 36768 19763 36771
rect 20254 36768 20260 36780
rect 19751 36740 20260 36768
rect 19751 36737 19763 36740
rect 19705 36731 19763 36737
rect 20254 36728 20260 36740
rect 20312 36728 20318 36780
rect 20441 36771 20499 36777
rect 20441 36737 20453 36771
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 20456 36700 20484 36731
rect 20530 36728 20536 36780
rect 20588 36768 20594 36780
rect 20901 36771 20959 36777
rect 20901 36768 20913 36771
rect 20588 36740 20913 36768
rect 20588 36728 20594 36740
rect 20901 36737 20913 36740
rect 20947 36737 20959 36771
rect 20901 36731 20959 36737
rect 20990 36728 20996 36780
rect 21048 36768 21054 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21048 36740 21833 36768
rect 21048 36728 21054 36740
rect 21821 36737 21833 36740
rect 21867 36737 21879 36771
rect 22554 36768 22560 36780
rect 22515 36740 22560 36768
rect 21821 36731 21879 36737
rect 22554 36728 22560 36740
rect 22612 36728 22618 36780
rect 23198 36728 23204 36780
rect 23256 36768 23262 36780
rect 23474 36768 23480 36780
rect 23256 36740 23480 36768
rect 23256 36728 23262 36740
rect 23474 36728 23480 36740
rect 23532 36768 23538 36780
rect 24044 36777 24072 36808
rect 24118 36796 24124 36848
rect 24176 36836 24182 36848
rect 31110 36836 31116 36848
rect 24176 36808 31116 36836
rect 24176 36796 24182 36808
rect 31110 36796 31116 36808
rect 31168 36796 31174 36848
rect 34882 36796 34888 36848
rect 34940 36836 34946 36848
rect 35710 36836 35716 36848
rect 34940 36808 35716 36836
rect 34940 36796 34946 36808
rect 35710 36796 35716 36808
rect 35768 36836 35774 36848
rect 37277 36839 37335 36845
rect 37277 36836 37289 36839
rect 35768 36808 37289 36836
rect 35768 36796 35774 36808
rect 37277 36805 37289 36808
rect 37323 36805 37335 36839
rect 37277 36799 37335 36805
rect 37921 36839 37979 36845
rect 37921 36805 37933 36839
rect 37967 36836 37979 36839
rect 38010 36836 38016 36848
rect 37967 36808 38016 36836
rect 37967 36805 37979 36808
rect 37921 36799 37979 36805
rect 38010 36796 38016 36808
rect 38068 36796 38074 36848
rect 23569 36771 23627 36777
rect 23569 36768 23581 36771
rect 23532 36740 23581 36768
rect 23532 36728 23538 36740
rect 23569 36737 23581 36740
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 24029 36771 24087 36777
rect 24029 36737 24041 36771
rect 24075 36737 24087 36771
rect 24029 36731 24087 36737
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36737 24823 36771
rect 24765 36731 24823 36737
rect 21082 36700 21088 36712
rect 20456 36672 21088 36700
rect 21082 36660 21088 36672
rect 21140 36660 21146 36712
rect 21174 36660 21180 36712
rect 21232 36700 21238 36712
rect 24780 36700 24808 36731
rect 25406 36728 25412 36780
rect 25464 36768 25470 36780
rect 25501 36771 25559 36777
rect 25501 36768 25513 36771
rect 25464 36740 25513 36768
rect 25464 36728 25470 36740
rect 25501 36737 25513 36740
rect 25547 36737 25559 36771
rect 26418 36768 26424 36780
rect 26379 36740 26424 36768
rect 25501 36731 25559 36737
rect 26418 36728 26424 36740
rect 26476 36728 26482 36780
rect 26878 36728 26884 36780
rect 26936 36768 26942 36780
rect 26973 36771 27031 36777
rect 26973 36768 26985 36771
rect 26936 36740 26985 36768
rect 26936 36728 26942 36740
rect 26973 36737 26985 36740
rect 27019 36737 27031 36771
rect 26973 36731 27031 36737
rect 27246 36728 27252 36780
rect 27304 36768 27310 36780
rect 27709 36771 27767 36777
rect 27709 36768 27721 36771
rect 27304 36740 27721 36768
rect 27304 36728 27310 36740
rect 27709 36737 27721 36740
rect 27755 36737 27767 36771
rect 27709 36731 27767 36737
rect 28626 36728 28632 36780
rect 28684 36768 28690 36780
rect 28721 36771 28779 36777
rect 28721 36768 28733 36771
rect 28684 36740 28733 36768
rect 28684 36728 28690 36740
rect 28721 36737 28733 36740
rect 28767 36737 28779 36771
rect 29270 36768 29276 36780
rect 29231 36740 29276 36768
rect 28721 36731 28779 36737
rect 29270 36728 29276 36740
rect 29328 36728 29334 36780
rect 30006 36768 30012 36780
rect 29967 36740 30012 36768
rect 30006 36728 30012 36740
rect 30064 36728 30070 36780
rect 31018 36768 31024 36780
rect 30979 36740 31024 36768
rect 31018 36728 31024 36740
rect 31076 36728 31082 36780
rect 31938 36728 31944 36780
rect 31996 36768 32002 36780
rect 32125 36771 32183 36777
rect 32125 36768 32137 36771
rect 31996 36740 32137 36768
rect 31996 36728 32002 36740
rect 32125 36737 32137 36740
rect 32171 36737 32183 36771
rect 33134 36768 33140 36780
rect 33095 36740 33140 36768
rect 32125 36731 32183 36737
rect 33134 36728 33140 36740
rect 33192 36728 33198 36780
rect 34238 36768 34244 36780
rect 34199 36740 34244 36768
rect 34238 36728 34244 36740
rect 34296 36728 34302 36780
rect 34514 36728 34520 36780
rect 34572 36768 34578 36780
rect 35253 36771 35311 36777
rect 35253 36768 35265 36771
rect 34572 36740 35265 36768
rect 34572 36728 34578 36740
rect 35253 36737 35265 36740
rect 35299 36737 35311 36771
rect 35253 36731 35311 36737
rect 36262 36728 36268 36780
rect 36320 36768 36326 36780
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 36320 36740 36369 36768
rect 36320 36728 36326 36740
rect 36357 36737 36369 36740
rect 36403 36737 36415 36771
rect 36357 36731 36415 36737
rect 21232 36672 24808 36700
rect 21232 36660 21238 36672
rect 24854 36660 24860 36712
rect 24912 36700 24918 36712
rect 37550 36700 37556 36712
rect 24912 36672 37556 36700
rect 24912 36660 24918 36672
rect 37550 36660 37556 36672
rect 37608 36660 37614 36712
rect 18598 36632 18604 36644
rect 18064 36604 18604 36632
rect 18598 36592 18604 36604
rect 18656 36632 18662 36644
rect 18656 36604 23520 36632
rect 18656 36592 18662 36604
rect 1486 36524 1492 36576
rect 1544 36564 1550 36576
rect 2593 36567 2651 36573
rect 2593 36564 2605 36567
rect 1544 36536 2605 36564
rect 1544 36524 1550 36536
rect 2593 36533 2605 36536
rect 2639 36533 2651 36567
rect 2593 36527 2651 36533
rect 6362 36524 6368 36576
rect 6420 36564 6426 36576
rect 6730 36564 6736 36576
rect 6420 36536 6736 36564
rect 6420 36524 6426 36536
rect 6730 36524 6736 36536
rect 6788 36524 6794 36576
rect 23382 36564 23388 36576
rect 23343 36536 23388 36564
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 23492 36564 23520 36604
rect 23658 36592 23664 36644
rect 23716 36632 23722 36644
rect 23716 36604 24808 36632
rect 23716 36592 23722 36604
rect 24670 36564 24676 36576
rect 23492 36536 24676 36564
rect 24670 36524 24676 36536
rect 24728 36524 24734 36576
rect 24780 36564 24808 36604
rect 26326 36592 26332 36644
rect 26384 36632 26390 36644
rect 27157 36635 27215 36641
rect 27157 36632 27169 36635
rect 26384 36604 27169 36632
rect 26384 36592 26390 36604
rect 27157 36601 27169 36604
rect 27203 36601 27215 36635
rect 27157 36595 27215 36601
rect 38105 36635 38163 36641
rect 38105 36601 38117 36635
rect 38151 36632 38163 36635
rect 38194 36632 38200 36644
rect 38151 36604 38200 36632
rect 38151 36601 38163 36604
rect 38105 36595 38163 36601
rect 38194 36592 38200 36604
rect 38252 36592 38258 36644
rect 26237 36567 26295 36573
rect 26237 36564 26249 36567
rect 24780 36536 26249 36564
rect 26237 36533 26249 36536
rect 26283 36533 26295 36567
rect 26237 36527 26295 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 382 36320 388 36372
rect 440 36360 446 36372
rect 1489 36363 1547 36369
rect 1489 36360 1501 36363
rect 440 36332 1501 36360
rect 440 36320 446 36332
rect 1489 36329 1501 36332
rect 1535 36329 1547 36363
rect 1489 36323 1547 36329
rect 1854 36320 1860 36372
rect 1912 36360 1918 36372
rect 2225 36363 2283 36369
rect 2225 36360 2237 36363
rect 1912 36332 2237 36360
rect 1912 36320 1918 36332
rect 2225 36329 2237 36332
rect 2271 36329 2283 36363
rect 2225 36323 2283 36329
rect 2866 36320 2872 36372
rect 2924 36360 2930 36372
rect 3053 36363 3111 36369
rect 3053 36360 3065 36363
rect 2924 36332 3065 36360
rect 2924 36320 2930 36332
rect 3053 36329 3065 36332
rect 3099 36329 3111 36363
rect 3053 36323 3111 36329
rect 3878 36320 3884 36372
rect 3936 36360 3942 36372
rect 4065 36363 4123 36369
rect 4065 36360 4077 36363
rect 3936 36332 4077 36360
rect 3936 36320 3942 36332
rect 4065 36329 4077 36332
rect 4111 36329 4123 36363
rect 5350 36360 5356 36372
rect 5311 36332 5356 36360
rect 4065 36323 4123 36329
rect 5350 36320 5356 36332
rect 5408 36320 5414 36372
rect 5994 36320 6000 36372
rect 6052 36360 6058 36372
rect 6181 36363 6239 36369
rect 6181 36360 6193 36363
rect 6052 36332 6193 36360
rect 6052 36320 6058 36332
rect 6181 36329 6193 36332
rect 6227 36329 6239 36363
rect 6181 36323 6239 36329
rect 7190 36320 7196 36372
rect 7248 36360 7254 36372
rect 7285 36363 7343 36369
rect 7285 36360 7297 36363
rect 7248 36332 7297 36360
rect 7248 36320 7254 36332
rect 7285 36329 7297 36332
rect 7331 36329 7343 36363
rect 7926 36360 7932 36372
rect 7887 36332 7932 36360
rect 7285 36323 7343 36329
rect 7926 36320 7932 36332
rect 7984 36320 7990 36372
rect 8294 36320 8300 36372
rect 8352 36360 8358 36372
rect 9033 36363 9091 36369
rect 9033 36360 9045 36363
rect 8352 36332 9045 36360
rect 8352 36320 8358 36332
rect 9033 36329 9045 36332
rect 9079 36329 9091 36363
rect 9033 36323 9091 36329
rect 9858 36320 9864 36372
rect 9916 36360 9922 36372
rect 10045 36363 10103 36369
rect 10045 36360 10057 36363
rect 9916 36332 10057 36360
rect 9916 36320 9922 36332
rect 10045 36329 10057 36332
rect 10091 36329 10103 36363
rect 10045 36323 10103 36329
rect 10226 36320 10232 36372
rect 10284 36360 10290 36372
rect 10781 36363 10839 36369
rect 10781 36360 10793 36363
rect 10284 36332 10793 36360
rect 10284 36320 10290 36332
rect 10781 36329 10793 36332
rect 10827 36329 10839 36363
rect 10781 36323 10839 36329
rect 11330 36320 11336 36372
rect 11388 36360 11394 36372
rect 11517 36363 11575 36369
rect 11517 36360 11529 36363
rect 11388 36332 11529 36360
rect 11388 36320 11394 36332
rect 11517 36329 11529 36332
rect 11563 36329 11575 36363
rect 11517 36323 11575 36329
rect 12434 36320 12440 36372
rect 12492 36360 12498 36372
rect 12529 36363 12587 36369
rect 12529 36360 12541 36363
rect 12492 36332 12541 36360
rect 12492 36320 12498 36332
rect 12529 36329 12541 36332
rect 12575 36329 12587 36363
rect 12529 36323 12587 36329
rect 13446 36320 13452 36372
rect 13504 36360 13510 36372
rect 14277 36363 14335 36369
rect 14277 36360 14289 36363
rect 13504 36332 14289 36360
rect 13504 36320 13510 36332
rect 14277 36329 14289 36332
rect 14323 36329 14335 36363
rect 14277 36323 14335 36329
rect 14458 36320 14464 36372
rect 14516 36360 14522 36372
rect 15197 36363 15255 36369
rect 15197 36360 15209 36363
rect 14516 36332 15209 36360
rect 14516 36320 14522 36332
rect 15197 36329 15209 36332
rect 15243 36329 15255 36363
rect 15197 36323 15255 36329
rect 15933 36363 15991 36369
rect 15933 36329 15945 36363
rect 15979 36360 15991 36363
rect 16206 36360 16212 36372
rect 15979 36332 16212 36360
rect 15979 36329 15991 36332
rect 15933 36323 15991 36329
rect 16206 36320 16212 36332
rect 16264 36320 16270 36372
rect 16574 36320 16580 36372
rect 16632 36360 16638 36372
rect 16761 36363 16819 36369
rect 16761 36360 16773 36363
rect 16632 36332 16773 36360
rect 16632 36320 16638 36332
rect 16761 36329 16773 36332
rect 16807 36329 16819 36363
rect 16761 36323 16819 36329
rect 17586 36320 17592 36372
rect 17644 36360 17650 36372
rect 17773 36363 17831 36369
rect 17773 36360 17785 36363
rect 17644 36332 17785 36360
rect 17644 36320 17650 36332
rect 17773 36329 17785 36332
rect 17819 36329 17831 36363
rect 17773 36323 17831 36329
rect 18690 36320 18696 36372
rect 18748 36360 18754 36372
rect 19337 36363 19395 36369
rect 19337 36360 19349 36363
rect 18748 36332 19349 36360
rect 18748 36320 18754 36332
rect 19337 36329 19349 36332
rect 19383 36329 19395 36363
rect 19337 36323 19395 36329
rect 20165 36363 20223 36369
rect 20165 36329 20177 36363
rect 20211 36360 20223 36363
rect 20530 36360 20536 36372
rect 20211 36332 20536 36360
rect 20211 36329 20223 36332
rect 20165 36323 20223 36329
rect 20530 36320 20536 36332
rect 20588 36320 20594 36372
rect 20809 36363 20867 36369
rect 20809 36329 20821 36363
rect 20855 36360 20867 36363
rect 20990 36360 20996 36372
rect 20855 36332 20996 36360
rect 20855 36329 20867 36332
rect 20809 36323 20867 36329
rect 20990 36320 20996 36332
rect 21048 36320 21054 36372
rect 21729 36363 21787 36369
rect 21729 36329 21741 36363
rect 21775 36360 21787 36363
rect 21818 36360 21824 36372
rect 21775 36332 21824 36360
rect 21775 36329 21787 36332
rect 21729 36323 21787 36329
rect 21818 36320 21824 36332
rect 21876 36320 21882 36372
rect 22066 36332 23796 36360
rect 13541 36295 13599 36301
rect 13541 36261 13553 36295
rect 13587 36292 13599 36295
rect 14918 36292 14924 36304
rect 13587 36264 14924 36292
rect 13587 36261 13599 36264
rect 13541 36255 13599 36261
rect 14918 36252 14924 36264
rect 14976 36252 14982 36304
rect 15102 36252 15108 36304
rect 15160 36292 15166 36304
rect 18417 36295 18475 36301
rect 18417 36292 18429 36295
rect 15160 36264 18429 36292
rect 15160 36252 15166 36264
rect 18417 36261 18429 36264
rect 18463 36261 18475 36295
rect 18417 36255 18475 36261
rect 12894 36224 12900 36236
rect 12728 36196 12900 36224
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 2409 36159 2467 36165
rect 2409 36125 2421 36159
rect 2455 36125 2467 36159
rect 3234 36156 3240 36168
rect 3195 36128 3240 36156
rect 2409 36119 2467 36125
rect 2424 36088 2452 36119
rect 3234 36116 3240 36128
rect 3292 36116 3298 36168
rect 4249 36159 4307 36165
rect 4249 36125 4261 36159
rect 4295 36156 4307 36159
rect 4706 36156 4712 36168
rect 4295 36128 4712 36156
rect 4295 36125 4307 36128
rect 4249 36119 4307 36125
rect 4706 36116 4712 36128
rect 4764 36116 4770 36168
rect 5537 36159 5595 36165
rect 5537 36125 5549 36159
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 6365 36159 6423 36165
rect 6365 36125 6377 36159
rect 6411 36156 6423 36159
rect 7006 36156 7012 36168
rect 6411 36128 7012 36156
rect 6411 36125 6423 36128
rect 6365 36119 6423 36125
rect 3142 36088 3148 36100
rect 2424 36060 3148 36088
rect 3142 36048 3148 36060
rect 3200 36048 3206 36100
rect 4893 36091 4951 36097
rect 4893 36057 4905 36091
rect 4939 36088 4951 36091
rect 5552 36088 5580 36119
rect 7006 36116 7012 36128
rect 7064 36116 7070 36168
rect 7466 36156 7472 36168
rect 7427 36128 7472 36156
rect 7466 36116 7472 36128
rect 7524 36116 7530 36168
rect 8018 36116 8024 36168
rect 8076 36156 8082 36168
rect 8113 36159 8171 36165
rect 8113 36156 8125 36159
rect 8076 36128 8125 36156
rect 8076 36116 8082 36128
rect 8113 36125 8125 36128
rect 8159 36125 8171 36159
rect 9214 36156 9220 36168
rect 9175 36128 9220 36156
rect 8113 36119 8171 36125
rect 9214 36116 9220 36128
rect 9272 36116 9278 36168
rect 10226 36156 10232 36168
rect 10187 36128 10232 36156
rect 10226 36116 10232 36128
rect 10284 36116 10290 36168
rect 10965 36159 11023 36165
rect 10965 36125 10977 36159
rect 11011 36125 11023 36159
rect 11698 36156 11704 36168
rect 11659 36128 11704 36156
rect 10965 36119 11023 36125
rect 6454 36088 6460 36100
rect 4939 36060 6460 36088
rect 4939 36057 4951 36060
rect 4893 36051 4951 36057
rect 6454 36048 6460 36060
rect 6512 36048 6518 36100
rect 10980 36088 11008 36119
rect 11698 36116 11704 36128
rect 11756 36116 11762 36168
rect 12728 36165 12756 36196
rect 12894 36184 12900 36196
rect 12952 36224 12958 36236
rect 22066 36224 22094 36332
rect 22741 36295 22799 36301
rect 22741 36261 22753 36295
rect 22787 36261 22799 36295
rect 23658 36292 23664 36304
rect 23619 36264 23664 36292
rect 22741 36255 22799 36261
rect 12952 36196 22094 36224
rect 22756 36224 22784 36255
rect 23658 36252 23664 36264
rect 23716 36252 23722 36304
rect 23768 36292 23796 36332
rect 23934 36320 23940 36372
rect 23992 36360 23998 36372
rect 24489 36363 24547 36369
rect 24489 36360 24501 36363
rect 23992 36332 24501 36360
rect 23992 36320 23998 36332
rect 24489 36329 24501 36332
rect 24535 36329 24547 36363
rect 25314 36360 25320 36372
rect 25275 36332 25320 36360
rect 24489 36323 24547 36329
rect 25314 36320 25320 36332
rect 25372 36320 25378 36372
rect 26326 36360 26332 36372
rect 25424 36332 26332 36360
rect 25424 36292 25452 36332
rect 26326 36320 26332 36332
rect 26384 36320 26390 36372
rect 26602 36360 26608 36372
rect 26563 36332 26608 36360
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 27246 36360 27252 36372
rect 27207 36332 27252 36360
rect 27246 36320 27252 36332
rect 27304 36320 27310 36372
rect 28626 36360 28632 36372
rect 28587 36332 28632 36360
rect 28626 36320 28632 36332
rect 28684 36320 28690 36372
rect 28810 36320 28816 36372
rect 28868 36360 28874 36372
rect 29549 36363 29607 36369
rect 29549 36360 29561 36363
rect 28868 36332 29561 36360
rect 28868 36320 28874 36332
rect 29549 36329 29561 36332
rect 29595 36329 29607 36363
rect 29549 36323 29607 36329
rect 31294 36320 31300 36372
rect 31352 36360 31358 36372
rect 31849 36363 31907 36369
rect 31849 36360 31861 36363
rect 31352 36332 31861 36360
rect 31352 36320 31358 36332
rect 31849 36329 31861 36332
rect 31895 36329 31907 36363
rect 31849 36323 31907 36329
rect 34422 36320 34428 36372
rect 34480 36360 34486 36372
rect 34885 36363 34943 36369
rect 34885 36360 34897 36363
rect 34480 36332 34897 36360
rect 34480 36320 34486 36332
rect 34885 36329 34897 36332
rect 34931 36329 34943 36363
rect 35434 36360 35440 36372
rect 35395 36332 35440 36360
rect 34885 36323 34943 36329
rect 35434 36320 35440 36332
rect 35492 36320 35498 36372
rect 23768 36264 25452 36292
rect 25961 36295 26019 36301
rect 25961 36261 25973 36295
rect 26007 36292 26019 36295
rect 26418 36292 26424 36304
rect 26007 36264 26424 36292
rect 26007 36261 26019 36264
rect 25961 36255 26019 36261
rect 26418 36252 26424 36264
rect 26476 36252 26482 36304
rect 28169 36295 28227 36301
rect 28169 36261 28181 36295
rect 28215 36292 28227 36295
rect 29270 36292 29276 36304
rect 28215 36264 29276 36292
rect 28215 36261 28227 36264
rect 28169 36255 28227 36261
rect 29270 36252 29276 36264
rect 29328 36252 29334 36304
rect 29362 36252 29368 36304
rect 29420 36292 29426 36304
rect 32401 36295 32459 36301
rect 32401 36292 32413 36295
rect 29420 36264 32413 36292
rect 29420 36252 29426 36264
rect 32401 36261 32413 36264
rect 32447 36261 32459 36295
rect 32401 36255 32459 36261
rect 28442 36224 28448 36236
rect 22756 36196 28448 36224
rect 12952 36184 12958 36196
rect 28442 36184 28448 36196
rect 28500 36184 28506 36236
rect 30929 36227 30987 36233
rect 30929 36224 30941 36227
rect 28644 36196 30941 36224
rect 12713 36159 12771 36165
rect 12713 36125 12725 36159
rect 12759 36125 12771 36159
rect 12713 36119 12771 36125
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36156 13415 36159
rect 13446 36156 13452 36168
rect 13403 36128 13452 36156
rect 13403 36125 13415 36128
rect 13357 36119 13415 36125
rect 13446 36116 13452 36128
rect 13504 36116 13510 36168
rect 13906 36116 13912 36168
rect 13964 36156 13970 36168
rect 14093 36159 14151 36165
rect 14093 36156 14105 36159
rect 13964 36128 14105 36156
rect 13964 36116 13970 36128
rect 14093 36125 14105 36128
rect 14139 36125 14151 36159
rect 14093 36119 14151 36125
rect 14182 36116 14188 36168
rect 14240 36156 14246 36168
rect 15013 36159 15071 36165
rect 15013 36156 15025 36159
rect 14240 36128 15025 36156
rect 14240 36116 14246 36128
rect 15013 36125 15025 36128
rect 15059 36125 15071 36159
rect 15013 36119 15071 36125
rect 16117 36159 16175 36165
rect 16117 36125 16129 36159
rect 16163 36156 16175 36159
rect 16482 36156 16488 36168
rect 16163 36128 16488 36156
rect 16163 36125 16175 36128
rect 16117 36119 16175 36125
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 16945 36159 17003 36165
rect 16945 36125 16957 36159
rect 16991 36156 17003 36159
rect 17126 36156 17132 36168
rect 16991 36128 17132 36156
rect 16991 36125 17003 36128
rect 16945 36119 17003 36125
rect 17126 36116 17132 36128
rect 17184 36116 17190 36168
rect 17957 36159 18015 36165
rect 17957 36125 17969 36159
rect 18003 36156 18015 36159
rect 18046 36156 18052 36168
rect 18003 36128 18052 36156
rect 18003 36125 18015 36128
rect 17957 36119 18015 36125
rect 18046 36116 18052 36128
rect 18104 36116 18110 36168
rect 19521 36159 19579 36165
rect 19521 36125 19533 36159
rect 19567 36125 19579 36159
rect 19521 36119 19579 36125
rect 19981 36159 20039 36165
rect 19981 36125 19993 36159
rect 20027 36156 20039 36159
rect 20162 36156 20168 36168
rect 20027 36128 20168 36156
rect 20027 36125 20039 36128
rect 19981 36119 20039 36125
rect 12066 36088 12072 36100
rect 10980 36060 12072 36088
rect 12066 36048 12072 36060
rect 12124 36048 12130 36100
rect 19536 36088 19564 36119
rect 20162 36116 20168 36128
rect 20220 36116 20226 36168
rect 20625 36159 20683 36165
rect 20625 36125 20637 36159
rect 20671 36156 20683 36159
rect 20714 36156 20720 36168
rect 20671 36128 20720 36156
rect 20671 36125 20683 36128
rect 20625 36119 20683 36125
rect 20714 36116 20720 36128
rect 20772 36116 20778 36168
rect 21913 36159 21971 36165
rect 21913 36125 21925 36159
rect 21959 36156 21971 36159
rect 22002 36156 22008 36168
rect 21959 36128 22008 36156
rect 21959 36125 21971 36128
rect 21913 36119 21971 36125
rect 22002 36116 22008 36128
rect 22060 36116 22066 36168
rect 24673 36159 24731 36165
rect 24673 36125 24685 36159
rect 24719 36156 24731 36159
rect 24854 36156 24860 36168
rect 24719 36128 24860 36156
rect 24719 36125 24731 36128
rect 24673 36119 24731 36125
rect 24854 36116 24860 36128
rect 24912 36116 24918 36168
rect 26421 36159 26479 36165
rect 26421 36125 26433 36159
rect 26467 36156 26479 36159
rect 26510 36156 26516 36168
rect 26467 36128 26516 36156
rect 26467 36125 26479 36128
rect 26421 36119 26479 36125
rect 26510 36116 26516 36128
rect 26568 36116 26574 36168
rect 27062 36156 27068 36168
rect 27023 36128 27068 36156
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 27982 36156 27988 36168
rect 27943 36128 27988 36156
rect 27982 36116 27988 36128
rect 28040 36116 28046 36168
rect 20438 36088 20444 36100
rect 19536 36060 20444 36088
rect 20438 36048 20444 36060
rect 20496 36048 20502 36100
rect 22373 36091 22431 36097
rect 22373 36057 22385 36091
rect 22419 36088 22431 36091
rect 23290 36088 23296 36100
rect 22419 36060 23296 36088
rect 22419 36057 22431 36060
rect 22373 36051 22431 36057
rect 23290 36048 23296 36060
rect 23348 36048 23354 36100
rect 24946 36048 24952 36100
rect 25004 36088 25010 36100
rect 28644 36088 28672 36196
rect 30929 36193 30941 36196
rect 30975 36193 30987 36227
rect 30929 36187 30987 36193
rect 31110 36184 31116 36236
rect 31168 36224 31174 36236
rect 36541 36227 36599 36233
rect 36541 36224 36553 36227
rect 31168 36196 36553 36224
rect 31168 36184 31174 36196
rect 36541 36193 36553 36196
rect 36587 36193 36599 36227
rect 37550 36224 37556 36236
rect 37511 36196 37556 36224
rect 36541 36187 36599 36193
rect 37550 36184 37556 36196
rect 37608 36184 37614 36236
rect 28810 36156 28816 36168
rect 28771 36128 28816 36156
rect 28810 36116 28816 36128
rect 28868 36116 28874 36168
rect 30190 36156 30196 36168
rect 30151 36128 30196 36156
rect 30190 36116 30196 36128
rect 30248 36116 30254 36168
rect 31662 36156 31668 36168
rect 31623 36128 31668 36156
rect 31662 36116 31668 36128
rect 31720 36116 31726 36168
rect 34698 36156 34704 36168
rect 34659 36128 34704 36156
rect 34698 36116 34704 36128
rect 34756 36116 34762 36168
rect 36817 36159 36875 36165
rect 36817 36125 36829 36159
rect 36863 36125 36875 36159
rect 36817 36119 36875 36125
rect 37277 36159 37335 36165
rect 37277 36125 37289 36159
rect 37323 36156 37335 36159
rect 38562 36156 38568 36168
rect 37323 36128 38568 36156
rect 37323 36125 37335 36128
rect 37277 36119 37335 36125
rect 25004 36060 28672 36088
rect 30377 36091 30435 36097
rect 25004 36048 25010 36060
rect 30377 36057 30389 36091
rect 30423 36088 30435 36091
rect 30466 36088 30472 36100
rect 30423 36060 30472 36088
rect 30423 36057 30435 36060
rect 30377 36051 30435 36057
rect 30466 36048 30472 36060
rect 30524 36048 30530 36100
rect 30926 36048 30932 36100
rect 30984 36088 30990 36100
rect 31113 36091 31171 36097
rect 31113 36088 31125 36091
rect 30984 36060 31125 36088
rect 30984 36048 30990 36060
rect 31113 36057 31125 36060
rect 31159 36057 31171 36091
rect 31113 36051 31171 36057
rect 32585 36091 32643 36097
rect 32585 36057 32597 36091
rect 32631 36088 32643 36091
rect 33226 36088 33232 36100
rect 32631 36060 33232 36088
rect 32631 36057 32643 36060
rect 32585 36051 32643 36057
rect 33226 36048 33232 36060
rect 33284 36048 33290 36100
rect 33505 36091 33563 36097
rect 33505 36057 33517 36091
rect 33551 36088 33563 36091
rect 33962 36088 33968 36100
rect 33551 36060 33968 36088
rect 33551 36057 33563 36060
rect 33505 36051 33563 36057
rect 33962 36048 33968 36060
rect 34020 36088 34026 36100
rect 34057 36091 34115 36097
rect 34057 36088 34069 36091
rect 34020 36060 34069 36088
rect 34020 36048 34026 36060
rect 34057 36057 34069 36060
rect 34103 36057 34115 36091
rect 36832 36088 36860 36119
rect 38562 36116 38568 36128
rect 38620 36116 38626 36168
rect 38838 36088 38844 36100
rect 36832 36060 38844 36088
rect 34057 36051 34115 36057
rect 38838 36048 38844 36060
rect 38896 36048 38902 36100
rect 22830 36020 22836 36032
rect 22791 35992 22836 36020
rect 22830 35980 22836 35992
rect 22888 35980 22894 36032
rect 23658 35980 23664 36032
rect 23716 36020 23722 36032
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 23716 35992 23765 36020
rect 23716 35980 23722 35992
rect 23753 35989 23765 35992
rect 23799 35989 23811 36023
rect 23753 35983 23811 35989
rect 26326 35980 26332 36032
rect 26384 36020 26390 36032
rect 33413 36023 33471 36029
rect 33413 36020 33425 36023
rect 26384 35992 33425 36020
rect 26384 35980 26390 35992
rect 33413 35989 33425 35992
rect 33459 35989 33471 36023
rect 33413 35983 33471 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 750 35776 756 35828
rect 808 35816 814 35828
rect 1489 35819 1547 35825
rect 1489 35816 1501 35819
rect 808 35788 1501 35816
rect 808 35776 814 35788
rect 1489 35785 1501 35788
rect 1535 35785 1547 35819
rect 1489 35779 1547 35785
rect 2685 35819 2743 35825
rect 2685 35785 2697 35819
rect 2731 35785 2743 35819
rect 2685 35779 2743 35785
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 2700 35680 2728 35779
rect 3142 35776 3148 35828
rect 3200 35816 3206 35828
rect 3329 35819 3387 35825
rect 3329 35816 3341 35819
rect 3200 35788 3341 35816
rect 3200 35776 3206 35788
rect 3329 35785 3341 35788
rect 3375 35785 3387 35819
rect 3329 35779 3387 35785
rect 4062 35776 4068 35828
rect 4120 35816 4126 35828
rect 4525 35819 4583 35825
rect 4525 35816 4537 35819
rect 4120 35788 4537 35816
rect 4120 35776 4126 35788
rect 4525 35785 4537 35788
rect 4571 35785 4583 35819
rect 5074 35816 5080 35828
rect 5035 35788 5080 35816
rect 4525 35779 4583 35785
rect 5074 35776 5080 35788
rect 5132 35776 5138 35828
rect 6641 35819 6699 35825
rect 6641 35785 6653 35819
rect 6687 35816 6699 35819
rect 7098 35816 7104 35828
rect 6687 35788 7104 35816
rect 6687 35785 6699 35788
rect 6641 35779 6699 35785
rect 7098 35776 7104 35788
rect 7156 35776 7162 35828
rect 8570 35816 8576 35828
rect 8531 35788 8576 35816
rect 8570 35776 8576 35788
rect 8628 35776 8634 35828
rect 9306 35776 9312 35828
rect 9364 35816 9370 35828
rect 9769 35819 9827 35825
rect 9769 35816 9781 35819
rect 9364 35788 9781 35816
rect 9364 35776 9370 35788
rect 9769 35785 9781 35788
rect 9815 35785 9827 35819
rect 9769 35779 9827 35785
rect 10686 35776 10692 35828
rect 10744 35816 10750 35828
rect 10781 35819 10839 35825
rect 10781 35816 10793 35819
rect 10744 35788 10793 35816
rect 10744 35776 10750 35788
rect 10781 35785 10793 35788
rect 10827 35785 10839 35819
rect 10781 35779 10839 35785
rect 11698 35776 11704 35828
rect 11756 35816 11762 35828
rect 12253 35819 12311 35825
rect 12253 35816 12265 35819
rect 11756 35788 12265 35816
rect 11756 35776 11762 35788
rect 12253 35785 12265 35788
rect 12299 35785 12311 35819
rect 12253 35779 12311 35785
rect 14185 35819 14243 35825
rect 14185 35785 14197 35819
rect 14231 35816 14243 35819
rect 14274 35816 14280 35828
rect 14231 35788 14280 35816
rect 14231 35785 14243 35788
rect 14185 35779 14243 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 14826 35816 14832 35828
rect 14787 35788 14832 35816
rect 14826 35776 14832 35788
rect 14884 35776 14890 35828
rect 15470 35776 15476 35828
rect 15528 35816 15534 35828
rect 15657 35819 15715 35825
rect 15657 35816 15669 35819
rect 15528 35788 15669 35816
rect 15528 35776 15534 35788
rect 15657 35785 15669 35788
rect 15703 35785 15715 35819
rect 15657 35779 15715 35785
rect 15930 35776 15936 35828
rect 15988 35816 15994 35828
rect 16669 35819 16727 35825
rect 16669 35816 16681 35819
rect 15988 35788 16681 35816
rect 15988 35776 15994 35788
rect 16669 35785 16681 35788
rect 16715 35785 16727 35819
rect 16669 35779 16727 35785
rect 19705 35819 19763 35825
rect 19705 35785 19717 35819
rect 19751 35816 19763 35819
rect 20898 35816 20904 35828
rect 19751 35788 20904 35816
rect 19751 35785 19763 35788
rect 19705 35779 19763 35785
rect 20898 35776 20904 35788
rect 20956 35776 20962 35828
rect 22186 35776 22192 35828
rect 22244 35816 22250 35828
rect 22465 35819 22523 35825
rect 22465 35816 22477 35819
rect 22244 35788 22477 35816
rect 22244 35776 22250 35788
rect 22465 35785 22477 35788
rect 22511 35785 22523 35819
rect 22465 35779 22523 35785
rect 22922 35776 22928 35828
rect 22980 35816 22986 35828
rect 23201 35819 23259 35825
rect 23201 35816 23213 35819
rect 22980 35788 23213 35816
rect 22980 35776 22986 35788
rect 23201 35785 23213 35788
rect 23247 35785 23259 35819
rect 23201 35779 23259 35785
rect 23474 35776 23480 35828
rect 23532 35816 23538 35828
rect 23753 35819 23811 35825
rect 23753 35816 23765 35819
rect 23532 35788 23765 35816
rect 23532 35776 23538 35788
rect 23753 35785 23765 35788
rect 23799 35785 23811 35819
rect 24302 35816 24308 35828
rect 24263 35788 24308 35816
rect 23753 35779 23811 35785
rect 24302 35776 24308 35788
rect 24360 35776 24366 35828
rect 26421 35819 26479 35825
rect 26421 35785 26433 35819
rect 26467 35816 26479 35819
rect 26970 35816 26976 35828
rect 26467 35788 26976 35816
rect 26467 35785 26479 35788
rect 26421 35779 26479 35785
rect 26970 35776 26976 35788
rect 27028 35776 27034 35828
rect 28902 35776 28908 35828
rect 28960 35816 28966 35828
rect 29730 35816 29736 35828
rect 28960 35788 29736 35816
rect 28960 35776 28966 35788
rect 29730 35776 29736 35788
rect 29788 35776 29794 35828
rect 30282 35776 30288 35828
rect 30340 35816 30346 35828
rect 30469 35819 30527 35825
rect 30469 35816 30481 35819
rect 30340 35788 30481 35816
rect 30340 35776 30346 35788
rect 30469 35785 30481 35788
rect 30515 35785 30527 35819
rect 31202 35816 31208 35828
rect 31163 35788 31208 35816
rect 30469 35779 30527 35785
rect 31202 35776 31208 35788
rect 31260 35776 31266 35828
rect 33410 35776 33416 35828
rect 33468 35816 33474 35828
rect 34241 35819 34299 35825
rect 34241 35816 34253 35819
rect 33468 35788 34253 35816
rect 33468 35776 33474 35788
rect 34241 35785 34253 35788
rect 34287 35785 34299 35819
rect 34241 35779 34299 35785
rect 35618 35776 35624 35828
rect 35676 35816 35682 35828
rect 35805 35819 35863 35825
rect 35805 35816 35817 35819
rect 35676 35788 35817 35816
rect 35676 35776 35682 35788
rect 35805 35785 35817 35788
rect 35851 35785 35863 35819
rect 37274 35816 37280 35828
rect 37235 35788 37280 35816
rect 35805 35779 35863 35785
rect 37274 35776 37280 35788
rect 37332 35776 37338 35828
rect 22554 35748 22560 35760
rect 11716 35720 22560 35748
rect 1719 35652 2728 35680
rect 2869 35683 2927 35689
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 2869 35649 2881 35683
rect 2915 35649 2927 35683
rect 3510 35680 3516 35692
rect 3471 35652 3516 35680
rect 2869 35643 2927 35649
rect 2225 35615 2283 35621
rect 2225 35581 2237 35615
rect 2271 35612 2283 35615
rect 2884 35612 2912 35643
rect 3510 35640 3516 35652
rect 3568 35680 3574 35692
rect 3973 35683 4031 35689
rect 3973 35680 3985 35683
rect 3568 35652 3985 35680
rect 3568 35640 3574 35652
rect 3973 35649 3985 35652
rect 4019 35649 4031 35683
rect 3973 35643 4031 35649
rect 6457 35683 6515 35689
rect 6457 35649 6469 35683
rect 6503 35680 6515 35683
rect 8757 35683 8815 35689
rect 6503 35652 6914 35680
rect 6503 35649 6515 35652
rect 6457 35643 6515 35649
rect 5166 35612 5172 35624
rect 2271 35584 5172 35612
rect 2271 35581 2283 35584
rect 2225 35575 2283 35581
rect 5166 35572 5172 35584
rect 5224 35572 5230 35624
rect 5718 35476 5724 35488
rect 5679 35448 5724 35476
rect 5718 35436 5724 35448
rect 5776 35436 5782 35488
rect 6886 35476 6914 35652
rect 8757 35649 8769 35683
rect 8803 35680 8815 35683
rect 9030 35680 9036 35692
rect 8803 35652 9036 35680
rect 8803 35649 8815 35652
rect 8757 35643 8815 35649
rect 9030 35640 9036 35652
rect 9088 35640 9094 35692
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35649 10011 35683
rect 10962 35680 10968 35692
rect 10923 35652 10968 35680
rect 9953 35643 10011 35649
rect 9968 35612 9996 35643
rect 10962 35640 10968 35652
rect 11020 35640 11026 35692
rect 11422 35640 11428 35692
rect 11480 35680 11486 35692
rect 11517 35683 11575 35689
rect 11517 35680 11529 35683
rect 11480 35652 11529 35680
rect 11480 35640 11486 35652
rect 11517 35649 11529 35652
rect 11563 35649 11575 35683
rect 11517 35643 11575 35649
rect 11238 35612 11244 35624
rect 9968 35584 11244 35612
rect 11238 35572 11244 35584
rect 11296 35572 11302 35624
rect 11716 35553 11744 35720
rect 22554 35708 22560 35720
rect 22612 35708 22618 35760
rect 27430 35708 27436 35760
rect 27488 35748 27494 35760
rect 29917 35751 29975 35757
rect 27488 35720 28396 35748
rect 27488 35708 27494 35720
rect 12437 35683 12495 35689
rect 12437 35649 12449 35683
rect 12483 35680 12495 35683
rect 14369 35683 14427 35689
rect 12483 35652 13032 35680
rect 12483 35649 12495 35652
rect 12437 35643 12495 35649
rect 13004 35553 13032 35652
rect 14369 35649 14381 35683
rect 14415 35680 14427 35683
rect 14458 35680 14464 35692
rect 14415 35652 14464 35680
rect 14415 35649 14427 35652
rect 14369 35643 14427 35649
rect 14458 35640 14464 35652
rect 14516 35640 14522 35692
rect 14918 35640 14924 35692
rect 14976 35680 14982 35692
rect 15013 35683 15071 35689
rect 15013 35680 15025 35683
rect 14976 35652 15025 35680
rect 14976 35640 14982 35652
rect 15013 35649 15025 35652
rect 15059 35649 15071 35683
rect 15013 35643 15071 35649
rect 15841 35683 15899 35689
rect 15841 35649 15853 35683
rect 15887 35680 15899 35683
rect 16114 35680 16120 35692
rect 15887 35652 16120 35680
rect 15887 35649 15899 35652
rect 15841 35643 15899 35649
rect 16114 35640 16120 35652
rect 16172 35640 16178 35692
rect 16758 35640 16764 35692
rect 16816 35680 16822 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16816 35652 16865 35680
rect 16816 35640 16822 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 17497 35683 17555 35689
rect 17497 35649 17509 35683
rect 17543 35680 17555 35683
rect 17862 35680 17868 35692
rect 17543 35652 17868 35680
rect 17543 35649 17555 35652
rect 17497 35643 17555 35649
rect 17862 35640 17868 35652
rect 17920 35640 17926 35692
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 23014 35680 23020 35692
rect 22975 35652 23020 35680
rect 19521 35643 19579 35649
rect 16574 35572 16580 35624
rect 16632 35612 16638 35624
rect 18969 35615 19027 35621
rect 18969 35612 18981 35615
rect 16632 35584 18981 35612
rect 16632 35572 16638 35584
rect 18969 35581 18981 35584
rect 19015 35612 19027 35615
rect 19536 35612 19564 35643
rect 23014 35640 23020 35652
rect 23072 35640 23078 35692
rect 26237 35683 26295 35689
rect 26237 35649 26249 35683
rect 26283 35680 26295 35683
rect 26326 35680 26332 35692
rect 26283 35652 26332 35680
rect 26283 35649 26295 35652
rect 26237 35643 26295 35649
rect 26326 35640 26332 35652
rect 26384 35640 26390 35692
rect 27522 35680 27528 35692
rect 27483 35652 27528 35680
rect 27522 35640 27528 35652
rect 27580 35640 27586 35692
rect 28368 35689 28396 35720
rect 29917 35717 29929 35751
rect 29963 35748 29975 35751
rect 30558 35748 30564 35760
rect 29963 35720 30564 35748
rect 29963 35717 29975 35720
rect 29917 35711 29975 35717
rect 30558 35708 30564 35720
rect 30616 35708 30622 35760
rect 28353 35683 28411 35689
rect 28353 35649 28365 35683
rect 28399 35680 28411 35683
rect 28813 35683 28871 35689
rect 28813 35680 28825 35683
rect 28399 35652 28825 35680
rect 28399 35649 28411 35652
rect 28353 35643 28411 35649
rect 28813 35649 28825 35652
rect 28859 35649 28871 35683
rect 28813 35643 28871 35649
rect 30653 35683 30711 35689
rect 30653 35649 30665 35683
rect 30699 35680 30711 35683
rect 31294 35680 31300 35692
rect 30699 35652 31300 35680
rect 30699 35649 30711 35652
rect 30653 35643 30711 35649
rect 31294 35640 31300 35652
rect 31352 35640 31358 35692
rect 32769 35683 32827 35689
rect 32769 35649 32781 35683
rect 32815 35680 32827 35683
rect 32950 35680 32956 35692
rect 32815 35652 32956 35680
rect 32815 35649 32827 35652
rect 32769 35643 32827 35649
rect 32950 35640 32956 35652
rect 33008 35640 33014 35692
rect 33597 35683 33655 35689
rect 33597 35649 33609 35683
rect 33643 35680 33655 35683
rect 33686 35680 33692 35692
rect 33643 35652 33692 35680
rect 33643 35649 33655 35652
rect 33597 35643 33655 35649
rect 33686 35640 33692 35652
rect 33744 35640 33750 35692
rect 33870 35640 33876 35692
rect 33928 35680 33934 35692
rect 34057 35683 34115 35689
rect 34057 35680 34069 35683
rect 33928 35652 34069 35680
rect 33928 35640 33934 35652
rect 34057 35649 34069 35652
rect 34103 35649 34115 35683
rect 34057 35643 34115 35649
rect 35161 35683 35219 35689
rect 35161 35649 35173 35683
rect 35207 35680 35219 35683
rect 35342 35680 35348 35692
rect 35207 35652 35348 35680
rect 35207 35649 35219 35652
rect 35161 35643 35219 35649
rect 35342 35640 35348 35652
rect 35400 35640 35406 35692
rect 35618 35680 35624 35692
rect 35579 35652 35624 35680
rect 35618 35640 35624 35652
rect 35676 35640 35682 35692
rect 36354 35640 36360 35692
rect 36412 35680 36418 35692
rect 36449 35683 36507 35689
rect 36449 35680 36461 35683
rect 36412 35652 36461 35680
rect 36412 35640 36418 35652
rect 36449 35649 36461 35652
rect 36495 35649 36507 35683
rect 36449 35643 36507 35649
rect 37918 35640 37924 35692
rect 37976 35680 37982 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37976 35652 38025 35680
rect 37976 35640 37982 35652
rect 38013 35649 38025 35652
rect 38059 35680 38071 35683
rect 39022 35680 39028 35692
rect 38059 35652 39028 35680
rect 38059 35649 38071 35652
rect 38013 35643 38071 35649
rect 39022 35640 39028 35652
rect 39080 35640 39086 35692
rect 19015 35584 19564 35612
rect 19015 35581 19027 35584
rect 18969 35575 19027 35581
rect 11701 35547 11759 35553
rect 11701 35513 11713 35547
rect 11747 35513 11759 35547
rect 11701 35507 11759 35513
rect 12989 35547 13047 35553
rect 12989 35513 13001 35547
rect 13035 35544 13047 35547
rect 13354 35544 13360 35556
rect 13035 35516 13360 35544
rect 13035 35513 13047 35516
rect 12989 35507 13047 35513
rect 13354 35504 13360 35516
rect 13412 35504 13418 35556
rect 16482 35504 16488 35556
rect 16540 35544 16546 35556
rect 17313 35547 17371 35553
rect 17313 35544 17325 35547
rect 16540 35516 17325 35544
rect 16540 35504 16546 35516
rect 17313 35513 17325 35516
rect 17359 35513 17371 35547
rect 17313 35507 17371 35513
rect 27709 35547 27767 35553
rect 27709 35513 27721 35547
rect 27755 35544 27767 35547
rect 29546 35544 29552 35556
rect 27755 35516 29552 35544
rect 27755 35513 27767 35516
rect 27709 35507 27767 35513
rect 29546 35504 29552 35516
rect 29604 35504 29610 35556
rect 32398 35504 32404 35556
rect 32456 35544 32462 35556
rect 33413 35547 33471 35553
rect 33413 35544 33425 35547
rect 32456 35516 33425 35544
rect 32456 35504 32462 35516
rect 33413 35513 33425 35516
rect 33459 35513 33471 35547
rect 33413 35507 33471 35513
rect 34977 35547 35035 35553
rect 34977 35513 34989 35547
rect 35023 35544 35035 35547
rect 36538 35544 36544 35556
rect 35023 35516 36544 35544
rect 35023 35513 35035 35516
rect 34977 35507 35035 35513
rect 36538 35504 36544 35516
rect 36596 35504 36602 35556
rect 36633 35547 36691 35553
rect 36633 35513 36645 35547
rect 36679 35544 36691 35547
rect 37366 35544 37372 35556
rect 36679 35516 37372 35544
rect 36679 35513 36691 35516
rect 36633 35507 36691 35513
rect 37366 35504 37372 35516
rect 37424 35504 37430 35556
rect 37826 35544 37832 35556
rect 37787 35516 37832 35544
rect 37826 35504 37832 35516
rect 37884 35504 37890 35556
rect 7193 35479 7251 35485
rect 7193 35476 7205 35479
rect 6886 35448 7205 35476
rect 7193 35445 7205 35448
rect 7239 35476 7251 35479
rect 7742 35476 7748 35488
rect 7239 35448 7748 35476
rect 7239 35445 7251 35448
rect 7193 35439 7251 35445
rect 7742 35436 7748 35448
rect 7800 35436 7806 35488
rect 8110 35476 8116 35488
rect 8071 35448 8116 35476
rect 8110 35436 8116 35448
rect 8168 35436 8174 35488
rect 13446 35476 13452 35488
rect 13407 35448 13452 35476
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 17862 35436 17868 35488
rect 17920 35476 17926 35488
rect 17957 35479 18015 35485
rect 17957 35476 17969 35479
rect 17920 35448 17969 35476
rect 17920 35436 17926 35448
rect 17957 35445 17969 35448
rect 18003 35445 18015 35479
rect 20162 35476 20168 35488
rect 20123 35448 20168 35476
rect 17957 35439 18015 35445
rect 20162 35436 20168 35448
rect 20220 35436 20226 35488
rect 20714 35476 20720 35488
rect 20675 35448 20720 35476
rect 20714 35436 20720 35448
rect 20772 35436 20778 35488
rect 22002 35476 22008 35488
rect 21963 35448 22008 35476
rect 22002 35436 22008 35448
rect 22060 35436 22066 35488
rect 24854 35476 24860 35488
rect 24815 35448 24860 35476
rect 24854 35436 24860 35448
rect 24912 35436 24918 35488
rect 25406 35476 25412 35488
rect 25367 35448 25412 35476
rect 25406 35436 25412 35448
rect 25464 35436 25470 35488
rect 26970 35476 26976 35488
rect 26931 35448 26976 35476
rect 26970 35436 26976 35448
rect 27028 35436 27034 35488
rect 28166 35476 28172 35488
rect 28127 35448 28172 35476
rect 28166 35436 28172 35448
rect 28224 35436 28230 35488
rect 29454 35436 29460 35488
rect 29512 35476 29518 35488
rect 32677 35479 32735 35485
rect 32677 35476 32689 35479
rect 29512 35448 32689 35476
rect 29512 35436 29518 35448
rect 32677 35445 32689 35448
rect 32723 35445 32735 35479
rect 32677 35439 32735 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1578 35272 1584 35284
rect 1539 35244 1584 35272
rect 1578 35232 1584 35244
rect 1636 35232 1642 35284
rect 1946 35232 1952 35284
rect 2004 35272 2010 35284
rect 2133 35275 2191 35281
rect 2133 35272 2145 35275
rect 2004 35244 2145 35272
rect 2004 35232 2010 35244
rect 2133 35241 2145 35244
rect 2179 35241 2191 35275
rect 6178 35272 6184 35284
rect 6139 35244 6184 35272
rect 2133 35235 2191 35241
rect 6178 35232 6184 35244
rect 6236 35232 6242 35284
rect 6730 35272 6736 35284
rect 6691 35244 6736 35272
rect 6730 35232 6736 35244
rect 6788 35232 6794 35284
rect 7466 35232 7472 35284
rect 7524 35272 7530 35284
rect 7837 35275 7895 35281
rect 7837 35272 7849 35275
rect 7524 35244 7849 35272
rect 7524 35232 7530 35244
rect 7837 35241 7849 35244
rect 7883 35241 7895 35275
rect 7837 35235 7895 35241
rect 9582 35232 9588 35284
rect 9640 35272 9646 35284
rect 9953 35275 10011 35281
rect 9953 35272 9965 35275
rect 9640 35244 9965 35272
rect 9640 35232 9646 35244
rect 9953 35241 9965 35244
rect 9999 35272 10011 35275
rect 10134 35272 10140 35284
rect 9999 35244 10140 35272
rect 9999 35241 10011 35244
rect 9953 35235 10011 35241
rect 10134 35232 10140 35244
rect 10192 35232 10198 35284
rect 10226 35232 10232 35284
rect 10284 35272 10290 35284
rect 10413 35275 10471 35281
rect 10413 35272 10425 35275
rect 10284 35244 10425 35272
rect 10284 35232 10290 35244
rect 10413 35241 10425 35244
rect 10459 35241 10471 35275
rect 12158 35272 12164 35284
rect 12119 35244 12164 35272
rect 10413 35235 10471 35241
rect 12158 35232 12164 35244
rect 12216 35232 12222 35284
rect 12710 35272 12716 35284
rect 12671 35244 12716 35272
rect 12710 35232 12716 35244
rect 12768 35232 12774 35284
rect 17494 35272 17500 35284
rect 17455 35244 17500 35272
rect 17494 35232 17500 35244
rect 17552 35232 17558 35284
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18049 35275 18107 35281
rect 18049 35272 18061 35275
rect 18012 35244 18061 35272
rect 18012 35232 18018 35244
rect 18049 35241 18061 35244
rect 18095 35241 18107 35275
rect 18598 35272 18604 35284
rect 18559 35244 18604 35272
rect 18049 35235 18107 35241
rect 18598 35232 18604 35244
rect 18656 35232 18662 35284
rect 19058 35232 19064 35284
rect 19116 35272 19122 35284
rect 19337 35275 19395 35281
rect 19337 35272 19349 35275
rect 19116 35244 19349 35272
rect 19116 35232 19122 35244
rect 19337 35241 19349 35244
rect 19383 35241 19395 35275
rect 20070 35272 20076 35284
rect 20031 35244 20076 35272
rect 19337 35235 19395 35241
rect 20070 35232 20076 35244
rect 20128 35232 20134 35284
rect 28810 35232 28816 35284
rect 28868 35272 28874 35284
rect 29549 35275 29607 35281
rect 29549 35272 29561 35275
rect 28868 35244 29561 35272
rect 28868 35232 28874 35244
rect 29549 35241 29561 35244
rect 29595 35241 29607 35275
rect 33502 35272 33508 35284
rect 33463 35244 33508 35272
rect 29549 35235 29607 35241
rect 33502 35232 33508 35244
rect 33560 35232 33566 35284
rect 35345 35275 35403 35281
rect 35345 35241 35357 35275
rect 35391 35272 35403 35275
rect 35802 35272 35808 35284
rect 35391 35244 35808 35272
rect 35391 35241 35403 35244
rect 35345 35235 35403 35241
rect 35802 35232 35808 35244
rect 35860 35232 35866 35284
rect 38013 35275 38071 35281
rect 38013 35241 38025 35275
rect 38059 35272 38071 35275
rect 38286 35272 38292 35284
rect 38059 35244 38292 35272
rect 38059 35241 38071 35244
rect 38013 35235 38071 35241
rect 38286 35232 38292 35244
rect 38344 35232 38350 35284
rect 1670 35164 1676 35216
rect 1728 35204 1734 35216
rect 2685 35207 2743 35213
rect 2685 35204 2697 35207
rect 1728 35176 2697 35204
rect 1728 35164 1734 35176
rect 2685 35173 2697 35176
rect 2731 35173 2743 35207
rect 2685 35167 2743 35173
rect 15289 35207 15347 35213
rect 15289 35173 15301 35207
rect 15335 35204 15347 35207
rect 17218 35204 17224 35216
rect 15335 35176 17224 35204
rect 15335 35173 15347 35176
rect 15289 35167 15347 35173
rect 17218 35164 17224 35176
rect 17276 35164 17282 35216
rect 18782 35164 18788 35216
rect 18840 35204 18846 35216
rect 20530 35204 20536 35216
rect 18840 35176 20536 35204
rect 18840 35164 18846 35176
rect 20530 35164 20536 35176
rect 20588 35164 20594 35216
rect 26329 35207 26387 35213
rect 26329 35173 26341 35207
rect 26375 35204 26387 35207
rect 28166 35204 28172 35216
rect 26375 35176 28172 35204
rect 26375 35173 26387 35176
rect 26329 35167 26387 35173
rect 28166 35164 28172 35176
rect 28224 35164 28230 35216
rect 28902 35164 28908 35216
rect 28960 35204 28966 35216
rect 34514 35204 34520 35216
rect 28960 35176 34520 35204
rect 28960 35164 28966 35176
rect 34514 35164 34520 35176
rect 34572 35204 34578 35216
rect 34701 35207 34759 35213
rect 34701 35204 34713 35207
rect 34572 35176 34713 35204
rect 34572 35164 34578 35176
rect 34701 35173 34713 35176
rect 34747 35173 34759 35207
rect 34701 35167 34759 35173
rect 12526 35096 12532 35148
rect 12584 35136 12590 35148
rect 13357 35139 13415 35145
rect 13357 35136 13369 35139
rect 12584 35108 13369 35136
rect 12584 35096 12590 35108
rect 13357 35105 13369 35108
rect 13403 35136 13415 35139
rect 18414 35136 18420 35148
rect 13403 35108 18420 35136
rect 13403 35105 13415 35108
rect 13357 35099 13415 35105
rect 18414 35096 18420 35108
rect 18472 35096 18478 35148
rect 18598 35096 18604 35148
rect 18656 35136 18662 35148
rect 29454 35136 29460 35148
rect 18656 35108 29460 35136
rect 18656 35096 18662 35108
rect 29454 35096 29460 35108
rect 29512 35096 29518 35148
rect 30101 35139 30159 35145
rect 30101 35105 30113 35139
rect 30147 35105 30159 35139
rect 30101 35099 30159 35105
rect 2869 35071 2927 35077
rect 2869 35037 2881 35071
rect 2915 35068 2927 35071
rect 10597 35071 10655 35077
rect 2915 35040 3924 35068
rect 2915 35037 2927 35040
rect 2869 35031 2927 35037
rect 3896 34944 3924 35040
rect 10597 35037 10609 35071
rect 10643 35068 10655 35071
rect 10778 35068 10784 35080
rect 10643 35040 10784 35068
rect 10643 35037 10655 35040
rect 10597 35031 10655 35037
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 15102 35068 15108 35080
rect 15063 35040 15108 35068
rect 15102 35028 15108 35040
rect 15160 35028 15166 35080
rect 15746 35068 15752 35080
rect 15707 35040 15752 35068
rect 15746 35028 15752 35040
rect 15804 35068 15810 35080
rect 16393 35071 16451 35077
rect 16393 35068 16405 35071
rect 15804 35040 16405 35068
rect 15804 35028 15810 35040
rect 16393 35037 16405 35040
rect 16439 35037 16451 35071
rect 16393 35031 16451 35037
rect 17218 35028 17224 35080
rect 17276 35068 17282 35080
rect 21174 35068 21180 35080
rect 17276 35040 21180 35068
rect 17276 35028 17282 35040
rect 21174 35028 21180 35040
rect 21232 35028 21238 35080
rect 28442 35028 28448 35080
rect 28500 35068 28506 35080
rect 30116 35068 30144 35099
rect 28500 35040 30144 35068
rect 28500 35028 28506 35040
rect 30558 35028 30564 35080
rect 30616 35068 30622 35080
rect 31389 35071 31447 35077
rect 31389 35068 31401 35071
rect 30616 35040 31401 35068
rect 30616 35028 30622 35040
rect 31389 35037 31401 35040
rect 31435 35068 31447 35071
rect 31662 35068 31668 35080
rect 31435 35040 31668 35068
rect 31435 35037 31447 35040
rect 31389 35031 31447 35037
rect 31662 35028 31668 35040
rect 31720 35028 31726 35080
rect 35529 35071 35587 35077
rect 35529 35037 35541 35071
rect 35575 35037 35587 35071
rect 35529 35031 35587 35037
rect 10962 34960 10968 35012
rect 11020 35000 11026 35012
rect 11149 35003 11207 35009
rect 11149 35000 11161 35003
rect 11020 34972 11161 35000
rect 11020 34960 11026 34972
rect 11149 34969 11161 34972
rect 11195 35000 11207 35003
rect 13170 35000 13176 35012
rect 11195 34972 13176 35000
rect 11195 34969 11207 34972
rect 11149 34963 11207 34969
rect 13170 34960 13176 34972
rect 13228 34960 13234 35012
rect 25498 35000 25504 35012
rect 15948 34972 25504 35000
rect 3878 34932 3884 34944
rect 3839 34904 3884 34932
rect 3878 34892 3884 34904
rect 3936 34892 3942 34944
rect 4433 34935 4491 34941
rect 4433 34901 4445 34935
rect 4479 34932 4491 34935
rect 4706 34932 4712 34944
rect 4479 34904 4712 34932
rect 4479 34901 4491 34904
rect 4433 34895 4491 34901
rect 4706 34892 4712 34904
rect 4764 34892 4770 34944
rect 4798 34892 4804 34944
rect 4856 34932 4862 34944
rect 4893 34935 4951 34941
rect 4893 34932 4905 34935
rect 4856 34904 4905 34932
rect 4856 34892 4862 34904
rect 4893 34901 4905 34904
rect 4939 34901 4951 34935
rect 5534 34932 5540 34944
rect 5495 34904 5540 34932
rect 4893 34895 4951 34901
rect 5534 34892 5540 34904
rect 5592 34892 5598 34944
rect 7098 34892 7104 34944
rect 7156 34932 7162 34944
rect 7285 34935 7343 34941
rect 7285 34932 7297 34935
rect 7156 34904 7297 34932
rect 7156 34892 7162 34904
rect 7285 34901 7297 34904
rect 7331 34901 7343 34935
rect 9030 34932 9036 34944
rect 8991 34904 9036 34932
rect 7285 34895 7343 34901
rect 9030 34892 9036 34904
rect 9088 34892 9094 34944
rect 11422 34892 11428 34944
rect 11480 34932 11486 34944
rect 11609 34935 11667 34941
rect 11609 34932 11621 34935
rect 11480 34904 11621 34932
rect 11480 34892 11486 34904
rect 11609 34901 11621 34904
rect 11655 34901 11667 34935
rect 14458 34932 14464 34944
rect 14419 34904 14464 34932
rect 11609 34895 11667 34901
rect 14458 34892 14464 34904
rect 14516 34892 14522 34944
rect 15948 34941 15976 34972
rect 25498 34960 25504 34972
rect 25556 34960 25562 35012
rect 25961 35003 26019 35009
rect 25961 34969 25973 35003
rect 26007 35000 26019 35003
rect 26234 35000 26240 35012
rect 26007 34972 26240 35000
rect 26007 34969 26019 34972
rect 25961 34963 26019 34969
rect 26234 34960 26240 34972
rect 26292 34960 26298 35012
rect 30009 35003 30067 35009
rect 30009 34969 30021 35003
rect 30055 35000 30067 35003
rect 33134 35000 33140 35012
rect 30055 34972 33140 35000
rect 30055 34969 30067 34972
rect 30009 34963 30067 34969
rect 33134 34960 33140 34972
rect 33192 34960 33198 35012
rect 15933 34935 15991 34941
rect 15933 34901 15945 34935
rect 15979 34901 15991 34935
rect 15933 34895 15991 34901
rect 16758 34892 16764 34944
rect 16816 34932 16822 34944
rect 16945 34935 17003 34941
rect 16945 34932 16957 34935
rect 16816 34904 16957 34932
rect 16816 34892 16822 34904
rect 16945 34901 16957 34904
rect 16991 34901 17003 34935
rect 21082 34932 21088 34944
rect 21043 34904 21088 34932
rect 16945 34895 17003 34901
rect 21082 34892 21088 34904
rect 21140 34892 21146 34944
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22833 34935 22891 34941
rect 22833 34932 22845 34935
rect 22520 34904 22845 34932
rect 22520 34892 22526 34904
rect 22833 34901 22845 34904
rect 22879 34932 22891 34935
rect 23014 34932 23020 34944
rect 22879 34904 23020 34932
rect 22879 34901 22891 34904
rect 22833 34895 22891 34901
rect 23014 34892 23020 34904
rect 23072 34892 23078 34944
rect 26418 34932 26424 34944
rect 26379 34904 26424 34932
rect 26418 34892 26424 34904
rect 26476 34892 26482 34944
rect 28994 34932 29000 34944
rect 28955 34904 29000 34932
rect 28994 34892 29000 34904
rect 29052 34932 29058 34944
rect 29917 34935 29975 34941
rect 29917 34932 29929 34935
rect 29052 34904 29929 34932
rect 29052 34892 29058 34904
rect 29917 34901 29929 34904
rect 29963 34901 29975 34935
rect 29917 34895 29975 34901
rect 30374 34892 30380 34944
rect 30432 34932 30438 34944
rect 30837 34935 30895 34941
rect 30837 34932 30849 34935
rect 30432 34904 30849 34932
rect 30432 34892 30438 34904
rect 30837 34901 30849 34904
rect 30883 34932 30895 34935
rect 31018 34932 31024 34944
rect 30883 34904 31024 34932
rect 30883 34901 30895 34904
rect 30837 34895 30895 34901
rect 31018 34892 31024 34904
rect 31076 34892 31082 34944
rect 31938 34932 31944 34944
rect 31899 34904 31944 34932
rect 31938 34892 31944 34904
rect 31996 34892 32002 34944
rect 32950 34932 32956 34944
rect 32911 34904 32956 34932
rect 32950 34892 32956 34904
rect 33008 34892 33014 34944
rect 33594 34892 33600 34944
rect 33652 34932 33658 34944
rect 34057 34935 34115 34941
rect 34057 34932 34069 34935
rect 33652 34904 34069 34932
rect 33652 34892 33658 34904
rect 34057 34901 34069 34904
rect 34103 34932 34115 34935
rect 34238 34932 34244 34944
rect 34103 34904 34244 34932
rect 34103 34901 34115 34904
rect 34057 34895 34115 34901
rect 34238 34892 34244 34904
rect 34296 34892 34302 34944
rect 35544 34932 35572 35031
rect 35894 35028 35900 35080
rect 35952 35068 35958 35080
rect 35989 35071 36047 35077
rect 35989 35068 36001 35071
rect 35952 35040 36001 35068
rect 35952 35028 35958 35040
rect 35989 35037 36001 35040
rect 36035 35037 36047 35071
rect 35989 35031 36047 35037
rect 37274 35028 37280 35080
rect 37332 35068 37338 35080
rect 37829 35071 37887 35077
rect 37829 35068 37841 35071
rect 37332 35040 37841 35068
rect 37332 35028 37338 35040
rect 37829 35037 37841 35040
rect 37875 35068 37887 35071
rect 38746 35068 38752 35080
rect 37875 35040 38752 35068
rect 37875 35037 37887 35040
rect 37829 35031 37887 35037
rect 38746 35028 38752 35040
rect 38804 35028 38810 35080
rect 36256 35003 36314 35009
rect 36256 34969 36268 35003
rect 36302 35000 36314 35003
rect 36446 35000 36452 35012
rect 36302 34972 36452 35000
rect 36302 34969 36314 34972
rect 36256 34963 36314 34969
rect 36446 34960 36452 34972
rect 36504 34960 36510 35012
rect 37369 34935 37427 34941
rect 37369 34932 37381 34935
rect 35544 34904 37381 34932
rect 37369 34901 37381 34904
rect 37415 34901 37427 34935
rect 37369 34895 37427 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2590 34728 2596 34740
rect 2551 34700 2596 34728
rect 2590 34688 2596 34700
rect 2648 34688 2654 34740
rect 12066 34728 12072 34740
rect 12027 34700 12072 34728
rect 12066 34688 12072 34700
rect 12124 34688 12130 34740
rect 12894 34728 12900 34740
rect 12855 34700 12900 34728
rect 12894 34688 12900 34700
rect 12952 34688 12958 34740
rect 13538 34688 13544 34740
rect 13596 34728 13602 34740
rect 15102 34728 15108 34740
rect 13596 34700 15108 34728
rect 13596 34688 13602 34700
rect 15102 34688 15108 34700
rect 15160 34728 15166 34740
rect 15657 34731 15715 34737
rect 15657 34728 15669 34731
rect 15160 34700 15669 34728
rect 15160 34688 15166 34700
rect 15657 34697 15669 34700
rect 15703 34697 15715 34731
rect 16942 34728 16948 34740
rect 16903 34700 16948 34728
rect 15657 34691 15715 34697
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 23293 34731 23351 34737
rect 23293 34697 23305 34731
rect 23339 34697 23351 34731
rect 23293 34691 23351 34697
rect 24213 34731 24271 34737
rect 24213 34697 24225 34731
rect 24259 34728 24271 34731
rect 27522 34728 27528 34740
rect 24259 34700 27528 34728
rect 24259 34697 24271 34700
rect 24213 34691 24271 34697
rect 6365 34663 6423 34669
rect 6365 34660 6377 34663
rect 4448 34632 6377 34660
rect 2774 34552 2780 34604
rect 2832 34592 2838 34604
rect 3234 34592 3240 34604
rect 2832 34564 3240 34592
rect 2832 34552 2838 34564
rect 3234 34552 3240 34564
rect 3292 34592 3298 34604
rect 4448 34601 4476 34632
rect 6365 34629 6377 34632
rect 6411 34660 6423 34663
rect 9490 34660 9496 34672
rect 6411 34632 9496 34660
rect 6411 34629 6423 34632
rect 6365 34623 6423 34629
rect 9490 34620 9496 34632
rect 9548 34620 9554 34672
rect 23308 34660 23336 34691
rect 27522 34688 27528 34700
rect 27580 34688 27586 34740
rect 36541 34731 36599 34737
rect 36541 34697 36553 34731
rect 36587 34728 36599 34731
rect 36630 34728 36636 34740
rect 36587 34700 36636 34728
rect 36587 34697 36599 34700
rect 36541 34691 36599 34697
rect 36630 34688 36636 34700
rect 36688 34688 36694 34740
rect 37274 34728 37280 34740
rect 37108 34700 37280 34728
rect 27982 34660 27988 34672
rect 12406 34632 22094 34660
rect 23308 34632 27988 34660
rect 3605 34595 3663 34601
rect 3605 34592 3617 34595
rect 3292 34564 3617 34592
rect 3292 34552 3298 34564
rect 3605 34561 3617 34564
rect 3651 34561 3663 34595
rect 3605 34555 3663 34561
rect 4433 34595 4491 34601
rect 4433 34561 4445 34595
rect 4479 34561 4491 34595
rect 4433 34555 4491 34561
rect 4700 34595 4758 34601
rect 4700 34561 4712 34595
rect 4746 34592 4758 34595
rect 5258 34592 5264 34604
rect 4746 34564 5264 34592
rect 4746 34561 4758 34564
rect 4700 34555 4758 34561
rect 5258 34552 5264 34564
rect 5316 34552 5322 34604
rect 9214 34592 9220 34604
rect 9127 34564 9220 34592
rect 9214 34552 9220 34564
rect 9272 34592 9278 34604
rect 12406 34592 12434 34632
rect 13906 34592 13912 34604
rect 9272 34564 12434 34592
rect 13867 34564 13912 34592
rect 9272 34552 9278 34564
rect 13906 34552 13912 34564
rect 13964 34552 13970 34604
rect 14182 34552 14188 34604
rect 14240 34592 14246 34604
rect 14553 34595 14611 34601
rect 14553 34592 14565 34595
rect 14240 34564 14565 34592
rect 14240 34552 14246 34564
rect 14553 34561 14565 34564
rect 14599 34561 14611 34595
rect 14553 34555 14611 34561
rect 14918 34552 14924 34604
rect 14976 34592 14982 34604
rect 18322 34601 18328 34604
rect 15105 34595 15163 34601
rect 15105 34592 15117 34595
rect 14976 34564 15117 34592
rect 14976 34552 14982 34564
rect 15105 34561 15117 34564
rect 15151 34561 15163 34595
rect 15105 34555 15163 34561
rect 18316 34555 18328 34601
rect 18380 34592 18386 34604
rect 18380 34564 18416 34592
rect 18322 34552 18328 34555
rect 18380 34552 18386 34564
rect 2866 34484 2872 34536
rect 2924 34524 2930 34536
rect 3053 34527 3111 34533
rect 3053 34524 3065 34527
rect 2924 34496 3065 34524
rect 2924 34484 2930 34496
rect 3053 34493 3065 34496
rect 3099 34493 3111 34527
rect 3053 34487 3111 34493
rect 9674 34484 9680 34536
rect 9732 34524 9738 34536
rect 9769 34527 9827 34533
rect 9769 34524 9781 34527
rect 9732 34496 9781 34524
rect 9732 34484 9738 34496
rect 9769 34493 9781 34496
rect 9815 34524 9827 34527
rect 9858 34524 9864 34536
rect 9815 34496 9864 34524
rect 9815 34493 9827 34496
rect 9769 34487 9827 34493
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 10778 34524 10784 34536
rect 10739 34496 10784 34524
rect 10778 34484 10784 34496
rect 10836 34484 10842 34536
rect 11238 34484 11244 34536
rect 11296 34524 11302 34536
rect 11517 34527 11575 34533
rect 11517 34524 11529 34527
rect 11296 34496 11529 34524
rect 11296 34484 11302 34496
rect 11517 34493 11529 34496
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 13722 34484 13728 34536
rect 13780 34524 13786 34536
rect 17589 34527 17647 34533
rect 17589 34524 17601 34527
rect 13780 34496 17601 34524
rect 13780 34484 13786 34496
rect 17589 34493 17601 34496
rect 17635 34524 17647 34527
rect 18049 34527 18107 34533
rect 18049 34524 18061 34527
rect 17635 34496 18061 34524
rect 17635 34493 17647 34496
rect 17589 34487 17647 34493
rect 18049 34493 18061 34496
rect 18095 34493 18107 34527
rect 18049 34487 18107 34493
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20254 34524 20260 34536
rect 20027 34496 20260 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 20254 34484 20260 34496
rect 20312 34484 20318 34536
rect 20438 34524 20444 34536
rect 20399 34496 20444 34524
rect 20438 34484 20444 34496
rect 20496 34484 20502 34536
rect 22066 34524 22094 34632
rect 27982 34620 27988 34632
rect 28040 34620 28046 34672
rect 34793 34663 34851 34669
rect 34793 34629 34805 34663
rect 34839 34660 34851 34663
rect 37108 34660 37136 34700
rect 37274 34688 37280 34700
rect 37332 34688 37338 34740
rect 37369 34731 37427 34737
rect 37369 34697 37381 34731
rect 37415 34728 37427 34731
rect 38010 34728 38016 34740
rect 37415 34700 38016 34728
rect 37415 34697 37427 34700
rect 37369 34691 37427 34697
rect 38010 34688 38016 34700
rect 38068 34688 38074 34740
rect 34839 34632 37136 34660
rect 34839 34629 34851 34632
rect 34793 34623 34851 34629
rect 37182 34620 37188 34672
rect 37240 34660 37246 34672
rect 39758 34660 39764 34672
rect 37240 34632 39764 34660
rect 37240 34620 37246 34632
rect 39758 34620 39764 34632
rect 39816 34620 39822 34672
rect 22833 34595 22891 34601
rect 22833 34561 22845 34595
rect 22879 34592 22891 34595
rect 23290 34592 23296 34604
rect 22879 34564 23296 34592
rect 22879 34561 22891 34564
rect 22833 34555 22891 34561
rect 23290 34552 23296 34564
rect 23348 34592 23354 34604
rect 23753 34595 23811 34601
rect 23753 34592 23765 34595
rect 23348 34564 23765 34592
rect 23348 34552 23354 34564
rect 23753 34561 23765 34564
rect 23799 34592 23811 34595
rect 26234 34592 26240 34604
rect 23799 34564 26240 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 26234 34552 26240 34564
rect 26292 34592 26298 34604
rect 27522 34592 27528 34604
rect 26292 34564 27528 34592
rect 26292 34552 26298 34564
rect 27522 34552 27528 34564
rect 27580 34552 27586 34604
rect 36725 34595 36783 34601
rect 36725 34561 36737 34595
rect 36771 34592 36783 34595
rect 37550 34592 37556 34604
rect 36771 34564 37556 34592
rect 36771 34561 36783 34564
rect 36725 34555 36783 34561
rect 37550 34552 37556 34564
rect 37608 34552 37614 34604
rect 37829 34595 37887 34601
rect 37829 34561 37841 34595
rect 37875 34561 37887 34595
rect 37829 34555 37887 34561
rect 24946 34524 24952 34536
rect 22066 34496 24952 34524
rect 24946 34484 24952 34496
rect 25004 34484 25010 34536
rect 32858 34484 32864 34536
rect 32916 34524 32922 34536
rect 32953 34527 33011 34533
rect 32953 34524 32965 34527
rect 32916 34496 32965 34524
rect 32916 34484 32922 34496
rect 32953 34493 32965 34496
rect 32999 34524 33011 34527
rect 33042 34524 33048 34536
rect 32999 34496 33048 34524
rect 32999 34493 33011 34496
rect 32953 34487 33011 34493
rect 33042 34484 33048 34496
rect 33100 34484 33106 34536
rect 33686 34524 33692 34536
rect 33647 34496 33692 34524
rect 33686 34484 33692 34496
rect 33744 34484 33750 34536
rect 34422 34484 34428 34536
rect 34480 34524 34486 34536
rect 35253 34527 35311 34533
rect 35253 34524 35265 34527
rect 34480 34496 35265 34524
rect 34480 34484 34486 34496
rect 35253 34493 35265 34496
rect 35299 34524 35311 34527
rect 36262 34524 36268 34536
rect 35299 34496 36268 34524
rect 35299 34493 35311 34496
rect 35253 34487 35311 34493
rect 36262 34484 36268 34496
rect 36320 34484 36326 34536
rect 37090 34484 37096 34536
rect 37148 34524 37154 34536
rect 37844 34524 37872 34555
rect 39390 34524 39396 34536
rect 37148 34496 37872 34524
rect 38028 34496 39396 34524
rect 37148 34484 37154 34496
rect 23109 34459 23167 34465
rect 23109 34425 23121 34459
rect 23155 34425 23167 34459
rect 24026 34456 24032 34468
rect 23987 34428 24032 34456
rect 23109 34419 23167 34425
rect 5810 34388 5816 34400
rect 5771 34360 5816 34388
rect 5810 34348 5816 34360
rect 5868 34348 5874 34400
rect 19426 34388 19432 34400
rect 19387 34360 19432 34388
rect 19426 34348 19432 34360
rect 19484 34348 19490 34400
rect 19978 34348 19984 34400
rect 20036 34388 20042 34400
rect 22281 34391 22339 34397
rect 22281 34388 22293 34391
rect 20036 34360 22293 34388
rect 20036 34348 20042 34360
rect 22281 34357 22293 34360
rect 22327 34388 22339 34391
rect 23124 34388 23152 34419
rect 24026 34416 24032 34428
rect 24084 34416 24090 34468
rect 38028 34465 38056 34496
rect 39390 34484 39396 34496
rect 39448 34484 39454 34536
rect 38013 34459 38071 34465
rect 38013 34425 38025 34459
rect 38059 34425 38071 34459
rect 38013 34419 38071 34425
rect 22327 34360 23152 34388
rect 22327 34357 22339 34360
rect 22281 34351 22339 34357
rect 35802 34348 35808 34400
rect 35860 34388 35866 34400
rect 35989 34391 36047 34397
rect 35989 34388 36001 34391
rect 35860 34360 36001 34388
rect 35860 34348 35866 34360
rect 35989 34357 36001 34360
rect 36035 34357 36047 34391
rect 35989 34351 36047 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 18046 34184 18052 34196
rect 18007 34156 18052 34184
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 31294 34184 31300 34196
rect 31255 34156 31300 34184
rect 31294 34144 31300 34156
rect 31352 34144 31358 34196
rect 33134 34144 33140 34196
rect 33192 34184 33198 34196
rect 36357 34187 36415 34193
rect 36357 34184 36369 34187
rect 33192 34156 36369 34184
rect 33192 34144 33198 34156
rect 36357 34153 36369 34156
rect 36403 34153 36415 34187
rect 37182 34184 37188 34196
rect 37143 34156 37188 34184
rect 36357 34147 36415 34153
rect 37182 34144 37188 34156
rect 37240 34144 37246 34196
rect 37642 34144 37648 34196
rect 37700 34184 37706 34196
rect 37921 34187 37979 34193
rect 37921 34184 37933 34187
rect 37700 34156 37933 34184
rect 37700 34144 37706 34156
rect 37921 34153 37933 34156
rect 37967 34153 37979 34187
rect 37921 34147 37979 34153
rect 31478 34076 31484 34128
rect 31536 34116 31542 34128
rect 31662 34116 31668 34128
rect 31536 34088 31668 34116
rect 31536 34076 31542 34088
rect 31662 34076 31668 34088
rect 31720 34076 31726 34128
rect 35894 34076 35900 34128
rect 35952 34116 35958 34128
rect 35952 34088 35997 34116
rect 35952 34076 35958 34088
rect 28718 34008 28724 34060
rect 28776 34048 28782 34060
rect 35253 34051 35311 34057
rect 35253 34048 35265 34051
rect 28776 34020 35265 34048
rect 28776 34008 28782 34020
rect 35253 34017 35265 34020
rect 35299 34048 35311 34051
rect 35618 34048 35624 34060
rect 35299 34020 35624 34048
rect 35299 34017 35311 34020
rect 35253 34011 35311 34017
rect 35618 34008 35624 34020
rect 35676 34008 35682 34060
rect 9401 33983 9459 33989
rect 9401 33949 9413 33983
rect 9447 33980 9459 33983
rect 9490 33980 9496 33992
rect 9447 33952 9496 33980
rect 9447 33949 9459 33952
rect 9401 33943 9459 33949
rect 9490 33940 9496 33952
rect 9548 33980 9554 33992
rect 31478 33980 31484 33992
rect 9548 33952 11376 33980
rect 31439 33952 31484 33980
rect 9548 33940 9554 33952
rect 9668 33915 9726 33921
rect 9668 33881 9680 33915
rect 9714 33912 9726 33915
rect 10134 33912 10140 33924
rect 9714 33884 10140 33912
rect 9714 33881 9726 33884
rect 9668 33875 9726 33881
rect 10134 33872 10140 33884
rect 10192 33872 10198 33924
rect 10781 33847 10839 33853
rect 10781 33813 10793 33847
rect 10827 33844 10839 33847
rect 11054 33844 11060 33856
rect 10827 33816 11060 33844
rect 10827 33813 10839 33816
rect 10781 33807 10839 33813
rect 11054 33804 11060 33816
rect 11112 33804 11118 33856
rect 11348 33853 11376 33952
rect 31478 33940 31484 33952
rect 31536 33940 31542 33992
rect 33502 33940 33508 33992
rect 33560 33980 33566 33992
rect 34698 33980 34704 33992
rect 33560 33952 34704 33980
rect 33560 33940 33566 33952
rect 34698 33940 34704 33952
rect 34756 33940 34762 33992
rect 35710 33940 35716 33992
rect 35768 33980 35774 33992
rect 36541 33983 36599 33989
rect 36541 33980 36553 33983
rect 35768 33952 36553 33980
rect 35768 33940 35774 33952
rect 36541 33949 36553 33952
rect 36587 33949 36599 33983
rect 36541 33943 36599 33949
rect 36630 33940 36636 33992
rect 36688 33980 36694 33992
rect 37001 33983 37059 33989
rect 37001 33980 37013 33983
rect 36688 33952 37013 33980
rect 36688 33940 36694 33952
rect 37001 33949 37013 33952
rect 37047 33949 37059 33983
rect 37001 33943 37059 33949
rect 37737 33983 37795 33989
rect 37737 33949 37749 33983
rect 37783 33980 37795 33983
rect 38010 33980 38016 33992
rect 37783 33952 38016 33980
rect 37783 33949 37795 33952
rect 37737 33943 37795 33949
rect 38010 33940 38016 33952
rect 38068 33940 38074 33992
rect 20530 33872 20536 33924
rect 20588 33912 20594 33924
rect 38470 33912 38476 33924
rect 20588 33884 38476 33912
rect 20588 33872 20594 33884
rect 38470 33872 38476 33884
rect 38528 33872 38534 33924
rect 11333 33847 11391 33853
rect 11333 33813 11345 33847
rect 11379 33844 11391 33847
rect 13722 33844 13728 33856
rect 11379 33816 13728 33844
rect 11379 33813 11391 33816
rect 11333 33807 11391 33813
rect 13722 33804 13728 33816
rect 13780 33804 13786 33856
rect 16025 33847 16083 33853
rect 16025 33813 16037 33847
rect 16071 33844 16083 33847
rect 16114 33844 16120 33856
rect 16071 33816 16120 33844
rect 16071 33813 16083 33816
rect 16025 33807 16083 33813
rect 16114 33804 16120 33816
rect 16172 33804 16178 33856
rect 17126 33844 17132 33856
rect 17087 33816 17132 33844
rect 17126 33804 17132 33816
rect 17184 33804 17190 33856
rect 21266 33804 21272 33856
rect 21324 33844 21330 33856
rect 23569 33847 23627 33853
rect 23569 33844 23581 33847
rect 21324 33816 23581 33844
rect 21324 33804 21330 33816
rect 23569 33813 23581 33816
rect 23615 33844 23627 33847
rect 24026 33844 24032 33856
rect 23615 33816 24032 33844
rect 23615 33813 23627 33816
rect 23569 33807 23627 33813
rect 24026 33804 24032 33816
rect 24084 33804 24090 33856
rect 33870 33844 33876 33856
rect 33831 33816 33876 33844
rect 33870 33804 33876 33816
rect 33928 33804 33934 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 5258 33640 5264 33652
rect 5219 33612 5264 33640
rect 5258 33600 5264 33612
rect 5316 33600 5322 33652
rect 10134 33640 10140 33652
rect 10095 33612 10140 33640
rect 10134 33600 10140 33612
rect 10192 33600 10198 33652
rect 11054 33600 11060 33652
rect 11112 33640 11118 33652
rect 11609 33643 11667 33649
rect 11609 33640 11621 33643
rect 11112 33612 11621 33640
rect 11112 33600 11118 33612
rect 11609 33609 11621 33612
rect 11655 33640 11667 33643
rect 11698 33640 11704 33652
rect 11655 33612 11704 33640
rect 11655 33609 11667 33612
rect 11609 33603 11667 33609
rect 11698 33600 11704 33612
rect 11756 33600 11762 33652
rect 18322 33600 18328 33652
rect 18380 33640 18386 33652
rect 18417 33643 18475 33649
rect 18417 33640 18429 33643
rect 18380 33612 18429 33640
rect 18380 33600 18386 33612
rect 18417 33609 18429 33612
rect 18463 33609 18475 33643
rect 18417 33603 18475 33609
rect 29365 33643 29423 33649
rect 29365 33609 29377 33643
rect 29411 33640 29423 33643
rect 30006 33640 30012 33652
rect 29411 33612 30012 33640
rect 29411 33609 29423 33612
rect 29365 33603 29423 33609
rect 30006 33600 30012 33612
rect 30064 33600 30070 33652
rect 35710 33600 35716 33652
rect 35768 33640 35774 33652
rect 36633 33643 36691 33649
rect 36633 33640 36645 33643
rect 35768 33612 36645 33640
rect 35768 33600 35774 33612
rect 36633 33609 36645 33612
rect 36679 33609 36691 33643
rect 36633 33603 36691 33609
rect 37369 33643 37427 33649
rect 37369 33609 37381 33643
rect 37415 33640 37427 33643
rect 37918 33640 37924 33652
rect 37415 33612 37924 33640
rect 37415 33609 37427 33612
rect 37369 33603 37427 33609
rect 37918 33600 37924 33612
rect 37976 33600 37982 33652
rect 38013 33643 38071 33649
rect 38013 33609 38025 33643
rect 38059 33640 38071 33643
rect 38654 33640 38660 33652
rect 38059 33612 38660 33640
rect 38059 33609 38071 33612
rect 38013 33603 38071 33609
rect 38654 33600 38660 33612
rect 38712 33600 38718 33652
rect 5445 33507 5503 33513
rect 5445 33473 5457 33507
rect 5491 33504 5503 33507
rect 6914 33504 6920 33516
rect 5491 33476 6920 33504
rect 5491 33473 5503 33476
rect 5445 33467 5503 33473
rect 6914 33464 6920 33476
rect 6972 33464 6978 33516
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33473 10379 33507
rect 10321 33467 10379 33473
rect 10597 33507 10655 33513
rect 10597 33473 10609 33507
rect 10643 33504 10655 33507
rect 11054 33504 11060 33516
rect 10643 33476 11060 33504
rect 10643 33473 10655 33476
rect 10597 33467 10655 33473
rect 5721 33439 5779 33445
rect 5721 33405 5733 33439
rect 5767 33436 5779 33439
rect 5810 33436 5816 33448
rect 5767 33408 5816 33436
rect 5767 33405 5779 33408
rect 5721 33399 5779 33405
rect 5810 33396 5816 33408
rect 5868 33436 5874 33448
rect 6362 33436 6368 33448
rect 5868 33408 6368 33436
rect 5868 33396 5874 33408
rect 6362 33396 6368 33408
rect 6420 33396 6426 33448
rect 10336 33368 10364 33467
rect 11054 33464 11060 33476
rect 11112 33464 11118 33516
rect 11517 33507 11575 33513
rect 11517 33473 11529 33507
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 11793 33507 11851 33513
rect 11793 33473 11805 33507
rect 11839 33504 11851 33507
rect 18598 33504 18604 33516
rect 11839 33476 12388 33504
rect 18559 33476 18604 33504
rect 11839 33473 11851 33476
rect 11793 33467 11851 33473
rect 10502 33436 10508 33448
rect 10415 33408 10508 33436
rect 10502 33396 10508 33408
rect 10560 33436 10566 33448
rect 11532 33436 11560 33467
rect 10560 33408 11560 33436
rect 10560 33396 10566 33408
rect 12360 33377 12388 33476
rect 18598 33464 18604 33476
rect 18656 33464 18662 33516
rect 27522 33504 27528 33516
rect 27483 33476 27528 33504
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 29178 33504 29184 33516
rect 29139 33476 29184 33504
rect 29178 33464 29184 33476
rect 29236 33464 29242 33516
rect 37829 33507 37887 33513
rect 37829 33473 37841 33507
rect 37875 33504 37887 33507
rect 37875 33476 38792 33504
rect 37875 33473 37887 33476
rect 37829 33467 37887 33473
rect 38764 33448 38792 33476
rect 18877 33439 18935 33445
rect 18877 33405 18889 33439
rect 18923 33436 18935 33439
rect 19426 33436 19432 33448
rect 18923 33408 19432 33436
rect 18923 33405 18935 33408
rect 18877 33399 18935 33405
rect 19426 33396 19432 33408
rect 19484 33396 19490 33448
rect 27798 33436 27804 33448
rect 27759 33408 27804 33436
rect 27798 33396 27804 33408
rect 27856 33396 27862 33448
rect 38746 33396 38752 33448
rect 38804 33396 38810 33448
rect 11793 33371 11851 33377
rect 11793 33368 11805 33371
rect 10336 33340 11805 33368
rect 11793 33337 11805 33340
rect 11839 33337 11851 33371
rect 11793 33331 11851 33337
rect 12345 33371 12403 33377
rect 12345 33337 12357 33371
rect 12391 33368 12403 33371
rect 19518 33368 19524 33380
rect 12391 33340 19524 33368
rect 12391 33337 12403 33340
rect 12345 33331 12403 33337
rect 19518 33328 19524 33340
rect 19576 33328 19582 33380
rect 4890 33260 4896 33312
rect 4948 33300 4954 33312
rect 5629 33303 5687 33309
rect 5629 33300 5641 33303
rect 4948 33272 5641 33300
rect 4948 33260 4954 33272
rect 5629 33269 5641 33272
rect 5675 33269 5687 33303
rect 5629 33263 5687 33269
rect 8018 33260 8024 33312
rect 8076 33300 8082 33312
rect 10502 33300 10508 33312
rect 8076 33272 10508 33300
rect 8076 33260 8082 33272
rect 10502 33260 10508 33272
rect 10560 33260 10566 33312
rect 18785 33303 18843 33309
rect 18785 33269 18797 33303
rect 18831 33300 18843 33303
rect 19242 33300 19248 33312
rect 18831 33272 19248 33300
rect 18831 33269 18843 33272
rect 18785 33263 18843 33269
rect 19242 33260 19248 33272
rect 19300 33260 19306 33312
rect 27890 33260 27896 33312
rect 27948 33300 27954 33312
rect 35253 33303 35311 33309
rect 35253 33300 35265 33303
rect 27948 33272 35265 33300
rect 27948 33260 27954 33272
rect 35253 33269 35265 33272
rect 35299 33300 35311 33303
rect 35342 33300 35348 33312
rect 35299 33272 35348 33300
rect 35299 33269 35311 33272
rect 35253 33263 35311 33269
rect 35342 33260 35348 33272
rect 35400 33260 35406 33312
rect 36173 33303 36231 33309
rect 36173 33269 36185 33303
rect 36219 33300 36231 33303
rect 36354 33300 36360 33312
rect 36219 33272 36360 33300
rect 36219 33269 36231 33272
rect 36173 33263 36231 33269
rect 36354 33260 36360 33272
rect 36412 33260 36418 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 18598 33056 18604 33108
rect 18656 33096 18662 33108
rect 19521 33099 19579 33105
rect 19521 33096 19533 33099
rect 18656 33068 19533 33096
rect 18656 33056 18662 33068
rect 19521 33065 19533 33068
rect 19567 33065 19579 33099
rect 19521 33059 19579 33065
rect 28442 33028 28448 33040
rect 28403 33000 28448 33028
rect 28442 32988 28448 33000
rect 28500 32988 28506 33040
rect 36262 32920 36268 32972
rect 36320 32960 36326 32972
rect 36725 32963 36783 32969
rect 36725 32960 36737 32963
rect 36320 32932 36737 32960
rect 36320 32920 36326 32932
rect 36725 32929 36737 32932
rect 36771 32960 36783 32963
rect 37090 32960 37096 32972
rect 36771 32932 37096 32960
rect 36771 32929 36783 32932
rect 36725 32923 36783 32929
rect 37090 32920 37096 32932
rect 37148 32920 37154 32972
rect 19242 32892 19248 32904
rect 19203 32864 19248 32892
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 19518 32892 19524 32904
rect 19479 32864 19524 32892
rect 19518 32852 19524 32864
rect 19576 32892 19582 32904
rect 19981 32895 20039 32901
rect 19981 32892 19993 32895
rect 19576 32864 19993 32892
rect 19576 32852 19582 32864
rect 19981 32861 19993 32864
rect 20027 32892 20039 32895
rect 20530 32892 20536 32904
rect 20027 32864 20536 32892
rect 20027 32861 20039 32864
rect 19981 32855 20039 32861
rect 20530 32852 20536 32864
rect 20588 32852 20594 32904
rect 27798 32852 27804 32904
rect 27856 32892 27862 32904
rect 28261 32895 28319 32901
rect 28261 32892 28273 32895
rect 27856 32864 28273 32892
rect 27856 32852 27862 32864
rect 28261 32861 28273 32864
rect 28307 32892 28319 32895
rect 32766 32892 32772 32904
rect 28307 32864 32772 32892
rect 28307 32861 28319 32864
rect 28261 32855 28319 32861
rect 32766 32852 32772 32864
rect 32824 32892 32830 32904
rect 37829 32895 37887 32901
rect 37829 32892 37841 32895
rect 32824 32864 37841 32892
rect 32824 32852 32830 32864
rect 37829 32861 37841 32864
rect 37875 32861 37887 32895
rect 38102 32892 38108 32904
rect 38063 32864 38108 32892
rect 37829 32855 37887 32861
rect 38102 32852 38108 32864
rect 38160 32852 38166 32904
rect 9030 32716 9036 32768
rect 9088 32756 9094 32768
rect 18874 32756 18880 32768
rect 9088 32728 18880 32756
rect 9088 32716 9094 32728
rect 18874 32716 18880 32728
rect 18932 32716 18938 32768
rect 19337 32759 19395 32765
rect 19337 32725 19349 32759
rect 19383 32756 19395 32759
rect 19426 32756 19432 32768
rect 19383 32728 19432 32756
rect 19383 32725 19395 32728
rect 19337 32719 19395 32725
rect 19426 32716 19432 32728
rect 19484 32716 19490 32768
rect 36265 32759 36323 32765
rect 36265 32725 36277 32759
rect 36311 32756 36323 32759
rect 36538 32756 36544 32768
rect 36311 32728 36544 32756
rect 36311 32725 36323 32728
rect 36265 32719 36323 32725
rect 36538 32716 36544 32728
rect 36596 32716 36602 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 9766 32512 9772 32564
rect 9824 32552 9830 32564
rect 23106 32552 23112 32564
rect 9824 32524 23112 32552
rect 9824 32512 9830 32524
rect 23106 32512 23112 32524
rect 23164 32512 23170 32564
rect 26145 32555 26203 32561
rect 26145 32521 26157 32555
rect 26191 32552 26203 32555
rect 26326 32552 26332 32564
rect 26191 32524 26332 32552
rect 26191 32521 26203 32524
rect 26145 32515 26203 32521
rect 26326 32512 26332 32524
rect 26384 32512 26390 32564
rect 31478 32512 31484 32564
rect 31536 32552 31542 32564
rect 32125 32555 32183 32561
rect 32125 32552 32137 32555
rect 31536 32524 32137 32552
rect 31536 32512 31542 32524
rect 32125 32521 32137 32524
rect 32171 32521 32183 32555
rect 32125 32515 32183 32521
rect 10410 32444 10416 32496
rect 10468 32484 10474 32496
rect 27798 32484 27804 32496
rect 10468 32456 27804 32484
rect 10468 32444 10474 32456
rect 27798 32444 27804 32456
rect 27856 32444 27862 32496
rect 38102 32484 38108 32496
rect 38063 32456 38108 32484
rect 38102 32444 38108 32456
rect 38160 32444 38166 32496
rect 6733 32419 6791 32425
rect 6733 32385 6745 32419
rect 6779 32385 6791 32419
rect 6733 32379 6791 32385
rect 6917 32419 6975 32425
rect 6917 32385 6929 32419
rect 6963 32416 6975 32419
rect 8018 32416 8024 32428
rect 6963 32388 8024 32416
rect 6963 32385 6975 32388
rect 6917 32379 6975 32385
rect 6748 32348 6776 32379
rect 8018 32376 8024 32388
rect 8076 32376 8082 32428
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32416 13691 32419
rect 13722 32416 13728 32428
rect 13679 32388 13728 32416
rect 13679 32385 13691 32388
rect 13633 32379 13691 32385
rect 13722 32376 13728 32388
rect 13780 32416 13786 32428
rect 14366 32425 14372 32428
rect 14093 32419 14151 32425
rect 14093 32416 14105 32419
rect 13780 32388 14105 32416
rect 13780 32376 13786 32388
rect 14093 32385 14105 32388
rect 14139 32385 14151 32419
rect 14093 32379 14151 32385
rect 14360 32379 14372 32425
rect 14424 32416 14430 32428
rect 14424 32388 14460 32416
rect 14366 32376 14372 32379
rect 14424 32376 14430 32388
rect 25314 32376 25320 32428
rect 25372 32416 25378 32428
rect 25777 32419 25835 32425
rect 25777 32416 25789 32419
rect 25372 32388 25789 32416
rect 25372 32376 25378 32388
rect 25777 32385 25789 32388
rect 25823 32385 25835 32419
rect 25777 32379 25835 32385
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32416 26019 32419
rect 26234 32416 26240 32428
rect 26007 32388 26240 32416
rect 26007 32385 26019 32388
rect 25961 32379 26019 32385
rect 26234 32376 26240 32388
rect 26292 32376 26298 32428
rect 32493 32419 32551 32425
rect 32493 32416 32505 32419
rect 31496 32388 32505 32416
rect 6748 32320 7512 32348
rect 6914 32240 6920 32292
rect 6972 32280 6978 32292
rect 6972 32252 7017 32280
rect 6972 32240 6978 32252
rect 7484 32224 7512 32320
rect 7466 32212 7472 32224
rect 7427 32184 7472 32212
rect 7466 32172 7472 32184
rect 7524 32172 7530 32224
rect 14826 32172 14832 32224
rect 14884 32212 14890 32224
rect 15473 32215 15531 32221
rect 15473 32212 15485 32215
rect 14884 32184 15485 32212
rect 14884 32172 14890 32184
rect 15473 32181 15485 32184
rect 15519 32181 15531 32215
rect 25314 32212 25320 32224
rect 25275 32184 25320 32212
rect 15473 32175 15531 32181
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 26326 32172 26332 32224
rect 26384 32212 26390 32224
rect 31496 32221 31524 32388
rect 32493 32385 32505 32388
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32585 32419 32643 32425
rect 32585 32385 32597 32419
rect 32631 32416 32643 32419
rect 35342 32416 35348 32428
rect 32631 32388 35348 32416
rect 32631 32385 32643 32388
rect 32585 32379 32643 32385
rect 35342 32376 35348 32388
rect 35400 32376 35406 32428
rect 32766 32348 32772 32360
rect 32727 32320 32772 32348
rect 32766 32308 32772 32320
rect 32824 32308 32830 32360
rect 31481 32215 31539 32221
rect 31481 32212 31493 32215
rect 26384 32184 31493 32212
rect 26384 32172 26390 32184
rect 31481 32181 31493 32184
rect 31527 32181 31539 32215
rect 31481 32175 31539 32181
rect 37553 32215 37611 32221
rect 37553 32181 37565 32215
rect 37599 32212 37611 32215
rect 38010 32212 38016 32224
rect 37599 32184 38016 32212
rect 37599 32181 37611 32184
rect 37553 32175 37611 32181
rect 38010 32172 38016 32184
rect 38068 32172 38074 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 18506 31968 18512 32020
rect 18564 32008 18570 32020
rect 26326 32008 26332 32020
rect 18564 31980 26332 32008
rect 18564 31968 18570 31980
rect 26326 31968 26332 31980
rect 26384 31968 26390 32020
rect 26510 32008 26516 32020
rect 26471 31980 26516 32008
rect 26510 31968 26516 31980
rect 26568 31968 26574 32020
rect 28353 32011 28411 32017
rect 28353 31977 28365 32011
rect 28399 32008 28411 32011
rect 29178 32008 29184 32020
rect 28399 31980 29184 32008
rect 28399 31977 28411 31980
rect 28353 31971 28411 31977
rect 29178 31968 29184 31980
rect 29236 31968 29242 32020
rect 30098 31968 30104 32020
rect 30156 32008 30162 32020
rect 32858 32008 32864 32020
rect 30156 31980 32864 32008
rect 30156 31968 30162 31980
rect 32858 31968 32864 31980
rect 32916 31968 32922 32020
rect 27522 31900 27528 31952
rect 27580 31940 27586 31952
rect 27580 31912 28212 31940
rect 27580 31900 27586 31912
rect 21450 31832 21456 31884
rect 21508 31872 21514 31884
rect 27433 31875 27491 31881
rect 27433 31872 27445 31875
rect 21508 31844 27445 31872
rect 21508 31832 21514 31844
rect 27433 31841 27445 31844
rect 27479 31872 27491 31875
rect 27479 31844 28028 31872
rect 27479 31841 27491 31844
rect 27433 31835 27491 31841
rect 13262 31764 13268 31816
rect 13320 31804 13326 31816
rect 13630 31804 13636 31816
rect 13320 31776 13636 31804
rect 13320 31764 13326 31776
rect 13630 31764 13636 31776
rect 13688 31764 13694 31816
rect 25593 31807 25651 31813
rect 25593 31804 25605 31807
rect 16546 31776 25605 31804
rect 15102 31696 15108 31748
rect 15160 31736 15166 31748
rect 16546 31736 16574 31776
rect 25593 31773 25605 31776
rect 25639 31804 25651 31807
rect 26145 31807 26203 31813
rect 26145 31804 26157 31807
rect 25639 31776 26157 31804
rect 25639 31773 25651 31776
rect 25593 31767 25651 31773
rect 26145 31773 26157 31776
rect 26191 31773 26203 31807
rect 26145 31767 26203 31773
rect 26234 31764 26240 31816
rect 26292 31804 26298 31816
rect 26329 31807 26387 31813
rect 26329 31804 26341 31807
rect 26292 31776 26341 31804
rect 26292 31764 26298 31776
rect 26329 31773 26341 31776
rect 26375 31804 26387 31807
rect 27522 31804 27528 31816
rect 26375 31776 27528 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 27522 31764 27528 31776
rect 27580 31764 27586 31816
rect 28000 31813 28028 31844
rect 28184 31813 28212 31912
rect 27985 31807 28043 31813
rect 27985 31773 27997 31807
rect 28031 31773 28043 31807
rect 27985 31767 28043 31773
rect 28169 31807 28227 31813
rect 28169 31773 28181 31807
rect 28215 31804 28227 31807
rect 28442 31804 28448 31816
rect 28215 31776 28448 31804
rect 28215 31773 28227 31776
rect 28169 31767 28227 31773
rect 28442 31764 28448 31776
rect 28500 31764 28506 31816
rect 15160 31708 16574 31736
rect 15160 31696 15166 31708
rect 36170 31628 36176 31680
rect 36228 31668 36234 31680
rect 36446 31668 36452 31680
rect 36228 31640 36452 31668
rect 36228 31628 36234 31640
rect 36446 31628 36452 31640
rect 36504 31628 36510 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 34885 31467 34943 31473
rect 34885 31433 34897 31467
rect 34931 31433 34943 31467
rect 34885 31427 34943 31433
rect 34900 31396 34928 31427
rect 35342 31424 35348 31476
rect 35400 31464 35406 31476
rect 37921 31467 37979 31473
rect 37921 31464 37933 31467
rect 35400 31436 37933 31464
rect 35400 31424 35406 31436
rect 37921 31433 37933 31436
rect 37967 31433 37979 31467
rect 37921 31427 37979 31433
rect 36170 31396 36176 31408
rect 34900 31368 36176 31396
rect 36170 31356 36176 31368
rect 36228 31356 36234 31408
rect 36372 31368 36768 31396
rect 33042 31288 33048 31340
rect 33100 31328 33106 31340
rect 34701 31331 34759 31337
rect 34701 31328 34713 31331
rect 33100 31300 34713 31328
rect 33100 31288 33106 31300
rect 34701 31297 34713 31300
rect 34747 31297 34759 31331
rect 34701 31291 34759 31297
rect 35894 31288 35900 31340
rect 35952 31328 35958 31340
rect 36372 31328 36400 31368
rect 35952 31300 36400 31328
rect 35952 31288 35958 31300
rect 36446 31288 36452 31340
rect 36504 31337 36510 31340
rect 36740 31337 36768 31368
rect 36504 31328 36516 31337
rect 36725 31331 36783 31337
rect 36504 31300 36549 31328
rect 36504 31291 36516 31300
rect 36725 31297 36737 31331
rect 36771 31297 36783 31331
rect 36725 31291 36783 31297
rect 37461 31331 37519 31337
rect 37461 31297 37473 31331
rect 37507 31328 37519 31331
rect 38102 31328 38108 31340
rect 37507 31300 38108 31328
rect 37507 31297 37519 31300
rect 37461 31291 37519 31297
rect 36504 31288 36510 31291
rect 38102 31288 38108 31300
rect 38160 31288 38166 31340
rect 17310 31084 17316 31136
rect 17368 31124 17374 31136
rect 22646 31124 22652 31136
rect 17368 31096 22652 31124
rect 17368 31084 17374 31096
rect 22646 31084 22652 31096
rect 22704 31084 22710 31136
rect 33410 31084 33416 31136
rect 33468 31124 33474 31136
rect 35345 31127 35403 31133
rect 35345 31124 35357 31127
rect 33468 31096 35357 31124
rect 33468 31084 33474 31096
rect 35345 31093 35357 31096
rect 35391 31093 35403 31127
rect 35345 31087 35403 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 27062 30920 27068 30932
rect 27023 30892 27068 30920
rect 27062 30880 27068 30892
rect 27120 30880 27126 30932
rect 33042 30920 33048 30932
rect 33003 30892 33048 30920
rect 33042 30880 33048 30892
rect 33100 30880 33106 30932
rect 35253 30923 35311 30929
rect 35253 30889 35265 30923
rect 35299 30920 35311 30923
rect 35894 30920 35900 30932
rect 35299 30892 35900 30920
rect 35299 30889 35311 30892
rect 35253 30883 35311 30889
rect 35894 30880 35900 30892
rect 35952 30880 35958 30932
rect 32858 30852 32864 30864
rect 32819 30824 32864 30852
rect 32858 30812 32864 30824
rect 32916 30812 32922 30864
rect 27522 30744 27528 30796
rect 27580 30784 27586 30796
rect 27617 30787 27675 30793
rect 27617 30784 27629 30787
rect 27580 30756 27629 30784
rect 27580 30744 27586 30756
rect 27617 30753 27629 30756
rect 27663 30753 27675 30787
rect 27617 30747 27675 30753
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 1903 30688 3801 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 2124 30651 2182 30657
rect 2124 30617 2136 30651
rect 2170 30648 2182 30651
rect 2170 30620 2452 30648
rect 2170 30617 2182 30620
rect 2124 30611 2182 30617
rect 2424 30580 2452 30620
rect 2682 30608 2688 30660
rect 2740 30648 2746 30660
rect 2792 30648 2820 30688
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 4801 30719 4859 30725
rect 4801 30685 4813 30719
rect 4847 30716 4859 30719
rect 4890 30716 4896 30728
rect 4847 30688 4896 30716
rect 4847 30685 4859 30688
rect 4801 30679 4859 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 4985 30719 5043 30725
rect 4985 30685 4997 30719
rect 5031 30716 5043 30719
rect 23661 30719 23719 30725
rect 5031 30688 5580 30716
rect 5031 30685 5043 30688
rect 4985 30679 5043 30685
rect 2740 30620 2820 30648
rect 2740 30608 2746 30620
rect 3142 30580 3148 30592
rect 2424 30552 3148 30580
rect 3142 30540 3148 30552
rect 3200 30540 3206 30592
rect 3237 30583 3295 30589
rect 3237 30549 3249 30583
rect 3283 30580 3295 30583
rect 4062 30580 4068 30592
rect 3283 30552 4068 30580
rect 3283 30549 3295 30552
rect 3237 30543 3295 30549
rect 4062 30540 4068 30552
rect 4120 30540 4126 30592
rect 4890 30580 4896 30592
rect 4851 30552 4896 30580
rect 4890 30540 4896 30552
rect 4948 30540 4954 30592
rect 5552 30589 5580 30688
rect 23661 30685 23673 30719
rect 23707 30716 23719 30719
rect 23707 30688 24532 30716
rect 23707 30685 23719 30688
rect 23661 30679 23719 30685
rect 18782 30608 18788 30660
rect 18840 30648 18846 30660
rect 18840 30620 22416 30648
rect 18840 30608 18846 30620
rect 5537 30583 5595 30589
rect 5537 30549 5549 30583
rect 5583 30580 5595 30583
rect 7466 30580 7472 30592
rect 5583 30552 7472 30580
rect 5583 30549 5595 30552
rect 5537 30543 5595 30549
rect 7466 30540 7472 30552
rect 7524 30540 7530 30592
rect 22278 30580 22284 30592
rect 22239 30552 22284 30580
rect 22278 30540 22284 30552
rect 22336 30540 22342 30592
rect 22388 30580 22416 30620
rect 22738 30608 22744 30660
rect 22796 30648 22802 30660
rect 24504 30657 24532 30688
rect 23394 30651 23452 30657
rect 23394 30648 23406 30651
rect 22796 30620 23406 30648
rect 22796 30608 22802 30620
rect 23394 30617 23406 30620
rect 23440 30617 23452 30651
rect 23394 30611 23452 30617
rect 24489 30651 24547 30657
rect 24489 30617 24501 30651
rect 24535 30648 24547 30651
rect 27154 30648 27160 30660
rect 24535 30620 27160 30648
rect 24535 30617 24547 30620
rect 24489 30611 24547 30617
rect 27154 30608 27160 30620
rect 27212 30608 27218 30660
rect 32582 30648 32588 30660
rect 32543 30620 32588 30648
rect 32582 30608 32588 30620
rect 32640 30608 32646 30660
rect 26605 30583 26663 30589
rect 26605 30580 26617 30583
rect 22388 30552 26617 30580
rect 26605 30549 26617 30552
rect 26651 30580 26663 30583
rect 27433 30583 27491 30589
rect 27433 30580 27445 30583
rect 26651 30552 27445 30580
rect 26651 30549 26663 30552
rect 26605 30543 26663 30549
rect 27433 30549 27445 30552
rect 27479 30549 27491 30583
rect 27433 30543 27491 30549
rect 27525 30583 27583 30589
rect 27525 30549 27537 30583
rect 27571 30580 27583 30583
rect 37918 30580 37924 30592
rect 27571 30552 37924 30580
rect 27571 30549 27583 30552
rect 27525 30543 27583 30549
rect 37918 30540 37924 30552
rect 37976 30540 37982 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 4982 30376 4988 30388
rect 4943 30348 4988 30376
rect 4982 30336 4988 30348
rect 5040 30336 5046 30388
rect 5276 30348 5488 30376
rect 3142 30268 3148 30320
rect 3200 30308 3206 30320
rect 3605 30311 3663 30317
rect 3605 30308 3617 30311
rect 3200 30280 3617 30308
rect 3200 30268 3206 30280
rect 3605 30277 3617 30280
rect 3651 30277 3663 30311
rect 3605 30271 3663 30277
rect 5153 30311 5211 30317
rect 5153 30277 5165 30311
rect 5199 30308 5211 30311
rect 5276 30308 5304 30348
rect 5199 30280 5304 30308
rect 5353 30311 5411 30317
rect 5199 30277 5211 30280
rect 5153 30271 5211 30277
rect 5353 30277 5365 30311
rect 5399 30277 5411 30311
rect 5460 30308 5488 30348
rect 6196 30348 6500 30376
rect 5626 30308 5632 30320
rect 5460 30280 5632 30308
rect 5353 30271 5411 30277
rect 1578 30200 1584 30252
rect 1636 30240 1642 30252
rect 1857 30243 1915 30249
rect 1857 30240 1869 30243
rect 1636 30212 1869 30240
rect 1636 30200 1642 30212
rect 1857 30209 1869 30212
rect 1903 30209 1915 30243
rect 1857 30203 1915 30209
rect 3789 30243 3847 30249
rect 3789 30209 3801 30243
rect 3835 30240 3847 30243
rect 4890 30240 4896 30252
rect 3835 30212 4896 30240
rect 3835 30209 3847 30212
rect 3789 30203 3847 30209
rect 4890 30200 4896 30212
rect 4948 30200 4954 30252
rect 5368 30240 5396 30271
rect 5626 30268 5632 30280
rect 5684 30308 5690 30320
rect 6196 30308 6224 30348
rect 6362 30308 6368 30320
rect 5684 30280 6224 30308
rect 6323 30280 6368 30308
rect 5684 30268 5690 30280
rect 6362 30268 6368 30280
rect 6420 30268 6426 30320
rect 6472 30308 6500 30348
rect 11882 30336 11888 30388
rect 11940 30376 11946 30388
rect 12897 30379 12955 30385
rect 12897 30376 12909 30379
rect 11940 30348 12909 30376
rect 11940 30336 11946 30348
rect 12897 30345 12909 30348
rect 12943 30345 12955 30379
rect 22738 30376 22744 30388
rect 12897 30339 12955 30345
rect 18156 30348 20208 30376
rect 22699 30348 22744 30376
rect 6733 30311 6791 30317
rect 6733 30308 6745 30311
rect 6472 30280 6745 30308
rect 6733 30277 6745 30280
rect 6779 30277 6791 30311
rect 8018 30308 8024 30320
rect 7979 30280 8024 30308
rect 6733 30271 6791 30277
rect 8018 30268 8024 30280
rect 8076 30268 8082 30320
rect 11517 30311 11575 30317
rect 11517 30277 11529 30311
rect 11563 30308 11575 30311
rect 11606 30308 11612 30320
rect 11563 30280 11612 30308
rect 11563 30277 11575 30280
rect 11517 30271 11575 30277
rect 11606 30268 11612 30280
rect 11664 30268 11670 30320
rect 12986 30308 12992 30320
rect 11747 30277 11805 30283
rect 12947 30280 12992 30308
rect 11747 30274 11759 30277
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 5368 30212 6561 30240
rect 4062 30172 4068 30184
rect 4023 30144 4068 30172
rect 4062 30132 4068 30144
rect 4120 30172 4126 30184
rect 5368 30172 5396 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 6641 30243 6699 30249
rect 6641 30209 6653 30243
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30240 6975 30243
rect 7837 30243 7895 30249
rect 7837 30240 7849 30243
rect 6963 30212 7849 30240
rect 6963 30209 6975 30212
rect 6917 30203 6975 30209
rect 7837 30209 7849 30212
rect 7883 30240 7895 30243
rect 11330 30240 11336 30252
rect 7883 30212 11336 30240
rect 7883 30209 7895 30212
rect 7837 30203 7895 30209
rect 4120 30144 5396 30172
rect 4120 30132 4126 30144
rect 2133 30107 2191 30113
rect 2133 30073 2145 30107
rect 2179 30104 2191 30107
rect 6178 30104 6184 30116
rect 2179 30076 6184 30104
rect 2179 30073 2191 30076
rect 2133 30067 2191 30073
rect 6178 30064 6184 30076
rect 6236 30064 6242 30116
rect 3970 30036 3976 30048
rect 3931 30008 3976 30036
rect 3970 29996 3976 30008
rect 4028 29996 4034 30048
rect 4614 29996 4620 30048
rect 4672 30036 4678 30048
rect 5169 30039 5227 30045
rect 5169 30036 5181 30039
rect 4672 30008 5181 30036
rect 4672 29996 4678 30008
rect 5169 30005 5181 30008
rect 5215 30036 5227 30039
rect 6656 30036 6684 30203
rect 11330 30200 11336 30212
rect 11388 30200 11394 30252
rect 11732 30243 11759 30274
rect 11793 30252 11805 30277
rect 12986 30268 12992 30280
rect 13044 30268 13050 30320
rect 14366 30308 14372 30320
rect 14327 30280 14372 30308
rect 14366 30268 14372 30280
rect 14424 30268 14430 30320
rect 15473 30311 15531 30317
rect 15473 30308 15485 30311
rect 14568 30280 15485 30308
rect 11793 30243 11796 30252
rect 11732 30212 11796 30243
rect 11790 30200 11796 30212
rect 11848 30200 11854 30252
rect 14568 30249 14596 30280
rect 15473 30277 15485 30280
rect 15519 30277 15531 30311
rect 15473 30271 15531 30277
rect 15930 30268 15936 30320
rect 15988 30308 15994 30320
rect 18156 30308 18184 30348
rect 19137 30311 19195 30317
rect 19137 30308 19149 30311
rect 15988 30280 18184 30308
rect 18248 30280 19149 30308
rect 15988 30268 15994 30280
rect 12805 30243 12863 30249
rect 12805 30240 12817 30243
rect 11900 30212 12817 30240
rect 11606 30064 11612 30116
rect 11664 30104 11670 30116
rect 11900 30104 11928 30212
rect 12805 30209 12817 30212
rect 12851 30209 12863 30243
rect 12805 30203 12863 30209
rect 14553 30243 14611 30249
rect 14553 30209 14565 30243
rect 14599 30209 14611 30243
rect 14553 30203 14611 30209
rect 15381 30243 15439 30249
rect 15381 30209 15393 30243
rect 15427 30209 15439 30243
rect 15381 30203 15439 30209
rect 15565 30243 15623 30249
rect 15565 30209 15577 30243
rect 15611 30240 15623 30243
rect 17221 30243 17279 30249
rect 17221 30240 17233 30243
rect 15611 30212 17233 30240
rect 15611 30209 15623 30212
rect 15565 30203 15623 30209
rect 17221 30209 17233 30212
rect 17267 30240 17279 30243
rect 17267 30212 17448 30240
rect 17267 30209 17279 30212
rect 17221 30203 17279 30209
rect 14737 30175 14795 30181
rect 14737 30172 14749 30175
rect 11664 30076 11928 30104
rect 12406 30144 14749 30172
rect 11664 30064 11670 30076
rect 11698 30036 11704 30048
rect 5215 30008 6684 30036
rect 11659 30008 11704 30036
rect 5215 30005 5227 30008
rect 5169 29999 5227 30005
rect 11698 29996 11704 30008
rect 11756 29996 11762 30048
rect 11882 30036 11888 30048
rect 11843 30008 11888 30036
rect 11882 29996 11888 30008
rect 11940 30036 11946 30048
rect 12406 30036 12434 30144
rect 14737 30141 14749 30144
rect 14783 30141 14795 30175
rect 14737 30135 14795 30141
rect 14826 30132 14832 30184
rect 14884 30172 14890 30184
rect 15396 30172 15424 30203
rect 14884 30144 14977 30172
rect 15396 30144 16160 30172
rect 14884 30132 14890 30144
rect 12621 30107 12679 30113
rect 12621 30073 12633 30107
rect 12667 30104 12679 30107
rect 14844 30104 14872 30132
rect 12667 30076 14872 30104
rect 12667 30073 12679 30076
rect 12621 30067 12679 30073
rect 11940 30008 12434 30036
rect 13173 30039 13231 30045
rect 11940 29996 11946 30008
rect 13173 30005 13185 30039
rect 13219 30036 13231 30039
rect 15930 30036 15936 30048
rect 13219 30008 15936 30036
rect 13219 30005 13231 30008
rect 13173 29999 13231 30005
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 16132 30045 16160 30144
rect 17420 30104 17448 30212
rect 17512 30181 17540 30280
rect 18248 30249 18276 30280
rect 19137 30277 19149 30280
rect 19183 30308 19195 30311
rect 19242 30308 19248 30320
rect 19183 30280 19248 30308
rect 19183 30277 19195 30280
rect 19137 30271 19195 30277
rect 19242 30268 19248 30280
rect 19300 30268 19306 30320
rect 19337 30311 19395 30317
rect 19337 30277 19349 30311
rect 19383 30277 19395 30311
rect 19337 30271 19395 30277
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18325 30243 18383 30249
rect 18325 30209 18337 30243
rect 18371 30209 18383 30243
rect 18325 30203 18383 30209
rect 18509 30243 18567 30249
rect 18509 30209 18521 30243
rect 18555 30240 18567 30243
rect 18690 30240 18696 30252
rect 18555 30212 18696 30240
rect 18555 30209 18567 30212
rect 18509 30203 18567 30209
rect 17497 30175 17555 30181
rect 17497 30141 17509 30175
rect 17543 30141 17555 30175
rect 17497 30135 17555 30141
rect 18248 30104 18276 30203
rect 18340 30172 18368 30203
rect 18690 30200 18696 30212
rect 18748 30240 18754 30252
rect 19352 30240 19380 30271
rect 19426 30268 19432 30320
rect 19484 30308 19490 30320
rect 20180 30317 20208 30348
rect 22738 30336 22744 30348
rect 22796 30336 22802 30388
rect 32309 30379 32367 30385
rect 32309 30345 32321 30379
rect 32355 30345 32367 30379
rect 32309 30339 32367 30345
rect 20073 30311 20131 30317
rect 20073 30308 20085 30311
rect 19484 30280 20085 30308
rect 19484 30268 19490 30280
rect 20073 30277 20085 30280
rect 20119 30277 20131 30311
rect 20073 30271 20131 30277
rect 20165 30311 20223 30317
rect 20165 30277 20177 30311
rect 20211 30277 20223 30311
rect 20165 30271 20223 30277
rect 24946 30268 24952 30320
rect 25004 30308 25010 30320
rect 26970 30308 26976 30320
rect 25004 30280 26976 30308
rect 25004 30268 25010 30280
rect 26970 30268 26976 30280
rect 27028 30268 27034 30320
rect 32324 30308 32352 30339
rect 32582 30336 32588 30388
rect 32640 30376 32646 30388
rect 32769 30379 32827 30385
rect 32769 30376 32781 30379
rect 32640 30348 32781 30376
rect 32640 30336 32646 30348
rect 32769 30345 32781 30348
rect 32815 30345 32827 30379
rect 32769 30339 32827 30345
rect 32398 30308 32404 30320
rect 32324 30280 32404 30308
rect 32398 30268 32404 30280
rect 32456 30268 32462 30320
rect 32950 30268 32956 30320
rect 33008 30308 33014 30320
rect 33318 30308 33324 30320
rect 33008 30280 33324 30308
rect 33008 30268 33014 30280
rect 33318 30268 33324 30280
rect 33376 30268 33382 30320
rect 19981 30243 20039 30249
rect 19981 30240 19993 30243
rect 18748 30212 19993 30240
rect 18748 30200 18754 30212
rect 19981 30209 19993 30212
rect 20027 30209 20039 30243
rect 19981 30203 20039 30209
rect 22557 30243 22615 30249
rect 22557 30209 22569 30243
rect 22603 30240 22615 30243
rect 22922 30240 22928 30252
rect 22603 30212 22928 30240
rect 22603 30209 22615 30212
rect 22557 30203 22615 30209
rect 22922 30200 22928 30212
rect 22980 30200 22986 30252
rect 32214 30240 32220 30252
rect 32127 30212 32220 30240
rect 32214 30200 32220 30212
rect 32272 30240 32278 30252
rect 33410 30240 33416 30252
rect 32272 30212 33416 30240
rect 32272 30200 32278 30212
rect 33410 30200 33416 30212
rect 33468 30200 33474 30252
rect 19426 30172 19432 30184
rect 18340 30144 19432 30172
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 19797 30175 19855 30181
rect 19797 30141 19809 30175
rect 19843 30172 19855 30175
rect 22278 30172 22284 30184
rect 19843 30144 22284 30172
rect 19843 30141 19855 30144
rect 19797 30135 19855 30141
rect 22278 30132 22284 30144
rect 22336 30132 22342 30184
rect 32122 30172 32128 30184
rect 32083 30144 32128 30172
rect 32122 30132 32128 30144
rect 32180 30132 32186 30184
rect 32493 30175 32551 30181
rect 32493 30141 32505 30175
rect 32539 30141 32551 30175
rect 32493 30135 32551 30141
rect 32585 30175 32643 30181
rect 32585 30141 32597 30175
rect 32631 30141 32643 30175
rect 32585 30135 32643 30141
rect 17420 30076 18276 30104
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 18969 30107 19027 30113
rect 18969 30104 18981 30107
rect 18380 30076 18981 30104
rect 18380 30064 18386 30076
rect 18969 30073 18981 30076
rect 19015 30104 19027 30107
rect 22373 30107 22431 30113
rect 22373 30104 22385 30107
rect 19015 30076 22385 30104
rect 19015 30073 19027 30076
rect 18969 30067 19027 30073
rect 22373 30073 22385 30076
rect 22419 30073 22431 30107
rect 22373 30067 22431 30073
rect 30282 30064 30288 30116
rect 30340 30104 30346 30116
rect 32508 30104 32536 30135
rect 30340 30076 32536 30104
rect 30340 30064 30346 30076
rect 16117 30039 16175 30045
rect 16117 30005 16129 30039
rect 16163 30036 16175 30039
rect 16206 30036 16212 30048
rect 16163 30008 16212 30036
rect 16163 30005 16175 30008
rect 16117 29999 16175 30005
rect 16206 29996 16212 30008
rect 16264 29996 16270 30048
rect 18414 29996 18420 30048
rect 18472 30036 18478 30048
rect 18509 30039 18567 30045
rect 18509 30036 18521 30039
rect 18472 30008 18521 30036
rect 18472 29996 18478 30008
rect 18509 30005 18521 30008
rect 18555 30005 18567 30039
rect 18509 29999 18567 30005
rect 19153 30039 19211 30045
rect 19153 30005 19165 30039
rect 19199 30036 19211 30039
rect 19426 30036 19432 30048
rect 19199 30008 19432 30036
rect 19199 30005 19211 30008
rect 19153 29999 19211 30005
rect 19426 29996 19432 30008
rect 19484 29996 19490 30048
rect 20349 30039 20407 30045
rect 20349 30005 20361 30039
rect 20395 30036 20407 30039
rect 22278 30036 22284 30048
rect 20395 30008 22284 30036
rect 20395 30005 20407 30008
rect 20349 29999 20407 30005
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 30742 29996 30748 30048
rect 30800 30036 30806 30048
rect 31481 30039 31539 30045
rect 31481 30036 31493 30039
rect 30800 30008 31493 30036
rect 30800 29996 30806 30008
rect 31481 30005 31493 30008
rect 31527 30036 31539 30039
rect 32600 30036 32628 30135
rect 31527 30008 32628 30036
rect 31527 30005 31539 30008
rect 31481 29999 31539 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 6914 29792 6920 29844
rect 6972 29832 6978 29844
rect 7466 29832 7472 29844
rect 6972 29804 7472 29832
rect 6972 29792 6978 29804
rect 7466 29792 7472 29804
rect 7524 29832 7530 29844
rect 16206 29832 16212 29844
rect 7524 29804 16212 29832
rect 7524 29792 7530 29804
rect 16206 29792 16212 29804
rect 16264 29792 16270 29844
rect 32677 29835 32735 29841
rect 32677 29801 32689 29835
rect 32723 29832 32735 29835
rect 32858 29832 32864 29844
rect 32723 29804 32864 29832
rect 32723 29801 32735 29804
rect 32677 29795 32735 29801
rect 32858 29792 32864 29804
rect 32916 29792 32922 29844
rect 37918 29832 37924 29844
rect 37879 29804 37924 29832
rect 37918 29792 37924 29804
rect 37976 29792 37982 29844
rect 11333 29767 11391 29773
rect 11333 29733 11345 29767
rect 11379 29764 11391 29767
rect 11514 29764 11520 29776
rect 11379 29736 11520 29764
rect 11379 29733 11391 29736
rect 11333 29727 11391 29733
rect 11514 29724 11520 29736
rect 11572 29724 11578 29776
rect 32306 29724 32312 29776
rect 32364 29764 32370 29776
rect 33870 29764 33876 29776
rect 32364 29736 33876 29764
rect 32364 29724 32370 29736
rect 33870 29724 33876 29736
rect 33928 29724 33934 29776
rect 11790 29696 11796 29708
rect 11072 29668 11796 29696
rect 8018 29588 8024 29640
rect 8076 29628 8082 29640
rect 11072 29637 11100 29668
rect 11790 29656 11796 29668
rect 11848 29656 11854 29708
rect 15286 29656 15292 29708
rect 15344 29696 15350 29708
rect 25590 29696 25596 29708
rect 15344 29668 25596 29696
rect 15344 29656 15350 29668
rect 25590 29656 25596 29668
rect 25648 29656 25654 29708
rect 32122 29696 32128 29708
rect 26206 29668 32128 29696
rect 11057 29631 11115 29637
rect 11057 29628 11069 29631
rect 8076 29600 11069 29628
rect 8076 29588 8082 29600
rect 11057 29597 11069 29600
rect 11103 29597 11115 29631
rect 11057 29591 11115 29597
rect 11149 29631 11207 29637
rect 11149 29597 11161 29631
rect 11195 29628 11207 29631
rect 11698 29628 11704 29640
rect 11195 29600 11704 29628
rect 11195 29597 11207 29600
rect 11149 29591 11207 29597
rect 11698 29588 11704 29600
rect 11756 29588 11762 29640
rect 22278 29588 22284 29640
rect 22336 29628 22342 29640
rect 25409 29631 25467 29637
rect 25409 29628 25421 29631
rect 22336 29600 25421 29628
rect 22336 29588 22342 29600
rect 25409 29597 25421 29600
rect 25455 29628 25467 29631
rect 26206 29628 26234 29668
rect 32122 29656 32128 29668
rect 32180 29696 32186 29708
rect 32493 29699 32551 29705
rect 32493 29696 32505 29699
rect 32180 29668 32505 29696
rect 32180 29656 32186 29668
rect 32493 29665 32505 29668
rect 32539 29665 32551 29699
rect 32493 29659 32551 29665
rect 32214 29628 32220 29640
rect 25455 29600 26234 29628
rect 32175 29600 32220 29628
rect 25455 29597 25467 29600
rect 25409 29591 25467 29597
rect 32214 29588 32220 29600
rect 32272 29588 32278 29640
rect 32309 29631 32367 29637
rect 32309 29597 32321 29631
rect 32355 29597 32367 29631
rect 32309 29591 32367 29597
rect 8662 29520 8668 29572
rect 8720 29560 8726 29572
rect 9582 29560 9588 29572
rect 8720 29532 9588 29560
rect 8720 29520 8726 29532
rect 9582 29520 9588 29532
rect 9640 29560 9646 29572
rect 9861 29563 9919 29569
rect 9861 29560 9873 29563
rect 9640 29532 9873 29560
rect 9640 29520 9646 29532
rect 9861 29529 9873 29532
rect 9907 29529 9919 29563
rect 9861 29523 9919 29529
rect 10045 29563 10103 29569
rect 10045 29529 10057 29563
rect 10091 29560 10103 29563
rect 10134 29560 10140 29572
rect 10091 29532 10140 29560
rect 10091 29529 10103 29532
rect 10045 29523 10103 29529
rect 10134 29520 10140 29532
rect 10192 29520 10198 29572
rect 11330 29560 11336 29572
rect 11291 29532 11336 29560
rect 11330 29520 11336 29532
rect 11388 29560 11394 29572
rect 11606 29560 11612 29572
rect 11388 29532 11612 29560
rect 11388 29520 11394 29532
rect 11606 29520 11612 29532
rect 11664 29520 11670 29572
rect 25222 29560 25228 29572
rect 25183 29532 25228 29560
rect 25222 29520 25228 29532
rect 25280 29520 25286 29572
rect 31386 29520 31392 29572
rect 31444 29560 31450 29572
rect 32324 29560 32352 29591
rect 32398 29588 32404 29640
rect 32456 29628 32462 29640
rect 32582 29628 32588 29640
rect 32456 29600 32588 29628
rect 32456 29588 32462 29600
rect 32582 29588 32588 29600
rect 32640 29588 32646 29640
rect 37461 29631 37519 29637
rect 37461 29597 37473 29631
rect 37507 29628 37519 29631
rect 38102 29628 38108 29640
rect 37507 29600 38108 29628
rect 37507 29597 37519 29600
rect 37461 29591 37519 29597
rect 38102 29588 38108 29600
rect 38160 29588 38166 29640
rect 31444 29532 32352 29560
rect 31444 29520 31450 29532
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 9582 29248 9588 29300
rect 9640 29288 9646 29300
rect 10505 29291 10563 29297
rect 10505 29288 10517 29291
rect 9640 29260 10517 29288
rect 9640 29248 9646 29260
rect 10505 29257 10517 29260
rect 10551 29257 10563 29291
rect 10505 29251 10563 29257
rect 11517 29291 11575 29297
rect 11517 29257 11529 29291
rect 11563 29257 11575 29291
rect 22922 29288 22928 29300
rect 22883 29260 22928 29288
rect 11517 29251 11575 29257
rect 8932 29223 8990 29229
rect 8932 29189 8944 29223
rect 8978 29220 8990 29223
rect 11532 29220 11560 29251
rect 22922 29248 22928 29260
rect 22980 29248 22986 29300
rect 23477 29223 23535 29229
rect 23477 29220 23489 29223
rect 8978 29192 11560 29220
rect 22848 29192 23489 29220
rect 8978 29189 8990 29192
rect 8932 29183 8990 29189
rect 11514 29152 11520 29164
rect 11475 29124 11520 29152
rect 11514 29112 11520 29124
rect 11572 29112 11578 29164
rect 11609 29155 11667 29161
rect 11609 29121 11621 29155
rect 11655 29152 11667 29155
rect 11882 29152 11888 29164
rect 11655 29124 11888 29152
rect 11655 29121 11667 29124
rect 11609 29115 11667 29121
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 16206 29112 16212 29164
rect 16264 29152 16270 29164
rect 22848 29161 22876 29192
rect 23477 29189 23489 29192
rect 23523 29189 23535 29223
rect 23477 29183 23535 29189
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 16264 29124 22845 29152
rect 16264 29112 16270 29124
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 23017 29155 23075 29161
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 25222 29152 25228 29164
rect 23063 29124 25228 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 25222 29112 25228 29124
rect 25280 29112 25286 29164
rect 30282 29112 30288 29164
rect 30340 29152 30346 29164
rect 31113 29155 31171 29161
rect 31113 29152 31125 29155
rect 30340 29124 31125 29152
rect 30340 29112 30346 29124
rect 31113 29121 31125 29124
rect 31159 29121 31171 29155
rect 31113 29115 31171 29121
rect 8662 29084 8668 29096
rect 8623 29056 8668 29084
rect 8662 29044 8668 29056
rect 8720 29044 8726 29096
rect 11793 29087 11851 29093
rect 11793 29053 11805 29087
rect 11839 29084 11851 29087
rect 12253 29087 12311 29093
rect 12253 29084 12265 29087
rect 11839 29056 12265 29084
rect 11839 29053 11851 29056
rect 11793 29047 11851 29053
rect 12253 29053 12265 29056
rect 12299 29084 12311 29087
rect 13078 29084 13084 29096
rect 12299 29056 13084 29084
rect 12299 29053 12311 29056
rect 12253 29047 12311 29053
rect 13078 29044 13084 29056
rect 13136 29044 13142 29096
rect 10045 29019 10103 29025
rect 10045 28985 10057 29019
rect 10091 29016 10103 29019
rect 11330 29016 11336 29028
rect 10091 28988 11336 29016
rect 10091 28985 10103 28988
rect 10045 28979 10103 28985
rect 11330 28976 11336 28988
rect 11388 28976 11394 29028
rect 31297 29019 31355 29025
rect 31297 28985 31309 29019
rect 31343 29016 31355 29019
rect 31386 29016 31392 29028
rect 31343 28988 31392 29016
rect 31343 28985 31355 28988
rect 31297 28979 31355 28985
rect 31386 28976 31392 28988
rect 31444 28976 31450 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 6178 28744 6184 28756
rect 6139 28716 6184 28744
rect 6178 28704 6184 28716
rect 6236 28704 6242 28756
rect 6914 28744 6920 28756
rect 6875 28716 6920 28744
rect 6914 28704 6920 28716
rect 6972 28704 6978 28756
rect 18322 28676 18328 28688
rect 18283 28648 18328 28676
rect 18322 28636 18328 28648
rect 18380 28636 18386 28688
rect 15378 28568 15384 28620
rect 15436 28608 15442 28620
rect 28994 28608 29000 28620
rect 15436 28580 29000 28608
rect 15436 28568 15442 28580
rect 28994 28568 29000 28580
rect 29052 28568 29058 28620
rect 6178 28500 6184 28552
rect 6236 28540 6242 28552
rect 6730 28540 6736 28552
rect 6236 28512 6736 28540
rect 6236 28500 6242 28512
rect 6730 28500 6736 28512
rect 6788 28500 6794 28552
rect 9858 28500 9864 28552
rect 9916 28540 9922 28552
rect 9916 28512 18276 28540
rect 9916 28500 9922 28512
rect 18141 28475 18199 28481
rect 18141 28441 18153 28475
rect 18187 28441 18199 28475
rect 18248 28472 18276 28512
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 18472 28512 18517 28540
rect 18472 28500 18478 28512
rect 25774 28472 25780 28484
rect 18248 28444 25780 28472
rect 18141 28435 18199 28441
rect 17586 28404 17592 28416
rect 17547 28376 17592 28404
rect 17586 28364 17592 28376
rect 17644 28404 17650 28416
rect 18156 28404 18184 28435
rect 25774 28432 25780 28444
rect 25832 28432 25838 28484
rect 28994 28432 29000 28484
rect 29052 28472 29058 28484
rect 30653 28475 30711 28481
rect 30653 28472 30665 28475
rect 29052 28444 30665 28472
rect 29052 28432 29058 28444
rect 30653 28441 30665 28444
rect 30699 28441 30711 28475
rect 30653 28435 30711 28441
rect 30834 28432 30840 28484
rect 30892 28472 30898 28484
rect 35894 28472 35900 28484
rect 30892 28444 35900 28472
rect 30892 28432 30898 28444
rect 35894 28432 35900 28444
rect 35952 28432 35958 28484
rect 18414 28404 18420 28416
rect 17644 28376 18184 28404
rect 18375 28376 18420 28404
rect 17644 28364 17650 28376
rect 18414 28364 18420 28376
rect 18472 28364 18478 28416
rect 26418 28364 26424 28416
rect 26476 28404 26482 28416
rect 26513 28407 26571 28413
rect 26513 28404 26525 28407
rect 26476 28376 26525 28404
rect 26476 28364 26482 28376
rect 26513 28373 26525 28376
rect 26559 28373 26571 28407
rect 26513 28367 26571 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 29089 28203 29147 28209
rect 29089 28169 29101 28203
rect 29135 28200 29147 28203
rect 30834 28200 30840 28212
rect 29135 28172 30840 28200
rect 29135 28169 29147 28172
rect 29089 28163 29147 28169
rect 29104 28132 29132 28163
rect 30834 28160 30840 28172
rect 30892 28160 30898 28212
rect 27172 28104 29132 28132
rect 27172 28076 27200 28104
rect 31386 28092 31392 28144
rect 31444 28132 31450 28144
rect 32217 28135 32275 28141
rect 32217 28132 32229 28135
rect 31444 28104 32229 28132
rect 31444 28092 31450 28104
rect 32217 28101 32229 28104
rect 32263 28101 32275 28135
rect 32217 28095 32275 28101
rect 25222 28024 25228 28076
rect 25280 28064 25286 28076
rect 26142 28064 26148 28076
rect 25280 28036 26148 28064
rect 25280 28024 25286 28036
rect 26142 28024 26148 28036
rect 26200 28024 26206 28076
rect 26234 28024 26240 28076
rect 26292 28064 26298 28076
rect 26418 28064 26424 28076
rect 26292 28036 26337 28064
rect 26379 28036 26424 28064
rect 26292 28024 26298 28036
rect 26418 28024 26424 28036
rect 26476 28024 26482 28076
rect 27154 28064 27160 28076
rect 27067 28036 27160 28064
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27430 28073 27436 28076
rect 27424 28027 27436 28073
rect 27488 28064 27494 28076
rect 27488 28036 27524 28064
rect 27430 28024 27436 28027
rect 27488 28024 27494 28036
rect 31754 28024 31760 28076
rect 31812 28064 31818 28076
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31812 28036 32137 28064
rect 31812 28024 31818 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 32401 28067 32459 28073
rect 32401 28033 32413 28067
rect 32447 28064 32459 28067
rect 32582 28064 32588 28076
rect 32447 28036 32588 28064
rect 32447 28033 32459 28036
rect 32401 28027 32459 28033
rect 32582 28024 32588 28036
rect 32640 28024 32646 28076
rect 37461 28067 37519 28073
rect 37461 28033 37473 28067
rect 37507 28064 37519 28067
rect 38102 28064 38108 28076
rect 37507 28036 38108 28064
rect 37507 28033 37519 28036
rect 37461 28027 37519 28033
rect 38102 28024 38108 28036
rect 38160 28024 38166 28076
rect 28537 27931 28595 27937
rect 28537 27897 28549 27931
rect 28583 27928 28595 27931
rect 30282 27928 30288 27940
rect 28583 27900 30288 27928
rect 28583 27897 28595 27900
rect 28537 27891 28595 27897
rect 30282 27888 30288 27900
rect 30340 27888 30346 27940
rect 26421 27863 26479 27869
rect 26421 27829 26433 27863
rect 26467 27860 26479 27863
rect 27062 27860 27068 27872
rect 26467 27832 27068 27860
rect 26467 27829 26479 27832
rect 26421 27823 26479 27829
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 32398 27860 32404 27872
rect 32359 27832 32404 27860
rect 32398 27820 32404 27832
rect 32456 27820 32462 27872
rect 36078 27820 36084 27872
rect 36136 27860 36142 27872
rect 37921 27863 37979 27869
rect 37921 27860 37933 27863
rect 36136 27832 37933 27860
rect 36136 27820 36142 27832
rect 37921 27829 37933 27832
rect 37967 27829 37979 27863
rect 37921 27823 37979 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 27341 27659 27399 27665
rect 27341 27625 27353 27659
rect 27387 27656 27399 27659
rect 27430 27656 27436 27668
rect 27387 27628 27436 27656
rect 27387 27625 27399 27628
rect 27341 27619 27399 27625
rect 27430 27616 27436 27628
rect 27488 27616 27494 27668
rect 3970 27548 3976 27600
rect 4028 27588 4034 27600
rect 4801 27591 4859 27597
rect 4801 27588 4813 27591
rect 4028 27560 4813 27588
rect 4028 27548 4034 27560
rect 4801 27557 4813 27560
rect 4847 27557 4859 27591
rect 4801 27551 4859 27557
rect 5997 27591 6055 27597
rect 5997 27557 6009 27591
rect 6043 27588 6055 27591
rect 6914 27588 6920 27600
rect 6043 27560 6920 27588
rect 6043 27557 6055 27560
rect 5997 27551 6055 27557
rect 4522 27452 4528 27464
rect 4483 27424 4528 27452
rect 4522 27412 4528 27424
rect 4580 27412 4586 27464
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27421 4675 27455
rect 4816 27452 4844 27551
rect 5261 27455 5319 27461
rect 5261 27452 5273 27455
rect 4816 27424 5273 27452
rect 4617 27415 4675 27421
rect 5261 27421 5273 27424
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 5445 27455 5503 27461
rect 5445 27421 5457 27455
rect 5491 27452 5503 27455
rect 6012 27452 6040 27551
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 10778 27548 10784 27600
rect 10836 27588 10842 27600
rect 13538 27588 13544 27600
rect 10836 27560 13544 27588
rect 10836 27548 10842 27560
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 18690 27588 18696 27600
rect 18651 27560 18696 27588
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 26142 27548 26148 27600
rect 26200 27588 26206 27600
rect 37550 27588 37556 27600
rect 26200 27548 26234 27588
rect 37511 27560 37556 27588
rect 37550 27548 37556 27560
rect 37608 27548 37614 27600
rect 26206 27520 26234 27548
rect 26973 27523 27031 27529
rect 26973 27520 26985 27523
rect 26206 27492 26985 27520
rect 26973 27489 26985 27492
rect 27019 27520 27031 27523
rect 31754 27520 31760 27532
rect 27019 27492 31760 27520
rect 27019 27489 27031 27492
rect 26973 27483 27031 27489
rect 31754 27480 31760 27492
rect 31812 27480 31818 27532
rect 31941 27523 31999 27529
rect 31941 27489 31953 27523
rect 31987 27520 31999 27523
rect 35713 27523 35771 27529
rect 31987 27492 32628 27520
rect 31987 27489 31999 27492
rect 31941 27483 31999 27489
rect 17313 27455 17371 27461
rect 17313 27452 17325 27455
rect 5491 27424 6040 27452
rect 16776 27424 17325 27452
rect 5491 27421 5503 27424
rect 5445 27415 5503 27421
rect 4632 27384 4660 27415
rect 5626 27384 5632 27396
rect 4632 27356 5632 27384
rect 5626 27344 5632 27356
rect 5684 27344 5690 27396
rect 5350 27316 5356 27328
rect 5311 27288 5356 27316
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 8110 27276 8116 27328
rect 8168 27316 8174 27328
rect 14366 27316 14372 27328
rect 8168 27288 14372 27316
rect 8168 27276 8174 27288
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 15470 27276 15476 27328
rect 15528 27316 15534 27328
rect 16776 27325 16804 27424
rect 17313 27421 17325 27424
rect 17359 27421 17371 27455
rect 17313 27415 17371 27421
rect 17580 27455 17638 27461
rect 17580 27421 17592 27455
rect 17626 27452 17638 27455
rect 18414 27452 18420 27464
rect 17626 27424 18420 27452
rect 17626 27421 17638 27424
rect 17580 27415 17638 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 26234 27412 26240 27464
rect 26292 27452 26298 27464
rect 26881 27455 26939 27461
rect 26881 27452 26893 27455
rect 26292 27424 26893 27452
rect 26292 27412 26298 27424
rect 26881 27421 26893 27424
rect 26927 27421 26939 27455
rect 26881 27415 26939 27421
rect 26896 27384 26924 27415
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27157 27455 27215 27461
rect 27157 27452 27169 27455
rect 27120 27424 27169 27452
rect 27120 27412 27126 27424
rect 27157 27421 27169 27424
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 30834 27412 30840 27464
rect 30892 27452 30898 27464
rect 31481 27455 31539 27461
rect 31481 27452 31493 27455
rect 30892 27424 31493 27452
rect 30892 27412 30898 27424
rect 31481 27421 31493 27424
rect 31527 27421 31539 27455
rect 31481 27415 31539 27421
rect 31573 27455 31631 27461
rect 31573 27421 31585 27455
rect 31619 27421 31631 27455
rect 31573 27415 31631 27421
rect 31665 27455 31723 27461
rect 31665 27421 31677 27455
rect 31711 27421 31723 27455
rect 32398 27452 32404 27464
rect 32359 27424 32404 27452
rect 31665 27415 31723 27421
rect 31386 27384 31392 27396
rect 26896 27356 31392 27384
rect 31386 27344 31392 27356
rect 31444 27384 31450 27396
rect 31588 27384 31616 27415
rect 31444 27356 31616 27384
rect 31444 27344 31450 27356
rect 16761 27319 16819 27325
rect 16761 27316 16773 27319
rect 15528 27288 16773 27316
rect 15528 27276 15534 27288
rect 16761 27285 16773 27288
rect 16807 27285 16819 27319
rect 30834 27316 30840 27328
rect 30795 27288 30840 27316
rect 16761 27279 16819 27285
rect 30834 27276 30840 27288
rect 30892 27276 30898 27328
rect 31680 27316 31708 27415
rect 32398 27412 32404 27424
rect 32456 27412 32462 27464
rect 32600 27461 32628 27492
rect 35713 27489 35725 27523
rect 35759 27520 35771 27523
rect 35894 27520 35900 27532
rect 35759 27492 35900 27520
rect 35759 27489 35771 27492
rect 35713 27483 35771 27489
rect 35894 27480 35900 27492
rect 35952 27520 35958 27532
rect 36173 27523 36231 27529
rect 36173 27520 36185 27523
rect 35952 27492 36185 27520
rect 35952 27480 35958 27492
rect 36173 27489 36185 27492
rect 36219 27489 36231 27523
rect 36173 27483 36231 27489
rect 32585 27455 32643 27461
rect 32585 27421 32597 27455
rect 32631 27421 32643 27455
rect 32585 27415 32643 27421
rect 32493 27387 32551 27393
rect 32493 27353 32505 27387
rect 32539 27384 32551 27387
rect 35434 27384 35440 27396
rect 32539 27356 35440 27384
rect 32539 27353 32551 27356
rect 32493 27347 32551 27353
rect 35434 27344 35440 27356
rect 35492 27384 35498 27396
rect 36418 27387 36476 27393
rect 36418 27384 36430 27387
rect 35492 27356 36430 27384
rect 35492 27344 35498 27356
rect 36418 27353 36430 27356
rect 36464 27353 36476 27387
rect 36418 27347 36476 27353
rect 32582 27316 32588 27328
rect 31680 27288 32588 27316
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 19392 27084 31064 27112
rect 19392 27072 19398 27084
rect 14366 27004 14372 27056
rect 14424 27044 14430 27056
rect 26234 27044 26240 27056
rect 14424 27016 26240 27044
rect 14424 27004 14430 27016
rect 26234 27004 26240 27016
rect 26292 27004 26298 27056
rect 15013 26979 15071 26985
rect 15013 26945 15025 26979
rect 15059 26976 15071 26979
rect 15838 26976 15844 26988
rect 15059 26948 15844 26976
rect 15059 26945 15071 26948
rect 15013 26939 15071 26945
rect 15838 26936 15844 26948
rect 15896 26936 15902 26988
rect 16850 26936 16856 26988
rect 16908 26976 16914 26988
rect 19978 26976 19984 26988
rect 16908 26948 19984 26976
rect 16908 26936 16914 26948
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 31036 26976 31064 27084
rect 32582 27072 32588 27124
rect 32640 27112 32646 27124
rect 34333 27115 34391 27121
rect 34333 27112 34345 27115
rect 32640 27084 34345 27112
rect 32640 27072 32646 27084
rect 34333 27081 34345 27084
rect 34379 27081 34391 27115
rect 34333 27075 34391 27081
rect 33873 27047 33931 27053
rect 33873 27013 33885 27047
rect 33919 27044 33931 27047
rect 33919 27016 35756 27044
rect 33919 27013 33931 27016
rect 33873 27007 33931 27013
rect 31036 26948 34468 26976
rect 3878 26868 3884 26920
rect 3936 26908 3942 26920
rect 24670 26908 24676 26920
rect 3936 26880 24676 26908
rect 3936 26868 3942 26880
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 17218 26840 17224 26852
rect 15212 26812 17224 26840
rect 13078 26732 13084 26784
rect 13136 26772 13142 26784
rect 15212 26781 15240 26812
rect 17218 26800 17224 26812
rect 17276 26840 17282 26852
rect 17586 26840 17592 26852
rect 17276 26812 17592 26840
rect 17276 26800 17282 26812
rect 17586 26800 17592 26812
rect 17644 26800 17650 26852
rect 15197 26775 15255 26781
rect 15197 26772 15209 26775
rect 13136 26744 15209 26772
rect 13136 26732 13142 26744
rect 15197 26741 15209 26744
rect 15243 26741 15255 26775
rect 15838 26772 15844 26784
rect 15799 26744 15844 26772
rect 15197 26735 15255 26741
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 34440 26772 34468 26948
rect 35434 26936 35440 26988
rect 35492 26985 35498 26988
rect 35728 26985 35756 27016
rect 35492 26976 35504 26985
rect 35713 26979 35771 26985
rect 35492 26948 35537 26976
rect 35492 26939 35504 26948
rect 35713 26945 35725 26979
rect 35759 26976 35771 26979
rect 35894 26976 35900 26988
rect 35759 26948 35900 26976
rect 35759 26945 35771 26948
rect 35713 26939 35771 26945
rect 35492 26936 35498 26939
rect 35894 26936 35900 26948
rect 35952 26936 35958 26988
rect 37182 26772 37188 26784
rect 34440 26744 37188 26772
rect 37182 26732 37188 26744
rect 37240 26732 37246 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 15838 26528 15844 26580
rect 15896 26568 15902 26580
rect 30834 26568 30840 26580
rect 15896 26540 30840 26568
rect 15896 26528 15902 26540
rect 30834 26528 30840 26540
rect 30892 26528 30898 26580
rect 4157 26503 4215 26509
rect 4157 26469 4169 26503
rect 4203 26500 4215 26503
rect 5626 26500 5632 26512
rect 4203 26472 5632 26500
rect 4203 26469 4215 26472
rect 4157 26463 4215 26469
rect 5626 26460 5632 26472
rect 5684 26460 5690 26512
rect 5350 26432 5356 26444
rect 3988 26404 5356 26432
rect 3988 26373 4016 26404
rect 5350 26392 5356 26404
rect 5408 26392 5414 26444
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4249 26367 4307 26373
rect 4249 26333 4261 26367
rect 4295 26364 4307 26367
rect 4614 26364 4620 26376
rect 4295 26336 4620 26364
rect 4295 26333 4307 26336
rect 4249 26327 4307 26333
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 3786 26228 3792 26240
rect 3747 26200 3792 26228
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 3697 26027 3755 26033
rect 3697 25993 3709 26027
rect 3743 26024 3755 26027
rect 4614 26024 4620 26036
rect 3743 25996 4620 26024
rect 3743 25993 3755 25996
rect 3697 25987 3755 25993
rect 4614 25984 4620 25996
rect 4672 25984 4678 26036
rect 26418 25984 26424 26036
rect 26476 26024 26482 26036
rect 27065 26027 27123 26033
rect 27065 26024 27077 26027
rect 26476 25996 27077 26024
rect 26476 25984 26482 25996
rect 27065 25993 27077 25996
rect 27111 25993 27123 26027
rect 30834 26024 30840 26036
rect 30795 25996 30840 26024
rect 27065 25987 27123 25993
rect 30834 25984 30840 25996
rect 30892 25984 30898 26036
rect 2682 25956 2688 25968
rect 2332 25928 2688 25956
rect 2332 25897 2360 25928
rect 2682 25916 2688 25928
rect 2740 25956 2746 25968
rect 4157 25959 4215 25965
rect 4157 25956 4169 25959
rect 2740 25928 4169 25956
rect 2740 25916 2746 25928
rect 4157 25925 4169 25928
rect 4203 25956 4215 25959
rect 6914 25956 6920 25968
rect 4203 25928 6920 25956
rect 4203 25925 4215 25928
rect 4157 25919 4215 25925
rect 6914 25916 6920 25928
rect 6972 25956 6978 25968
rect 8389 25959 8447 25965
rect 8389 25956 8401 25959
rect 6972 25928 8401 25956
rect 6972 25916 6978 25928
rect 8389 25925 8401 25928
rect 8435 25956 8447 25959
rect 8662 25956 8668 25968
rect 8435 25928 8668 25956
rect 8435 25925 8447 25928
rect 8389 25919 8447 25925
rect 8662 25916 8668 25928
rect 8720 25916 8726 25968
rect 17034 25916 17040 25968
rect 17092 25956 17098 25968
rect 21450 25956 21456 25968
rect 17092 25928 21456 25956
rect 17092 25916 17098 25928
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 23753 25959 23811 25965
rect 23753 25956 23765 25959
rect 21836 25928 23765 25956
rect 2317 25891 2375 25897
rect 2317 25857 2329 25891
rect 2363 25857 2375 25891
rect 2317 25851 2375 25857
rect 2584 25891 2642 25897
rect 2584 25857 2596 25891
rect 2630 25888 2642 25891
rect 3786 25888 3792 25900
rect 2630 25860 3792 25888
rect 2630 25857 2642 25860
rect 2584 25851 2642 25857
rect 3786 25848 3792 25860
rect 3844 25848 3850 25900
rect 21836 25897 21864 25928
rect 23753 25925 23765 25928
rect 23799 25956 23811 25959
rect 27154 25956 27160 25968
rect 23799 25928 27160 25956
rect 23799 25925 23811 25928
rect 23753 25919 23811 25925
rect 27154 25916 27160 25928
rect 27212 25916 27218 25968
rect 30193 25959 30251 25965
rect 30193 25956 30205 25959
rect 27264 25928 30205 25956
rect 22094 25897 22100 25900
rect 21821 25891 21879 25897
rect 21821 25857 21833 25891
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 22088 25851 22100 25897
rect 22152 25888 22158 25900
rect 27264 25897 27292 25928
rect 30193 25925 30205 25928
rect 30239 25956 30251 25959
rect 30742 25956 30748 25968
rect 30239 25928 30748 25956
rect 30239 25925 30251 25928
rect 30193 25919 30251 25925
rect 30742 25916 30748 25928
rect 30800 25916 30806 25968
rect 26421 25891 26479 25897
rect 26421 25888 26433 25891
rect 22152 25860 22188 25888
rect 26206 25860 26433 25888
rect 22094 25848 22100 25851
rect 22152 25848 22158 25860
rect 8662 25712 8668 25764
rect 8720 25752 8726 25764
rect 13909 25755 13967 25761
rect 13909 25752 13921 25755
rect 8720 25724 13921 25752
rect 8720 25712 8726 25724
rect 13909 25721 13921 25724
rect 13955 25752 13967 25755
rect 15470 25752 15476 25764
rect 13955 25724 15476 25752
rect 13955 25721 13967 25724
rect 13909 25715 13967 25721
rect 15470 25712 15476 25724
rect 15528 25712 15534 25764
rect 26206 25752 26234 25860
rect 26421 25857 26433 25860
rect 26467 25888 26479 25891
rect 27249 25891 27307 25897
rect 27249 25888 27261 25891
rect 26467 25860 27261 25888
rect 26467 25857 26479 25860
rect 26421 25851 26479 25857
rect 27249 25857 27261 25860
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 38102 25752 38108 25764
rect 22756 25724 26234 25752
rect 38063 25724 38108 25752
rect 14366 25644 14372 25696
rect 14424 25684 14430 25696
rect 22756 25684 22784 25724
rect 38102 25712 38108 25724
rect 38160 25712 38166 25764
rect 14424 25656 22784 25684
rect 14424 25644 14430 25656
rect 23106 25644 23112 25696
rect 23164 25684 23170 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 23164 25656 23213 25684
rect 23164 25644 23170 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 6730 25440 6736 25492
rect 6788 25480 6794 25492
rect 9125 25483 9183 25489
rect 9125 25480 9137 25483
rect 6788 25452 9137 25480
rect 6788 25440 6794 25452
rect 9125 25449 9137 25452
rect 9171 25449 9183 25483
rect 13078 25480 13084 25492
rect 13039 25452 13084 25480
rect 9125 25443 9183 25449
rect 9140 25412 9168 25443
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 22005 25483 22063 25489
rect 22005 25449 22017 25483
rect 22051 25480 22063 25483
rect 22094 25480 22100 25492
rect 22051 25452 22100 25480
rect 22051 25449 22063 25452
rect 22005 25443 22063 25449
rect 22094 25440 22100 25452
rect 22152 25440 22158 25492
rect 22373 25483 22431 25489
rect 22373 25449 22385 25483
rect 22419 25480 22431 25483
rect 22419 25452 23244 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 9140 25384 12434 25412
rect 6914 25344 6920 25356
rect 6875 25316 6920 25344
rect 6914 25304 6920 25316
rect 6972 25304 6978 25356
rect 9140 25276 9168 25384
rect 12406 25344 12434 25384
rect 20530 25372 20536 25424
rect 20588 25412 20594 25424
rect 22830 25412 22836 25424
rect 20588 25384 22836 25412
rect 20588 25372 20594 25384
rect 22830 25372 22836 25384
rect 22888 25372 22894 25424
rect 22925 25415 22983 25421
rect 22925 25381 22937 25415
rect 22971 25381 22983 25415
rect 22925 25375 22983 25381
rect 14366 25344 14372 25356
rect 10060 25316 10364 25344
rect 12406 25316 14372 25344
rect 9861 25279 9919 25285
rect 9861 25276 9873 25279
rect 9140 25248 9873 25276
rect 9861 25245 9873 25248
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 7184 25211 7242 25217
rect 7184 25177 7196 25211
rect 7230 25208 7242 25211
rect 7926 25208 7932 25220
rect 7230 25180 7932 25208
rect 7230 25177 7242 25180
rect 7184 25171 7242 25177
rect 7926 25168 7932 25180
rect 7984 25168 7990 25220
rect 10060 25208 10088 25316
rect 10336 25285 10364 25316
rect 14366 25304 14372 25316
rect 14424 25304 14430 25356
rect 15470 25344 15476 25356
rect 15431 25316 15476 25344
rect 15470 25304 15476 25316
rect 15528 25304 15534 25356
rect 22940 25344 22968 25375
rect 22204 25316 22968 25344
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25276 10379 25279
rect 11606 25276 11612 25288
rect 10367 25248 11612 25276
rect 10367 25245 10379 25248
rect 10321 25239 10379 25245
rect 8312 25180 10088 25208
rect 10152 25208 10180 25239
rect 11606 25236 11612 25248
rect 11664 25236 11670 25288
rect 22204 25285 22232 25316
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 22465 25279 22523 25285
rect 22465 25245 22477 25279
rect 22511 25276 22523 25279
rect 23106 25276 23112 25288
rect 22511 25248 23112 25276
rect 22511 25245 22523 25248
rect 22465 25239 22523 25245
rect 11514 25208 11520 25220
rect 10152 25180 11520 25208
rect 8312 25149 8340 25180
rect 11514 25168 11520 25180
rect 11572 25168 11578 25220
rect 12986 25168 12992 25220
rect 13044 25208 13050 25220
rect 15206 25211 15264 25217
rect 15206 25208 15218 25211
rect 13044 25180 15218 25208
rect 13044 25168 13050 25180
rect 15206 25177 15218 25180
rect 15252 25177 15264 25211
rect 22480 25208 22508 25239
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23216 25285 23244 25452
rect 30926 25440 30932 25492
rect 30984 25480 30990 25492
rect 31021 25483 31079 25489
rect 31021 25480 31033 25483
rect 30984 25452 31033 25480
rect 30984 25440 30990 25452
rect 31021 25449 31033 25452
rect 31067 25449 31079 25483
rect 31021 25443 31079 25449
rect 31386 25304 31392 25356
rect 31444 25344 31450 25356
rect 31573 25347 31631 25353
rect 31573 25344 31585 25347
rect 31444 25316 31585 25344
rect 31444 25304 31450 25316
rect 31573 25313 31585 25316
rect 31619 25313 31631 25347
rect 31573 25307 31631 25313
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23382 25276 23388 25288
rect 23247 25248 23388 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25276 31539 25279
rect 36078 25276 36084 25288
rect 31527 25248 36084 25276
rect 31527 25245 31539 25248
rect 31481 25239 31539 25245
rect 36078 25236 36084 25248
rect 36136 25236 36142 25288
rect 15206 25171 15264 25177
rect 22204 25180 22508 25208
rect 22204 25152 22232 25180
rect 22830 25168 22836 25220
rect 22888 25208 22894 25220
rect 22925 25211 22983 25217
rect 22925 25208 22937 25211
rect 22888 25180 22937 25208
rect 22888 25168 22894 25180
rect 22925 25177 22937 25180
rect 22971 25208 22983 25211
rect 23661 25211 23719 25217
rect 23661 25208 23673 25211
rect 22971 25180 23673 25208
rect 22971 25177 22983 25180
rect 22925 25171 22983 25177
rect 23661 25177 23673 25180
rect 23707 25208 23719 25211
rect 25682 25208 25688 25220
rect 23707 25180 25688 25208
rect 23707 25177 23719 25180
rect 23661 25171 23719 25177
rect 25682 25168 25688 25180
rect 25740 25208 25746 25220
rect 26418 25208 26424 25220
rect 25740 25180 26424 25208
rect 25740 25168 25746 25180
rect 26418 25168 26424 25180
rect 26476 25168 26482 25220
rect 28813 25211 28871 25217
rect 28813 25177 28825 25211
rect 28859 25177 28871 25211
rect 28994 25208 29000 25220
rect 28955 25180 29000 25208
rect 28813 25171 28871 25177
rect 8297 25143 8355 25149
rect 8297 25109 8309 25143
rect 8343 25109 8355 25143
rect 9674 25140 9680 25152
rect 9635 25112 9680 25140
rect 8297 25103 8355 25109
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 14090 25140 14096 25152
rect 14051 25112 14096 25140
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 22186 25100 22192 25152
rect 22244 25100 22250 25152
rect 28166 25140 28172 25152
rect 28127 25112 28172 25140
rect 28166 25100 28172 25112
rect 28224 25140 28230 25152
rect 28828 25140 28856 25171
rect 28994 25168 29000 25180
rect 29052 25168 29058 25220
rect 28224 25112 28856 25140
rect 28224 25100 28230 25112
rect 31294 25100 31300 25152
rect 31352 25140 31358 25152
rect 31389 25143 31447 25149
rect 31389 25140 31401 25143
rect 31352 25112 31401 25140
rect 31352 25100 31358 25112
rect 31389 25109 31401 25112
rect 31435 25140 31447 25143
rect 32217 25143 32275 25149
rect 32217 25140 32229 25143
rect 31435 25112 32229 25140
rect 31435 25109 31447 25112
rect 31389 25103 31447 25109
rect 32217 25109 32229 25112
rect 32263 25109 32275 25143
rect 32217 25103 32275 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7926 24936 7932 24948
rect 7887 24908 7932 24936
rect 7926 24896 7932 24908
rect 7984 24896 7990 24948
rect 12986 24936 12992 24948
rect 12947 24908 12992 24936
rect 12986 24896 12992 24908
rect 13044 24896 13050 24948
rect 9674 24828 9680 24880
rect 9732 24828 9738 24880
rect 12618 24868 12624 24880
rect 11532 24840 12624 24868
rect 8113 24803 8171 24809
rect 8113 24769 8125 24803
rect 8159 24800 8171 24803
rect 9309 24803 9367 24809
rect 9309 24800 9321 24803
rect 8159 24772 9321 24800
rect 8159 24769 8171 24772
rect 8113 24763 8171 24769
rect 9309 24769 9321 24772
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24800 9551 24803
rect 9692 24800 9720 24828
rect 11532 24812 11560 24840
rect 12618 24828 12624 24840
rect 12676 24828 12682 24880
rect 12713 24871 12771 24877
rect 12713 24837 12725 24871
rect 12759 24837 12771 24871
rect 12713 24831 12771 24837
rect 10134 24800 10140 24812
rect 9539 24772 9720 24800
rect 10095 24772 10140 24800
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 11514 24800 11520 24812
rect 10367 24772 11008 24800
rect 11475 24772 11520 24800
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 10980 24741 11008 24772
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11664 24772 11713 24800
rect 11664 24760 11670 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 12526 24800 12532 24812
rect 12487 24772 12532 24800
rect 11701 24763 11759 24769
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24701 9735 24735
rect 9677 24695 9735 24701
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 12434 24732 12440 24744
rect 11011 24704 12440 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 9692 24664 9720 24695
rect 12434 24692 12440 24704
rect 12492 24692 12498 24744
rect 11609 24667 11667 24673
rect 11609 24664 11621 24667
rect 9692 24636 11621 24664
rect 11609 24633 11621 24636
rect 11655 24664 11667 24667
rect 11655 24636 12434 24664
rect 11655 24633 11667 24636
rect 11609 24627 11667 24633
rect 12406 24596 12434 24636
rect 12728 24596 12756 24831
rect 12897 24803 12955 24809
rect 12897 24769 12909 24803
rect 12943 24769 12955 24803
rect 12897 24763 12955 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24800 13047 24803
rect 13078 24800 13084 24812
rect 13035 24772 13084 24800
rect 13035 24769 13047 24772
rect 12989 24763 13047 24769
rect 12912 24732 12940 24763
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 14090 24800 14096 24812
rect 13679 24772 14096 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 12912 24704 13553 24732
rect 13541 24701 13553 24704
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 12406 24568 12756 24596
rect 20898 24556 20904 24608
rect 20956 24596 20962 24608
rect 28166 24596 28172 24608
rect 20956 24568 28172 24596
rect 20956 24556 20962 24568
rect 28166 24556 28172 24568
rect 28224 24556 28230 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 20898 24392 20904 24404
rect 12492 24364 20904 24392
rect 12492 24352 12498 24364
rect 20898 24352 20904 24364
rect 20956 24352 20962 24404
rect 25682 24392 25688 24404
rect 25643 24364 25688 24392
rect 25682 24352 25688 24364
rect 25740 24352 25746 24404
rect 12805 24259 12863 24265
rect 12805 24225 12817 24259
rect 12851 24256 12863 24259
rect 14090 24256 14096 24268
rect 12851 24228 14096 24256
rect 12851 24225 12863 24228
rect 12805 24219 12863 24225
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 11606 24148 11612 24200
rect 11664 24188 11670 24200
rect 12621 24191 12679 24197
rect 12621 24188 12633 24191
rect 11664 24160 12633 24188
rect 11664 24148 11670 24160
rect 12621 24157 12633 24160
rect 12667 24157 12679 24191
rect 12621 24151 12679 24157
rect 18874 24148 18880 24200
rect 18932 24188 18938 24200
rect 18932 24160 22094 24188
rect 18932 24148 18938 24160
rect 19426 24080 19432 24132
rect 19484 24120 19490 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 19484 24092 19625 24120
rect 19484 24080 19490 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 22066 24120 22094 24160
rect 23382 24148 23388 24200
rect 23440 24188 23446 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 23440 24160 25053 24188
rect 23440 24148 23446 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 25225 24191 25283 24197
rect 25225 24157 25237 24191
rect 25271 24188 25283 24191
rect 25700 24188 25728 24352
rect 26234 24284 26240 24336
rect 26292 24324 26298 24336
rect 29549 24327 29607 24333
rect 29549 24324 29561 24327
rect 26292 24296 29561 24324
rect 26292 24284 26298 24296
rect 29549 24293 29561 24296
rect 29595 24293 29607 24327
rect 29549 24287 29607 24293
rect 30377 24191 30435 24197
rect 30377 24188 30389 24191
rect 25271 24160 25728 24188
rect 25792 24160 30389 24188
rect 25271 24157 25283 24160
rect 25225 24151 25283 24157
rect 25792 24120 25820 24160
rect 30377 24157 30389 24160
rect 30423 24157 30435 24191
rect 30377 24151 30435 24157
rect 30561 24191 30619 24197
rect 30561 24157 30573 24191
rect 30607 24188 30619 24191
rect 31386 24188 31392 24200
rect 30607 24160 31392 24188
rect 30607 24157 30619 24160
rect 30561 24151 30619 24157
rect 22066 24092 25820 24120
rect 29733 24123 29791 24129
rect 19613 24083 19671 24089
rect 29733 24089 29745 24123
rect 29779 24089 29791 24123
rect 29914 24120 29920 24132
rect 29875 24092 29920 24120
rect 29733 24083 29791 24089
rect 12437 24055 12495 24061
rect 12437 24021 12449 24055
rect 12483 24052 12495 24055
rect 12526 24052 12532 24064
rect 12483 24024 12532 24052
rect 12483 24021 12495 24024
rect 12437 24015 12495 24021
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 25130 24052 25136 24064
rect 25091 24024 25136 24052
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 29748 24052 29776 24083
rect 29914 24080 29920 24092
rect 29972 24080 29978 24132
rect 30576 24052 30604 24151
rect 31386 24148 31392 24160
rect 31444 24148 31450 24200
rect 30745 24123 30803 24129
rect 30745 24089 30757 24123
rect 30791 24120 30803 24123
rect 30834 24120 30840 24132
rect 30791 24092 30840 24120
rect 30791 24089 30803 24092
rect 30745 24083 30803 24089
rect 30834 24080 30840 24092
rect 30892 24120 30898 24132
rect 31205 24123 31263 24129
rect 31205 24120 31217 24123
rect 30892 24092 31217 24120
rect 30892 24080 30898 24092
rect 31205 24089 31217 24092
rect 31251 24089 31263 24123
rect 31205 24083 31263 24089
rect 33778 24080 33784 24132
rect 33836 24120 33842 24132
rect 37829 24123 37887 24129
rect 37829 24120 37841 24123
rect 33836 24092 37841 24120
rect 33836 24080 33842 24092
rect 37829 24089 37841 24092
rect 37875 24089 37887 24123
rect 38010 24120 38016 24132
rect 37971 24092 38016 24120
rect 37829 24083 37887 24089
rect 38010 24080 38016 24092
rect 38068 24080 38074 24132
rect 29748 24024 30604 24052
rect 37369 24055 37427 24061
rect 37369 24021 37381 24055
rect 37415 24052 37427 24055
rect 38028 24052 38056 24080
rect 37415 24024 38056 24052
rect 37415 24021 37427 24024
rect 37369 24015 37427 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 37734 23848 37740 23860
rect 37695 23820 37740 23848
rect 37734 23808 37740 23820
rect 37792 23808 37798 23860
rect 13538 23740 13544 23792
rect 13596 23780 13602 23792
rect 31205 23783 31263 23789
rect 31205 23780 31217 23783
rect 13596 23752 31217 23780
rect 13596 23740 13602 23752
rect 31205 23749 31217 23752
rect 31251 23749 31263 23783
rect 31386 23780 31392 23792
rect 31347 23752 31392 23780
rect 31205 23743 31263 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 17586 23721 17592 23724
rect 17580 23675 17592 23721
rect 17644 23712 17650 23724
rect 31573 23715 31631 23721
rect 17644 23684 17680 23712
rect 17586 23672 17592 23675
rect 17644 23672 17650 23684
rect 31573 23681 31585 23715
rect 31619 23712 31631 23715
rect 31846 23712 31852 23724
rect 31619 23684 31852 23712
rect 31619 23681 31631 23684
rect 31573 23675 31631 23681
rect 31846 23672 31852 23684
rect 31904 23672 31910 23724
rect 37550 23672 37556 23724
rect 37608 23712 37614 23724
rect 37645 23715 37703 23721
rect 37645 23712 37657 23715
rect 37608 23684 37657 23712
rect 37608 23672 37614 23684
rect 37645 23681 37657 23684
rect 37691 23681 37703 23715
rect 37645 23675 37703 23681
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 16776 23616 17325 23644
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 16776 23517 16804 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 36630 23604 36636 23656
rect 36688 23644 36694 23656
rect 37829 23647 37887 23653
rect 37829 23644 37841 23647
rect 36688 23616 37841 23644
rect 36688 23604 36694 23616
rect 37829 23613 37841 23616
rect 37875 23613 37887 23647
rect 37829 23607 37887 23613
rect 18693 23579 18751 23585
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 20990 23576 20996 23588
rect 18739 23548 20996 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 20990 23536 20996 23548
rect 21048 23536 21054 23588
rect 37277 23579 37335 23585
rect 37277 23545 37289 23579
rect 37323 23576 37335 23579
rect 38838 23576 38844 23588
rect 37323 23548 38844 23576
rect 37323 23545 37335 23548
rect 37277 23539 37335 23545
rect 38838 23536 38844 23548
rect 38896 23536 38902 23588
rect 16761 23511 16819 23517
rect 16761 23508 16773 23511
rect 15988 23480 16773 23508
rect 15988 23468 15994 23480
rect 16761 23477 16773 23480
rect 16807 23477 16819 23511
rect 19426 23508 19432 23520
rect 19387 23480 19432 23508
rect 16761 23471 16819 23477
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 29914 23468 29920 23520
rect 29972 23508 29978 23520
rect 30009 23511 30067 23517
rect 30009 23508 30021 23511
rect 29972 23480 30021 23508
rect 29972 23468 29978 23480
rect 30009 23477 30021 23480
rect 30055 23477 30067 23511
rect 30009 23471 30067 23477
rect 31846 23468 31852 23520
rect 31904 23508 31910 23520
rect 32125 23511 32183 23517
rect 32125 23508 32137 23511
rect 31904 23480 32137 23508
rect 31904 23468 31910 23480
rect 32125 23477 32137 23480
rect 32171 23477 32183 23511
rect 32125 23471 32183 23477
rect 33962 23468 33968 23520
rect 34020 23508 34026 23520
rect 34514 23508 34520 23520
rect 34020 23480 34520 23508
rect 34020 23468 34026 23480
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 17218 23304 17224 23316
rect 17179 23276 17224 23304
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 17586 23264 17592 23316
rect 17644 23304 17650 23316
rect 18049 23307 18107 23313
rect 18049 23304 18061 23307
rect 17644 23276 18061 23304
rect 17644 23264 17650 23276
rect 18049 23273 18061 23276
rect 18095 23273 18107 23307
rect 18049 23267 18107 23273
rect 17236 23168 17264 23264
rect 20993 23239 21051 23245
rect 20993 23205 21005 23239
rect 21039 23205 21051 23239
rect 20993 23199 21051 23205
rect 17770 23168 17776 23180
rect 17236 23140 17776 23168
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 17954 23100 17960 23112
rect 17915 23072 17960 23100
rect 17954 23060 17960 23072
rect 18012 23060 18018 23112
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 21008 23100 21036 23199
rect 31386 23128 31392 23180
rect 31444 23168 31450 23180
rect 32493 23171 32551 23177
rect 32493 23168 32505 23171
rect 31444 23140 32505 23168
rect 31444 23128 31450 23140
rect 32493 23137 32505 23140
rect 32539 23137 32551 23171
rect 32493 23131 32551 23137
rect 18095 23072 21036 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 21174 23060 21180 23112
rect 21232 23100 21238 23112
rect 21269 23103 21327 23109
rect 21269 23100 21281 23103
rect 21232 23072 21281 23100
rect 21232 23060 21238 23072
rect 21269 23069 21281 23072
rect 21315 23069 21327 23103
rect 21269 23063 21327 23069
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23100 25835 23103
rect 27617 23103 27675 23109
rect 27617 23100 27629 23103
rect 25823 23072 27629 23100
rect 25823 23069 25835 23072
rect 25777 23063 25835 23069
rect 27617 23069 27629 23072
rect 27663 23100 27675 23103
rect 28258 23100 28264 23112
rect 27663 23072 28264 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 32217 23103 32275 23109
rect 32217 23069 32229 23103
rect 32263 23100 32275 23103
rect 33778 23100 33784 23112
rect 32263 23072 33784 23100
rect 32263 23069 32275 23072
rect 32217 23063 32275 23069
rect 33778 23060 33784 23072
rect 33836 23060 33842 23112
rect 37550 23060 37556 23112
rect 37608 23100 37614 23112
rect 38013 23103 38071 23109
rect 38013 23100 38025 23103
rect 37608 23072 38025 23100
rect 37608 23060 37614 23072
rect 38013 23069 38025 23072
rect 38059 23069 38071 23103
rect 38013 23063 38071 23069
rect 20990 23032 20996 23044
rect 20951 23004 20996 23032
rect 20990 22992 20996 23004
rect 21048 22992 21054 23044
rect 26050 23041 26056 23044
rect 26044 22995 26056 23041
rect 26108 23032 26114 23044
rect 26108 23004 26144 23032
rect 26050 22992 26056 22995
rect 26108 22992 26114 23004
rect 21177 22967 21235 22973
rect 21177 22933 21189 22967
rect 21223 22964 21235 22967
rect 22186 22964 22192 22976
rect 21223 22936 22192 22964
rect 21223 22933 21235 22936
rect 21177 22927 21235 22933
rect 22186 22924 22192 22936
rect 22244 22924 22250 22976
rect 27157 22967 27215 22973
rect 27157 22933 27169 22967
rect 27203 22964 27215 22967
rect 27246 22964 27252 22976
rect 27203 22936 27252 22964
rect 27203 22933 27215 22936
rect 27157 22927 27215 22933
rect 27246 22924 27252 22936
rect 27304 22924 27310 22976
rect 37553 22967 37611 22973
rect 37553 22933 37565 22967
rect 37599 22964 37611 22967
rect 37642 22964 37648 22976
rect 37599 22936 37648 22964
rect 37599 22933 37611 22936
rect 37553 22927 37611 22933
rect 37642 22924 37648 22936
rect 37700 22924 37706 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 10226 22720 10232 22772
rect 10284 22760 10290 22772
rect 20346 22760 20352 22772
rect 10284 22732 20352 22760
rect 10284 22720 10290 22732
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 25961 22763 26019 22769
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26050 22760 26056 22772
rect 26007 22732 26056 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 26050 22720 26056 22732
rect 26108 22720 26114 22772
rect 33226 22760 33232 22772
rect 33187 22732 33232 22760
rect 33226 22720 33232 22732
rect 33284 22720 33290 22772
rect 33689 22763 33747 22769
rect 33689 22729 33701 22763
rect 33735 22760 33747 22763
rect 37090 22760 37096 22772
rect 33735 22732 37096 22760
rect 33735 22729 33747 22732
rect 33689 22723 33747 22729
rect 37090 22720 37096 22732
rect 37148 22720 37154 22772
rect 37737 22763 37795 22769
rect 37737 22729 37749 22763
rect 37783 22760 37795 22763
rect 38470 22760 38476 22772
rect 37783 22732 38476 22760
rect 37783 22729 37795 22732
rect 37737 22723 37795 22729
rect 38470 22720 38476 22732
rect 38528 22720 38534 22772
rect 20990 22652 20996 22704
rect 21048 22692 21054 22704
rect 21048 22664 22140 22692
rect 21048 22652 21054 22664
rect 22112 22633 22140 22664
rect 22738 22652 22744 22704
rect 22796 22692 22802 22704
rect 35069 22695 35127 22701
rect 35069 22692 35081 22695
rect 22796 22664 35081 22692
rect 22796 22652 22802 22664
rect 35069 22661 35081 22664
rect 35115 22661 35127 22695
rect 35069 22655 35127 22661
rect 35621 22695 35679 22701
rect 35621 22661 35633 22695
rect 35667 22692 35679 22695
rect 35894 22692 35900 22704
rect 35667 22664 35900 22692
rect 35667 22661 35679 22664
rect 35621 22655 35679 22661
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 22020 22556 22048 22587
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 25188 22596 26157 22624
rect 25188 22584 25194 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 32950 22584 32956 22636
rect 33008 22624 33014 22636
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 33008 22596 33609 22624
rect 33008 22584 33014 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 22186 22556 22192 22568
rect 22020 22528 22192 22556
rect 22186 22516 22192 22528
rect 22244 22516 22250 22568
rect 26421 22559 26479 22565
rect 26421 22525 26433 22559
rect 26467 22556 26479 22559
rect 27246 22556 27252 22568
rect 26467 22528 27252 22556
rect 26467 22525 26479 22528
rect 26421 22519 26479 22525
rect 27246 22516 27252 22528
rect 27304 22516 27310 22568
rect 33778 22556 33784 22568
rect 33739 22528 33784 22556
rect 33778 22516 33784 22528
rect 33836 22516 33842 22568
rect 35084 22488 35112 22655
rect 35894 22652 35900 22664
rect 35952 22692 35958 22704
rect 36630 22692 36636 22704
rect 35952 22664 36636 22692
rect 35952 22652 35958 22664
rect 36630 22652 36636 22664
rect 36688 22652 36694 22704
rect 37642 22584 37648 22636
rect 37700 22624 37706 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37700 22596 37841 22624
rect 37700 22584 37706 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 35897 22491 35955 22497
rect 35897 22488 35909 22491
rect 35084 22460 35909 22488
rect 35897 22457 35909 22460
rect 35943 22457 35955 22491
rect 35897 22451 35955 22457
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21048 22392 21833 22420
rect 21048 22380 21054 22392
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 26329 22423 26387 22429
rect 26329 22389 26341 22423
rect 26375 22420 26387 22423
rect 26418 22420 26424 22432
rect 26375 22392 26424 22420
rect 26375 22389 26387 22392
rect 26329 22383 26387 22389
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 32769 22423 32827 22429
rect 32769 22389 32781 22423
rect 32815 22420 32827 22423
rect 32950 22420 32956 22432
rect 32815 22392 32956 22420
rect 32815 22389 32827 22392
rect 32769 22383 32827 22389
rect 32950 22380 32956 22392
rect 33008 22380 33014 22432
rect 36078 22420 36084 22432
rect 36039 22392 36084 22420
rect 36078 22380 36084 22392
rect 36136 22380 36142 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 31386 22148 31392 22160
rect 31220 22120 31392 22148
rect 17954 22040 17960 22092
rect 18012 22080 18018 22092
rect 20809 22083 20867 22089
rect 20809 22080 20821 22083
rect 18012 22052 20821 22080
rect 18012 22040 18018 22052
rect 20809 22049 20821 22052
rect 20855 22049 20867 22083
rect 21174 22080 21180 22092
rect 21135 22052 21180 22080
rect 20809 22043 20867 22049
rect 21174 22040 21180 22052
rect 21232 22080 21238 22092
rect 23382 22080 23388 22092
rect 21232 22052 23388 22080
rect 21232 22040 21238 22052
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 31220 22089 31248 22120
rect 31386 22108 31392 22120
rect 31444 22108 31450 22160
rect 31205 22083 31263 22089
rect 31205 22049 31217 22083
rect 31251 22049 31263 22083
rect 31205 22043 31263 22049
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 22012 4675 22015
rect 20990 22012 20996 22024
rect 4663 21984 6592 22012
rect 20951 21984 20996 22012
rect 4663 21981 4675 21984
rect 4617 21975 4675 21981
rect 4884 21947 4942 21953
rect 4884 21913 4896 21947
rect 4930 21944 4942 21947
rect 6362 21944 6368 21956
rect 4930 21916 6368 21944
rect 4930 21913 4942 21916
rect 4884 21907 4942 21913
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 6564 21888 6592 21984
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 37461 22015 37519 22021
rect 37461 21981 37473 22015
rect 37507 22012 37519 22015
rect 38102 22012 38108 22024
rect 37507 21984 38108 22012
rect 37507 21981 37519 21984
rect 37461 21975 37519 21981
rect 38102 21972 38108 21984
rect 38160 21972 38166 22024
rect 30929 21947 30987 21953
rect 30929 21944 30941 21947
rect 30024 21916 30941 21944
rect 5994 21876 6000 21888
rect 5955 21848 6000 21876
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6546 21876 6552 21888
rect 6507 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 29546 21836 29552 21888
rect 29604 21876 29610 21888
rect 30024 21885 30052 21916
rect 30929 21913 30941 21916
rect 30975 21913 30987 21947
rect 30929 21907 30987 21913
rect 37090 21904 37096 21956
rect 37148 21944 37154 21956
rect 37148 21916 37964 21944
rect 37148 21904 37154 21916
rect 30009 21879 30067 21885
rect 30009 21876 30021 21879
rect 29604 21848 30021 21876
rect 29604 21836 29610 21848
rect 30009 21845 30021 21848
rect 30055 21845 30067 21879
rect 30009 21839 30067 21845
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 30561 21879 30619 21885
rect 30561 21876 30573 21879
rect 30524 21848 30573 21876
rect 30524 21836 30530 21848
rect 30561 21845 30573 21848
rect 30607 21845 30619 21879
rect 30561 21839 30619 21845
rect 31021 21879 31079 21885
rect 31021 21845 31033 21879
rect 31067 21876 31079 21879
rect 37734 21876 37740 21888
rect 31067 21848 37740 21876
rect 31067 21845 31079 21848
rect 31021 21839 31079 21845
rect 37734 21836 37740 21848
rect 37792 21836 37798 21888
rect 37936 21885 37964 21916
rect 37921 21879 37979 21885
rect 37921 21845 37933 21879
rect 37967 21845 37979 21879
rect 37921 21839 37979 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 3568 21644 4108 21672
rect 3568 21632 3574 21644
rect 2056 21576 4016 21604
rect 2056 21545 2084 21576
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21505 2099 21539
rect 2041 21499 2099 21505
rect 2308 21539 2366 21545
rect 2308 21505 2320 21539
rect 2354 21536 2366 21539
rect 3050 21536 3056 21548
rect 2354 21508 3056 21536
rect 2354 21505 2366 21508
rect 2308 21499 2366 21505
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 3418 21332 3424 21344
rect 3379 21304 3424 21332
rect 3418 21292 3424 21304
rect 3476 21292 3482 21344
rect 3988 21341 4016 21576
rect 4080 21400 4108 21644
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 32214 21672 32220 21684
rect 13228 21644 32220 21672
rect 13228 21632 13234 21644
rect 32214 21632 32220 21644
rect 32272 21632 32278 21684
rect 11422 21564 11428 21616
rect 11480 21604 11486 21616
rect 31018 21604 31024 21616
rect 11480 21576 31024 21604
rect 11480 21564 11486 21576
rect 31018 21564 31024 21576
rect 31076 21564 31082 21616
rect 23382 21536 23388 21548
rect 23343 21508 23388 21536
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 23750 21536 23756 21548
rect 23615 21508 23756 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 7834 21428 7840 21480
rect 7892 21468 7898 21480
rect 27982 21468 27988 21480
rect 7892 21440 27988 21468
rect 7892 21428 7898 21440
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 25866 21400 25872 21412
rect 4080 21372 25872 21400
rect 25866 21360 25872 21372
rect 25924 21360 25930 21412
rect 3973 21335 4031 21341
rect 3973 21301 3985 21335
rect 4019 21332 4031 21335
rect 6546 21332 6552 21344
rect 4019 21304 6552 21332
rect 4019 21301 4031 21304
rect 3973 21295 4031 21301
rect 6546 21292 6552 21304
rect 6604 21332 6610 21344
rect 9950 21332 9956 21344
rect 6604 21304 9956 21332
rect 6604 21292 6610 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 6362 21128 6368 21140
rect 6323 21100 6368 21128
rect 6362 21088 6368 21100
rect 6420 21088 6426 21140
rect 26602 21088 26608 21140
rect 26660 21128 26666 21140
rect 35526 21128 35532 21140
rect 26660 21100 35532 21128
rect 26660 21088 26666 21100
rect 35526 21088 35532 21100
rect 35584 21088 35590 21140
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 6546 20992 6552 21004
rect 5684 20964 6552 20992
rect 5684 20952 5690 20964
rect 6546 20952 6552 20964
rect 6604 20952 6610 21004
rect 6641 20995 6699 21001
rect 6641 20961 6653 20995
rect 6687 20992 6699 20995
rect 7282 20992 7288 21004
rect 6687 20964 7288 20992
rect 6687 20961 6699 20964
rect 6641 20955 6699 20961
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 36078 20952 36084 21004
rect 36136 20992 36142 21004
rect 37001 20995 37059 21001
rect 37001 20992 37013 20995
rect 36136 20964 37013 20992
rect 36136 20952 36142 20964
rect 37001 20961 37013 20964
rect 37047 20961 37059 20995
rect 37001 20955 37059 20961
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 6788 20896 6833 20924
rect 10428 20896 10977 20924
rect 6788 20884 6794 20896
rect 9950 20748 9956 20800
rect 10008 20788 10014 20800
rect 10428 20797 10456 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 37090 20884 37096 20936
rect 37148 20924 37154 20936
rect 37277 20927 37335 20933
rect 37277 20924 37289 20927
rect 37148 20896 37289 20924
rect 37148 20884 37154 20896
rect 37277 20893 37289 20896
rect 37323 20893 37335 20927
rect 37277 20887 37335 20893
rect 11054 20816 11060 20868
rect 11112 20856 11118 20868
rect 11210 20859 11268 20865
rect 11210 20856 11222 20859
rect 11112 20828 11222 20856
rect 11112 20816 11118 20828
rect 11210 20825 11222 20828
rect 11256 20825 11268 20859
rect 11210 20819 11268 20825
rect 10413 20791 10471 20797
rect 10413 20788 10425 20791
rect 10008 20760 10425 20788
rect 10008 20748 10014 20760
rect 10413 20757 10425 20760
rect 10459 20757 10471 20791
rect 10413 20751 10471 20757
rect 12345 20791 12403 20797
rect 12345 20757 12357 20791
rect 12391 20788 12403 20791
rect 13078 20788 13084 20800
rect 12391 20760 13084 20788
rect 12391 20757 12403 20760
rect 12345 20751 12403 20757
rect 13078 20748 13084 20760
rect 13136 20748 13142 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 6733 20587 6791 20593
rect 6733 20553 6745 20587
rect 6779 20584 6791 20587
rect 7006 20584 7012 20596
rect 6779 20556 7012 20584
rect 6779 20553 6791 20556
rect 6733 20547 6791 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 11054 20584 11060 20596
rect 10183 20556 11060 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 37734 20544 37740 20596
rect 37792 20584 37798 20596
rect 37921 20587 37979 20593
rect 37921 20584 37933 20587
rect 37792 20556 37933 20584
rect 37792 20544 37798 20556
rect 37921 20553 37933 20556
rect 37967 20553 37979 20587
rect 37921 20547 37979 20553
rect 3418 20476 3424 20528
rect 3476 20516 3482 20528
rect 6917 20519 6975 20525
rect 6917 20516 6929 20519
rect 3476 20488 6929 20516
rect 3476 20476 3482 20488
rect 6917 20485 6929 20488
rect 6963 20485 6975 20519
rect 28258 20516 28264 20528
rect 28219 20488 28264 20516
rect 6917 20479 6975 20485
rect 28258 20476 28264 20488
rect 28316 20476 28322 20528
rect 28445 20519 28503 20525
rect 28445 20485 28457 20519
rect 28491 20516 28503 20519
rect 28994 20516 29000 20528
rect 28491 20488 29000 20516
rect 28491 20485 28503 20488
rect 28445 20479 28503 20485
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20448 6883 20451
rect 6871 20420 7236 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 5994 20340 6000 20392
rect 6052 20380 6058 20392
rect 7101 20383 7159 20389
rect 7101 20380 7113 20383
rect 6052 20352 7113 20380
rect 6052 20340 6058 20352
rect 6840 20324 6868 20352
rect 7101 20349 7113 20352
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 6822 20272 6828 20324
rect 6880 20272 6886 20324
rect 7208 20312 7236 20420
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 7340 20420 10425 20448
rect 7340 20408 7346 20420
rect 10413 20417 10425 20420
rect 10459 20448 10471 20451
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 10459 20420 11529 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 11517 20417 11529 20420
rect 11563 20448 11575 20451
rect 15194 20448 15200 20460
rect 11563 20420 12434 20448
rect 15155 20420 15200 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 7432 20352 10333 20380
rect 7432 20340 7438 20352
rect 10321 20349 10333 20352
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20380 10563 20383
rect 12250 20380 12256 20392
rect 10551 20352 12256 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 8202 20312 8208 20324
rect 7208 20284 8208 20312
rect 8202 20272 8208 20284
rect 8260 20272 8266 20324
rect 12406 20312 12434 20420
rect 15194 20408 15200 20420
rect 15252 20448 15258 20460
rect 15838 20448 15844 20460
rect 15252 20420 15844 20448
rect 15252 20408 15258 20420
rect 15838 20408 15844 20420
rect 15896 20448 15902 20460
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 15896 20420 15945 20448
rect 15896 20408 15902 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 37461 20451 37519 20457
rect 37461 20417 37473 20451
rect 37507 20448 37519 20451
rect 38102 20448 38108 20460
rect 37507 20420 38108 20448
rect 37507 20417 37519 20420
rect 37461 20411 37519 20417
rect 38102 20408 38108 20420
rect 38160 20408 38166 20460
rect 15381 20315 15439 20321
rect 15381 20312 15393 20315
rect 12406 20284 15393 20312
rect 15381 20281 15393 20284
rect 15427 20312 15439 20315
rect 25038 20312 25044 20324
rect 15427 20284 25044 20312
rect 15427 20281 15439 20284
rect 15381 20275 15439 20281
rect 25038 20272 25044 20284
rect 25096 20272 25102 20324
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 6730 20000 6736 20052
rect 6788 20040 6794 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6788 20012 6837 20040
rect 6788 20000 6794 20012
rect 6825 20009 6837 20012
rect 6871 20009 6883 20043
rect 6825 20003 6883 20009
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 6972 20012 7328 20040
rect 6972 20000 6978 20012
rect 4157 19975 4215 19981
rect 4157 19941 4169 19975
rect 4203 19972 4215 19975
rect 4614 19972 4620 19984
rect 4203 19944 4620 19972
rect 4203 19941 4215 19944
rect 4157 19935 4215 19941
rect 4614 19932 4620 19944
rect 4672 19972 4678 19984
rect 4672 19944 7236 19972
rect 4672 19932 4678 19944
rect 7208 19913 7236 19944
rect 7300 19913 7328 20012
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 18012 20012 18153 20040
rect 18012 20000 18018 20012
rect 18141 20009 18153 20012
rect 18187 20009 18199 20043
rect 18141 20003 18199 20009
rect 23750 20000 23756 20052
rect 23808 20040 23814 20052
rect 26697 20043 26755 20049
rect 26697 20040 26709 20043
rect 23808 20012 26709 20040
rect 23808 20000 23814 20012
rect 26697 20009 26709 20012
rect 26743 20009 26755 20043
rect 26697 20003 26755 20009
rect 27080 20012 31064 20040
rect 13078 19972 13084 19984
rect 13039 19944 13084 19972
rect 13078 19932 13084 19944
rect 13136 19932 13142 19984
rect 17313 19975 17371 19981
rect 17313 19941 17325 19975
rect 17359 19972 17371 19975
rect 23017 19975 23075 19981
rect 17359 19944 18276 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 7193 19907 7251 19913
rect 7193 19873 7205 19907
rect 7239 19873 7251 19907
rect 7193 19867 7251 19873
rect 7285 19907 7343 19913
rect 7285 19873 7297 19907
rect 7331 19873 7343 19907
rect 7285 19867 7343 19873
rect 9950 19864 9956 19916
rect 10008 19904 10014 19916
rect 10008 19876 15516 19904
rect 10008 19864 10014 19876
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 3476 19808 4353 19836
rect 3476 19796 3482 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 7006 19836 7012 19848
rect 6967 19808 7012 19836
rect 4341 19799 4399 19805
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7374 19836 7380 19848
rect 7147 19808 7380 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 10134 19836 10140 19848
rect 10095 19808 10140 19836
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12584 19808 12725 19836
rect 12584 19796 12590 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 15488 19836 15516 19876
rect 17770 19864 17776 19916
rect 17828 19904 17834 19916
rect 18248 19913 18276 19944
rect 23017 19941 23029 19975
rect 23063 19972 23075 19975
rect 23290 19972 23296 19984
rect 23063 19944 23296 19972
rect 23063 19941 23075 19944
rect 23017 19935 23075 19941
rect 23290 19932 23296 19944
rect 23348 19932 23354 19984
rect 27080 19972 27108 20012
rect 27246 19972 27252 19984
rect 26206 19944 27108 19972
rect 27207 19944 27252 19972
rect 18233 19907 18291 19913
rect 17828 19876 18092 19904
rect 17828 19864 17834 19876
rect 15930 19836 15936 19848
rect 15488 19808 15936 19836
rect 9950 19768 9956 19780
rect 9911 19740 9956 19768
rect 9950 19728 9956 19740
rect 10008 19728 10014 19780
rect 12618 19728 12624 19780
rect 12676 19768 12682 19780
rect 12897 19771 12955 19777
rect 12897 19768 12909 19771
rect 12676 19740 12909 19768
rect 12676 19728 12682 19740
rect 12897 19737 12909 19740
rect 12943 19737 12955 19771
rect 12897 19731 12955 19737
rect 15488 19712 15516 19808
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18064 19836 18092 19876
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 19978 19904 19984 19916
rect 18279 19876 19984 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 26050 19904 26056 19916
rect 25096 19876 26056 19904
rect 25096 19864 25102 19876
rect 26050 19864 26056 19876
rect 26108 19904 26114 19916
rect 26206 19904 26234 19944
rect 27246 19932 27252 19944
rect 27304 19932 27310 19984
rect 30190 19904 30196 19916
rect 26108 19876 26234 19904
rect 26896 19876 30196 19904
rect 26108 19864 26114 19876
rect 22465 19839 22523 19845
rect 22465 19836 22477 19839
rect 18064 19808 22477 19836
rect 22465 19805 22477 19808
rect 22511 19836 22523 19839
rect 23017 19839 23075 19845
rect 23017 19836 23029 19839
rect 22511 19808 23029 19836
rect 22511 19805 22523 19808
rect 22465 19799 22523 19805
rect 23017 19805 23029 19808
rect 23063 19805 23075 19839
rect 23017 19799 23075 19805
rect 23106 19796 23112 19848
rect 23164 19836 23170 19848
rect 26896 19845 26924 19876
rect 30190 19864 30196 19876
rect 30248 19904 30254 19916
rect 30377 19907 30435 19913
rect 30377 19904 30389 19907
rect 30248 19876 30389 19904
rect 30248 19864 30254 19876
rect 30377 19873 30389 19876
rect 30423 19873 30435 19907
rect 30377 19867 30435 19873
rect 23293 19839 23351 19845
rect 23293 19836 23305 19839
rect 23164 19808 23305 19836
rect 23164 19796 23170 19808
rect 23293 19805 23305 19808
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 26881 19839 26939 19845
rect 26881 19805 26893 19839
rect 26927 19805 26939 19839
rect 26881 19799 26939 19805
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 31036 19845 31064 20012
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 27304 19808 30113 19836
rect 27304 19796 27310 19808
rect 30101 19805 30113 19808
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 30837 19839 30895 19845
rect 30837 19805 30849 19839
rect 30883 19805 30895 19839
rect 30837 19799 30895 19805
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19836 31079 19839
rect 31481 19839 31539 19845
rect 31481 19836 31493 19839
rect 31067 19808 31493 19836
rect 31067 19805 31079 19808
rect 31021 19799 31079 19805
rect 31481 19805 31493 19808
rect 31527 19836 31539 19839
rect 33226 19836 33232 19848
rect 31527 19808 33232 19836
rect 31527 19805 31539 19808
rect 31481 19799 31539 19805
rect 16200 19771 16258 19777
rect 16200 19737 16212 19771
rect 16246 19768 16258 19771
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 16246 19740 17785 19768
rect 16246 19737 16258 19740
rect 16200 19731 16258 19737
rect 17773 19737 17785 19740
rect 17819 19737 17831 19771
rect 17773 19731 17831 19737
rect 27065 19771 27123 19777
rect 27065 19737 27077 19771
rect 27111 19768 27123 19771
rect 27338 19768 27344 19780
rect 27111 19740 27344 19768
rect 27111 19737 27123 19740
rect 27065 19731 27123 19737
rect 27338 19728 27344 19740
rect 27396 19728 27402 19780
rect 30116 19768 30144 19799
rect 30852 19768 30880 19799
rect 33226 19796 33232 19808
rect 33284 19796 33290 19848
rect 30116 19740 30880 19768
rect 8202 19660 8208 19712
rect 8260 19700 8266 19712
rect 12529 19703 12587 19709
rect 12529 19700 12541 19703
rect 8260 19672 12541 19700
rect 8260 19660 8266 19672
rect 12529 19669 12541 19672
rect 12575 19669 12587 19703
rect 12802 19700 12808 19712
rect 12763 19672 12808 19700
rect 12529 19663 12587 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 15470 19700 15476 19712
rect 15431 19672 15476 19700
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 23198 19700 23204 19712
rect 23159 19672 23204 19700
rect 23198 19660 23204 19672
rect 23256 19660 23262 19712
rect 26970 19660 26976 19712
rect 27028 19700 27034 19712
rect 30926 19700 30932 19712
rect 27028 19672 27073 19700
rect 30887 19672 30932 19700
rect 27028 19660 27034 19672
rect 30926 19660 30932 19672
rect 30984 19660 30990 19712
rect 34330 19660 34336 19712
rect 34388 19700 34394 19712
rect 35894 19700 35900 19712
rect 34388 19672 35900 19700
rect 34388 19660 34394 19672
rect 35894 19660 35900 19672
rect 35952 19660 35958 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 12250 19496 12256 19508
rect 12211 19468 12256 19496
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 19978 19496 19984 19508
rect 19939 19468 19984 19496
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 26142 19456 26148 19508
rect 26200 19496 26206 19508
rect 26237 19499 26295 19505
rect 26237 19496 26249 19499
rect 26200 19468 26249 19496
rect 26200 19456 26206 19468
rect 26237 19465 26249 19468
rect 26283 19496 26295 19499
rect 26970 19496 26976 19508
rect 26283 19468 26976 19496
rect 26283 19465 26295 19468
rect 26237 19459 26295 19465
rect 26970 19456 26976 19468
rect 27028 19456 27034 19508
rect 30190 19496 30196 19508
rect 30151 19468 30196 19496
rect 30190 19456 30196 19468
rect 30248 19456 30254 19508
rect 33226 19456 33232 19508
rect 33284 19496 33290 19508
rect 33413 19499 33471 19505
rect 33413 19496 33425 19499
rect 33284 19468 33425 19496
rect 33284 19456 33290 19468
rect 33413 19465 33425 19468
rect 33459 19465 33471 19499
rect 34330 19496 34336 19508
rect 34291 19468 34336 19496
rect 33413 19459 33471 19465
rect 34330 19456 34336 19468
rect 34388 19456 34394 19508
rect 35894 19456 35900 19508
rect 35952 19496 35958 19508
rect 36265 19499 36323 19505
rect 36265 19496 36277 19499
rect 35952 19468 36277 19496
rect 35952 19456 35958 19468
rect 36265 19465 36277 19468
rect 36311 19465 36323 19499
rect 36265 19459 36323 19465
rect 12526 19428 12532 19440
rect 12452 19400 12532 19428
rect 12452 19369 12480 19400
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 19886 19428 19892 19440
rect 19799 19400 19892 19428
rect 19886 19388 19892 19400
rect 19944 19428 19950 19440
rect 23750 19428 23756 19440
rect 19944 19400 22094 19428
rect 19944 19388 19950 19400
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13078 19360 13084 19372
rect 12759 19332 13084 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 17828 19332 19625 19360
rect 17828 19320 17834 19332
rect 19613 19329 19625 19332
rect 19659 19329 19671 19363
rect 19794 19360 19800 19372
rect 19755 19332 19800 19360
rect 19613 19323 19671 19329
rect 19794 19320 19800 19332
rect 19852 19360 19858 19372
rect 20990 19360 20996 19372
rect 19852 19332 20996 19360
rect 19852 19320 19858 19332
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 22066 19360 22094 19400
rect 22388 19400 23756 19428
rect 22388 19360 22416 19400
rect 23750 19388 23756 19400
rect 23808 19388 23814 19440
rect 27125 19431 27183 19437
rect 27125 19428 27137 19431
rect 26160 19400 27137 19428
rect 22066 19332 22416 19360
rect 23106 19320 23112 19372
rect 23164 19360 23170 19372
rect 26160 19369 26188 19400
rect 27125 19397 27137 19400
rect 27171 19428 27183 19431
rect 27246 19428 27252 19440
rect 27171 19400 27252 19428
rect 27171 19397 27183 19400
rect 27125 19391 27183 19397
rect 27246 19388 27252 19400
rect 27304 19388 27310 19440
rect 27338 19388 27344 19440
rect 27396 19428 27402 19440
rect 34698 19428 34704 19440
rect 27396 19400 27441 19428
rect 29656 19400 34704 19428
rect 27396 19388 27402 19400
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 23164 19332 26157 19360
rect 23164 19320 23170 19332
rect 26145 19329 26157 19332
rect 26191 19329 26203 19363
rect 26145 19323 26203 19329
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19360 26479 19363
rect 27356 19360 27384 19388
rect 26467 19332 27384 19360
rect 26467 19329 26479 19332
rect 26421 19323 26479 19329
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12544 19224 12572 19255
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 12676 19264 12721 19292
rect 12676 19252 12682 19264
rect 28258 19252 28264 19304
rect 28316 19292 28322 19304
rect 29656 19301 29684 19400
rect 30926 19320 30932 19372
rect 30984 19360 30990 19372
rect 31588 19369 31616 19400
rect 34698 19388 34704 19400
rect 34756 19428 34762 19440
rect 36280 19428 36308 19459
rect 37461 19431 37519 19437
rect 37461 19428 37473 19431
rect 34756 19400 34928 19428
rect 36280 19400 37473 19428
rect 34756 19388 34762 19400
rect 31306 19363 31364 19369
rect 31306 19360 31318 19363
rect 30984 19332 31318 19360
rect 30984 19320 30990 19332
rect 31306 19329 31318 19332
rect 31352 19329 31364 19363
rect 31306 19323 31364 19329
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19329 31631 19363
rect 31573 19323 31631 19329
rect 33226 19320 33232 19372
rect 33284 19360 33290 19372
rect 34149 19363 34207 19369
rect 34149 19360 34161 19363
rect 33284 19332 34161 19360
rect 33284 19320 33290 19332
rect 34149 19329 34161 19332
rect 34195 19329 34207 19363
rect 34149 19323 34207 19329
rect 34425 19363 34483 19369
rect 34425 19329 34437 19363
rect 34471 19360 34483 19363
rect 34790 19360 34796 19372
rect 34471 19332 34796 19360
rect 34471 19329 34483 19332
rect 34425 19323 34483 19329
rect 34790 19320 34796 19332
rect 34848 19320 34854 19372
rect 34900 19369 34928 19400
rect 37461 19397 37473 19400
rect 37507 19397 37519 19431
rect 37461 19391 37519 19397
rect 34885 19363 34943 19369
rect 34885 19329 34897 19363
rect 34931 19329 34943 19363
rect 35141 19363 35199 19369
rect 35141 19360 35153 19363
rect 34885 19323 34943 19329
rect 34992 19332 35153 19360
rect 29641 19295 29699 19301
rect 29641 19292 29653 19295
rect 28316 19264 29653 19292
rect 28316 19252 28322 19264
rect 29641 19261 29653 19264
rect 29687 19261 29699 19295
rect 29641 19255 29699 19261
rect 33965 19295 34023 19301
rect 33965 19261 33977 19295
rect 34011 19292 34023 19295
rect 34992 19292 35020 19332
rect 35141 19329 35153 19332
rect 35187 19329 35199 19363
rect 35141 19323 35199 19329
rect 37645 19363 37703 19369
rect 37645 19329 37657 19363
rect 37691 19360 37703 19363
rect 38838 19360 38844 19372
rect 37691 19332 38844 19360
rect 37691 19329 37703 19332
rect 37645 19323 37703 19329
rect 38838 19320 38844 19332
rect 38896 19320 38902 19372
rect 34011 19264 35020 19292
rect 37277 19295 37335 19301
rect 34011 19261 34023 19264
rect 33965 19255 34023 19261
rect 37277 19261 37289 19295
rect 37323 19292 37335 19295
rect 38562 19292 38568 19304
rect 37323 19264 38568 19292
rect 37323 19261 37335 19264
rect 37277 19255 37335 19261
rect 38562 19252 38568 19264
rect 38620 19252 38626 19304
rect 12802 19224 12808 19236
rect 12544 19196 12808 19224
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 20162 19224 20168 19236
rect 20123 19196 20168 19224
rect 20162 19184 20168 19196
rect 20220 19184 20226 19236
rect 23198 19184 23204 19236
rect 23256 19224 23262 19236
rect 26142 19224 26148 19236
rect 23256 19196 26148 19224
rect 23256 19184 23262 19196
rect 26142 19184 26148 19196
rect 26200 19224 26206 19236
rect 26200 19196 27200 19224
rect 26200 19184 26206 19196
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 25682 19156 25688 19168
rect 20312 19128 25688 19156
rect 20312 19116 20318 19128
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 26234 19116 26240 19168
rect 26292 19156 26298 19168
rect 26421 19159 26479 19165
rect 26421 19156 26433 19159
rect 26292 19128 26433 19156
rect 26292 19116 26298 19128
rect 26421 19125 26433 19128
rect 26467 19125 26479 19159
rect 26421 19119 26479 19125
rect 26510 19116 26516 19168
rect 26568 19156 26574 19168
rect 27172 19165 27200 19196
rect 26973 19159 27031 19165
rect 26973 19156 26985 19159
rect 26568 19128 26985 19156
rect 26568 19116 26574 19128
rect 26973 19125 26985 19128
rect 27019 19125 27031 19159
rect 26973 19119 27031 19125
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19125 27215 19159
rect 27157 19119 27215 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 19797 18955 19855 18961
rect 19797 18921 19809 18955
rect 19843 18952 19855 18955
rect 19886 18952 19892 18964
rect 19843 18924 19892 18952
rect 19843 18921 19855 18924
rect 19797 18915 19855 18921
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 23106 18952 23112 18964
rect 23067 18924 23112 18952
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 34698 18952 34704 18964
rect 34659 18924 34704 18952
rect 34698 18912 34704 18924
rect 34756 18912 34762 18964
rect 5166 18844 5172 18896
rect 5224 18884 5230 18896
rect 24210 18884 24216 18896
rect 5224 18856 24216 18884
rect 5224 18844 5230 18856
rect 24210 18844 24216 18856
rect 24268 18844 24274 18896
rect 26329 18887 26387 18893
rect 26329 18853 26341 18887
rect 26375 18884 26387 18887
rect 26418 18884 26424 18896
rect 26375 18856 26424 18884
rect 26375 18853 26387 18856
rect 26329 18847 26387 18853
rect 26418 18844 26424 18856
rect 26476 18844 26482 18896
rect 37366 18884 37372 18896
rect 35866 18856 37372 18884
rect 23198 18816 23204 18828
rect 23032 18788 23204 18816
rect 5718 18708 5724 18760
rect 5776 18748 5782 18760
rect 5776 18720 22094 18748
rect 5776 18708 5782 18720
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 18874 18680 18880 18692
rect 18104 18652 18880 18680
rect 18104 18640 18110 18652
rect 18874 18640 18880 18652
rect 18932 18680 18938 18692
rect 19794 18689 19800 18692
rect 19781 18683 19800 18689
rect 18932 18652 19656 18680
rect 18932 18640 18938 18652
rect 3142 18572 3148 18624
rect 3200 18612 3206 18624
rect 19426 18612 19432 18624
rect 3200 18584 19432 18612
rect 3200 18572 3206 18584
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 19628 18621 19656 18652
rect 19781 18649 19793 18683
rect 19781 18643 19800 18649
rect 19794 18640 19800 18643
rect 19852 18640 19858 18692
rect 19978 18680 19984 18692
rect 19939 18652 19984 18680
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 22066 18680 22094 18720
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 23032 18757 23060 18788
rect 23198 18776 23204 18788
rect 23256 18776 23262 18828
rect 25777 18819 25835 18825
rect 25777 18785 25789 18819
rect 25823 18816 25835 18819
rect 26050 18816 26056 18828
rect 25823 18788 26056 18816
rect 25823 18785 25835 18788
rect 25777 18779 25835 18785
rect 26050 18776 26056 18788
rect 26108 18816 26114 18828
rect 26513 18819 26571 18825
rect 26513 18816 26525 18819
rect 26108 18788 26525 18816
rect 26108 18776 26114 18788
rect 26513 18785 26525 18788
rect 26559 18785 26571 18819
rect 26513 18779 26571 18785
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22428 18720 23029 18748
rect 22428 18708 22434 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23290 18748 23296 18760
rect 23251 18720 23296 18748
rect 23017 18711 23075 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 26234 18708 26240 18760
rect 26292 18748 26298 18760
rect 26292 18720 26337 18748
rect 26292 18708 26298 18720
rect 25590 18680 25596 18692
rect 22066 18652 25596 18680
rect 25590 18640 25596 18652
rect 25648 18640 25654 18692
rect 25682 18640 25688 18692
rect 25740 18680 25746 18692
rect 35866 18680 35894 18856
rect 37366 18844 37372 18856
rect 37424 18844 37430 18896
rect 37461 18751 37519 18757
rect 37461 18717 37473 18751
rect 37507 18748 37519 18751
rect 38102 18748 38108 18760
rect 37507 18720 38108 18748
rect 37507 18717 37519 18720
rect 37461 18711 37519 18717
rect 38102 18708 38108 18720
rect 38160 18708 38166 18760
rect 25740 18652 35894 18680
rect 25740 18640 25746 18652
rect 19613 18615 19671 18621
rect 19613 18581 19625 18615
rect 19659 18581 19671 18615
rect 23474 18612 23480 18624
rect 23435 18584 23480 18612
rect 19613 18575 19671 18581
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 37918 18612 37924 18624
rect 26292 18584 26337 18612
rect 37879 18584 37924 18612
rect 26292 18572 26298 18584
rect 37918 18572 37924 18584
rect 37976 18572 37982 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 2961 18411 3019 18417
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 3050 18408 3056 18420
rect 3007 18380 3056 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 17773 18411 17831 18417
rect 17773 18377 17785 18411
rect 17819 18408 17831 18411
rect 17954 18408 17960 18420
rect 17819 18380 17960 18408
rect 17819 18377 17831 18380
rect 17773 18371 17831 18377
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 21082 18368 21088 18420
rect 21140 18408 21146 18420
rect 37274 18408 37280 18420
rect 21140 18380 37280 18408
rect 21140 18368 21146 18380
rect 37274 18368 37280 18380
rect 37332 18368 37338 18420
rect 3145 18275 3203 18281
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3234 18272 3240 18284
rect 3191 18244 3240 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 17678 18272 17684 18284
rect 17639 18244 17684 18272
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 18046 18272 18052 18284
rect 17911 18244 18052 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 4614 18204 4620 18216
rect 3467 18176 4620 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 3329 18071 3387 18077
rect 3329 18037 3341 18071
rect 3375 18068 3387 18071
rect 3970 18068 3976 18080
rect 3375 18040 3976 18068
rect 3375 18037 3387 18040
rect 3329 18031 3387 18037
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 3234 17864 3240 17876
rect 3195 17836 3240 17864
rect 3234 17824 3240 17836
rect 3292 17824 3298 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 8297 17867 8355 17873
rect 8297 17864 8309 17867
rect 7432 17836 8309 17864
rect 7432 17824 7438 17836
rect 8297 17833 8309 17836
rect 8343 17833 8355 17867
rect 8297 17827 8355 17833
rect 9769 17867 9827 17873
rect 9769 17833 9781 17867
rect 9815 17864 9827 17867
rect 15194 17864 15200 17876
rect 9815 17836 15200 17864
rect 9815 17833 9827 17836
rect 9769 17827 9827 17833
rect 4157 17731 4215 17737
rect 3068 17700 3924 17728
rect 3068 17669 3096 17700
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 3283 17632 3832 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 3804 17536 3832 17632
rect 3786 17524 3792 17536
rect 3747 17496 3792 17524
rect 3786 17484 3792 17496
rect 3844 17484 3850 17536
rect 3896 17524 3924 17700
rect 4157 17697 4169 17731
rect 4203 17728 4215 17731
rect 4614 17728 4620 17740
rect 4203 17700 4620 17728
rect 4203 17697 4215 17700
rect 4157 17691 4215 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 7374 17660 7380 17672
rect 4028 17632 7380 17660
rect 4028 17620 4034 17632
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 8202 17660 8208 17672
rect 8163 17632 8208 17660
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 8536 17632 8953 17660
rect 8536 17620 8542 17632
rect 8941 17629 8953 17632
rect 8987 17660 8999 17663
rect 9784 17660 9812 17827
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 22370 17864 22376 17876
rect 22331 17836 22376 17864
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 34606 17864 34612 17876
rect 22848 17836 34612 17864
rect 21542 17756 21548 17808
rect 21600 17796 21606 17808
rect 22848 17796 22876 17836
rect 34606 17824 34612 17836
rect 34664 17824 34670 17876
rect 21600 17768 22876 17796
rect 21600 17756 21606 17768
rect 8987 17632 9812 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 23474 17620 23480 17672
rect 23532 17669 23538 17672
rect 23532 17660 23544 17669
rect 23753 17663 23811 17669
rect 23532 17632 23577 17660
rect 23532 17623 23544 17632
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 38102 17660 38108 17672
rect 23799 17632 24532 17660
rect 38063 17632 38108 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 23532 17620 23538 17623
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 23382 17592 23388 17604
rect 12952 17564 23388 17592
rect 12952 17552 12958 17564
rect 23382 17552 23388 17564
rect 23440 17552 23446 17604
rect 4890 17524 4896 17536
rect 3896 17496 4896 17524
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 4948 17496 9137 17524
rect 4948 17484 4954 17496
rect 9125 17493 9137 17496
rect 9171 17524 9183 17527
rect 12434 17524 12440 17536
rect 9171 17496 12440 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 24504 17533 24532 17632
rect 38102 17620 38108 17632
rect 38160 17620 38166 17672
rect 24489 17527 24547 17533
rect 24489 17493 24501 17527
rect 24535 17524 24547 17527
rect 28258 17524 28264 17536
rect 24535 17496 28264 17524
rect 24535 17493 24547 17496
rect 24489 17487 24547 17493
rect 28258 17484 28264 17496
rect 28316 17484 28322 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8478 17320 8484 17332
rect 8439 17292 8484 17320
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 12710 17320 12716 17332
rect 12268 17292 12716 17320
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7653 17187 7711 17193
rect 7653 17184 7665 17187
rect 7432 17156 7665 17184
rect 7432 17144 7438 17156
rect 7653 17153 7665 17156
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 8496 17184 8524 17280
rect 12268 17193 12296 17292
rect 12710 17280 12716 17292
rect 12768 17320 12774 17332
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 12768 17292 13001 17320
rect 12768 17280 12774 17292
rect 12989 17289 13001 17292
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 13412 17292 17816 17320
rect 13412 17280 13418 17292
rect 17678 17252 17684 17264
rect 12728 17224 17684 17252
rect 7883 17156 8524 17184
rect 12253 17187 12311 17193
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12728 17184 12756 17224
rect 17678 17212 17684 17224
rect 17736 17212 17742 17264
rect 17788 17252 17816 17292
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 20496 17292 35894 17320
rect 20496 17280 20502 17292
rect 32122 17252 32128 17264
rect 17788 17224 32128 17252
rect 32122 17212 32128 17224
rect 32180 17212 32186 17264
rect 34238 17252 34244 17264
rect 32232 17224 34244 17252
rect 12492 17156 12756 17184
rect 12492 17144 12498 17156
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12860 17156 13185 17184
rect 12860 17144 12866 17156
rect 13173 17153 13185 17156
rect 13219 17184 13231 17187
rect 17770 17184 17776 17196
rect 13219 17156 17776 17184
rect 13219 17153 13231 17156
rect 13173 17147 13231 17153
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 32232 17184 32260 17224
rect 34238 17212 34244 17224
rect 34296 17212 34302 17264
rect 20588 17156 32260 17184
rect 20588 17144 20594 17156
rect 33686 17144 33692 17196
rect 33744 17184 33750 17196
rect 33873 17187 33931 17193
rect 33873 17184 33885 17187
rect 33744 17156 33885 17184
rect 33744 17144 33750 17156
rect 33873 17153 33885 17156
rect 33919 17153 33931 17187
rect 33873 17147 33931 17153
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7558 17116 7564 17128
rect 7064 17088 7564 17116
rect 7064 17076 7070 17088
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 13357 17119 13415 17125
rect 13357 17116 13369 17119
rect 12584 17088 13369 17116
rect 12584 17076 12590 17088
rect 13357 17085 13369 17088
rect 13403 17085 13415 17119
rect 34146 17116 34152 17128
rect 34107 17088 34152 17116
rect 13357 17079 13415 17085
rect 34146 17076 34152 17088
rect 34204 17076 34210 17128
rect 35866 17048 35894 17292
rect 37550 17048 37556 17060
rect 35866 17020 37556 17048
rect 37550 17008 37556 17020
rect 37608 17008 37614 17060
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 7377 16983 7435 16989
rect 7377 16980 7389 16983
rect 7340 16952 7389 16980
rect 7340 16940 7346 16952
rect 7377 16949 7389 16952
rect 7423 16949 7435 16983
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 7377 16943 7435 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 4614 16736 4620 16788
rect 4672 16776 4678 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 4672 16748 7021 16776
rect 4672 16736 4678 16748
rect 7009 16745 7021 16748
rect 7055 16776 7067 16779
rect 7742 16776 7748 16788
rect 7055 16748 7748 16776
rect 7055 16745 7067 16748
rect 7009 16739 7067 16745
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 12802 16776 12808 16788
rect 12483 16748 12808 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 31665 16643 31723 16649
rect 17828 16612 17908 16640
rect 17828 16600 17834 16612
rect 12250 16572 12256 16584
rect 12211 16544 12256 16572
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12584 16544 12629 16572
rect 12584 16532 12590 16544
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 15194 16572 15200 16584
rect 14516 16544 15200 16572
rect 14516 16532 14522 16544
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 17678 16532 17684 16584
rect 17736 16581 17742 16584
rect 17880 16581 17908 16612
rect 31665 16609 31677 16643
rect 31711 16640 31723 16643
rect 31938 16640 31944 16652
rect 31711 16612 31944 16640
rect 31711 16609 31723 16612
rect 31665 16603 31723 16609
rect 31938 16600 31944 16612
rect 31996 16600 32002 16652
rect 17736 16572 17745 16581
rect 17865 16575 17923 16581
rect 17736 16544 17781 16572
rect 17736 16535 17745 16544
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 31386 16572 31392 16584
rect 31347 16544 31392 16572
rect 17865 16535 17923 16541
rect 17736 16532 17742 16535
rect 31386 16532 31392 16544
rect 31444 16532 31450 16584
rect 7190 16504 7196 16516
rect 7151 16476 7196 16504
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 14734 16464 14740 16516
rect 14792 16504 14798 16516
rect 18782 16504 18788 16516
rect 14792 16476 18788 16504
rect 14792 16464 14798 16476
rect 18782 16464 18788 16476
rect 18840 16464 18846 16516
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6993 16439 7051 16445
rect 6993 16405 7005 16439
rect 7039 16436 7051 16439
rect 8202 16436 8208 16448
rect 7039 16408 8208 16436
rect 7039 16405 7051 16408
rect 6993 16399 7051 16405
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 17770 16436 17776 16448
rect 17731 16408 17776 16436
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 37458 16436 37464 16448
rect 37419 16408 37464 16436
rect 37458 16396 37464 16408
rect 37516 16396 37522 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 29917 16235 29975 16241
rect 29917 16201 29929 16235
rect 29963 16232 29975 16235
rect 30374 16232 30380 16244
rect 29963 16204 30380 16232
rect 29963 16201 29975 16204
rect 29917 16195 29975 16201
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 30558 16192 30564 16244
rect 30616 16232 30622 16244
rect 30653 16235 30711 16241
rect 30653 16232 30665 16235
rect 30616 16204 30665 16232
rect 30616 16192 30622 16204
rect 30653 16201 30665 16204
rect 30699 16201 30711 16235
rect 30653 16195 30711 16201
rect 33965 16235 34023 16241
rect 33965 16201 33977 16235
rect 34011 16232 34023 16235
rect 34146 16232 34152 16244
rect 34011 16204 34152 16232
rect 34011 16201 34023 16204
rect 33965 16195 34023 16201
rect 34146 16192 34152 16204
rect 34204 16192 34210 16244
rect 34425 16235 34483 16241
rect 34425 16201 34437 16235
rect 34471 16232 34483 16235
rect 38010 16232 38016 16244
rect 34471 16204 38016 16232
rect 34471 16201 34483 16204
rect 34425 16195 34483 16201
rect 38010 16192 38016 16204
rect 38068 16192 38074 16244
rect 4890 16164 4896 16176
rect 4264 16136 4896 16164
rect 4264 16105 4292 16136
rect 4890 16124 4896 16136
rect 4948 16124 4954 16176
rect 25498 16124 25504 16176
rect 25556 16164 25562 16176
rect 37458 16164 37464 16176
rect 25556 16136 37464 16164
rect 25556 16124 25562 16136
rect 37458 16124 37464 16136
rect 37516 16164 37522 16176
rect 37737 16167 37795 16173
rect 37737 16164 37749 16167
rect 37516 16136 37749 16164
rect 37516 16124 37522 16136
rect 37737 16133 37749 16136
rect 37783 16133 37795 16167
rect 37737 16127 37795 16133
rect 37921 16167 37979 16173
rect 37921 16133 37933 16167
rect 37967 16164 37979 16167
rect 38746 16164 38752 16176
rect 37967 16136 38752 16164
rect 37967 16133 37979 16136
rect 37921 16127 37979 16133
rect 38746 16124 38752 16136
rect 38804 16124 38810 16176
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 4249 16059 4307 16065
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 6822 16096 6828 16108
rect 4479 16068 6828 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 17770 16056 17776 16108
rect 17828 16096 17834 16108
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 17828 16068 18705 16096
rect 17828 16056 17834 16068
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 18874 16096 18880 16108
rect 18835 16068 18880 16096
rect 18693 16059 18751 16065
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 20162 16096 20168 16108
rect 19015 16068 20168 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 28994 16056 29000 16108
rect 29052 16096 29058 16108
rect 29825 16099 29883 16105
rect 29825 16096 29837 16099
rect 29052 16068 29837 16096
rect 29052 16056 29058 16068
rect 29825 16065 29837 16068
rect 29871 16065 29883 16099
rect 30558 16096 30564 16108
rect 30519 16068 30564 16096
rect 29825 16059 29883 16065
rect 30558 16056 30564 16068
rect 30616 16056 30622 16108
rect 34333 16099 34391 16105
rect 34333 16065 34345 16099
rect 34379 16065 34391 16099
rect 34333 16059 34391 16065
rect 3970 15852 3976 15904
rect 4028 15892 4034 15904
rect 4433 15895 4491 15901
rect 4433 15892 4445 15895
rect 4028 15864 4445 15892
rect 4028 15852 4034 15864
rect 4433 15861 4445 15864
rect 4479 15861 4491 15895
rect 18506 15892 18512 15904
rect 18467 15864 18512 15892
rect 4433 15855 4491 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 27246 15852 27252 15904
rect 27304 15892 27310 15904
rect 33413 15895 33471 15901
rect 33413 15892 33425 15895
rect 27304 15864 33425 15892
rect 27304 15852 27310 15864
rect 33413 15861 33425 15864
rect 33459 15892 33471 15895
rect 34348 15892 34376 16059
rect 34609 16031 34667 16037
rect 34609 15997 34621 16031
rect 34655 16028 34667 16031
rect 35342 16028 35348 16040
rect 34655 16000 35348 16028
rect 34655 15997 34667 16000
rect 34609 15991 34667 15997
rect 35342 15988 35348 16000
rect 35400 15988 35406 16040
rect 33459 15864 34376 15892
rect 33459 15861 33471 15864
rect 33413 15855 33471 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3786 15648 3792 15700
rect 3844 15688 3850 15700
rect 4157 15691 4215 15697
rect 4157 15688 4169 15691
rect 3844 15660 4169 15688
rect 3844 15648 3850 15660
rect 4157 15657 4169 15660
rect 4203 15657 4215 15691
rect 4157 15651 4215 15657
rect 12437 15691 12495 15697
rect 12437 15657 12449 15691
rect 12483 15688 12495 15691
rect 12526 15688 12532 15700
rect 12483 15660 12532 15688
rect 12483 15657 12495 15660
rect 12437 15651 12495 15657
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 20162 15648 20168 15700
rect 20220 15688 20226 15700
rect 20625 15691 20683 15697
rect 20625 15688 20637 15691
rect 20220 15660 20637 15688
rect 20220 15648 20226 15660
rect 20625 15657 20637 15660
rect 20671 15657 20683 15691
rect 27709 15691 27767 15697
rect 27709 15688 27721 15691
rect 20625 15651 20683 15657
rect 25792 15660 27721 15688
rect 15470 15552 15476 15564
rect 12406 15524 15476 15552
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10643 15456 11069 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 11057 15453 11069 15456
rect 11103 15484 11115 15487
rect 12406 15484 12434 15524
rect 15470 15512 15476 15524
rect 15528 15552 15534 15564
rect 25792 15561 25820 15660
rect 27709 15657 27721 15660
rect 27755 15688 27767 15691
rect 28258 15688 28264 15700
rect 27755 15660 28264 15688
rect 27755 15657 27767 15660
rect 27709 15651 27767 15657
rect 28258 15648 28264 15660
rect 28316 15648 28322 15700
rect 30653 15691 30711 15697
rect 30653 15657 30665 15691
rect 30699 15688 30711 15691
rect 31386 15688 31392 15700
rect 30699 15660 31392 15688
rect 30699 15657 30711 15660
rect 30653 15651 30711 15657
rect 31386 15648 31392 15660
rect 31444 15648 31450 15700
rect 32493 15691 32551 15697
rect 32493 15688 32505 15691
rect 31680 15660 32505 15688
rect 27157 15623 27215 15629
rect 27157 15589 27169 15623
rect 27203 15620 27215 15623
rect 27338 15620 27344 15632
rect 27203 15592 27344 15620
rect 27203 15589 27215 15592
rect 27157 15583 27215 15589
rect 27338 15580 27344 15592
rect 27396 15580 27402 15632
rect 31680 15629 31708 15660
rect 32493 15657 32505 15660
rect 32539 15688 32551 15691
rect 32582 15688 32588 15700
rect 32539 15660 32588 15688
rect 32539 15657 32551 15660
rect 32493 15651 32551 15657
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 34790 15688 34796 15700
rect 34751 15660 34796 15688
rect 34790 15648 34796 15660
rect 34848 15648 34854 15700
rect 35342 15648 35348 15700
rect 35400 15688 35406 15700
rect 37921 15691 37979 15697
rect 37921 15688 37933 15691
rect 35400 15660 37933 15688
rect 35400 15648 35406 15660
rect 37921 15657 37933 15660
rect 37967 15657 37979 15691
rect 37921 15651 37979 15657
rect 31665 15623 31723 15629
rect 31665 15589 31677 15623
rect 31711 15589 31723 15623
rect 31665 15583 31723 15589
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 15528 15524 18705 15552
rect 15528 15512 15534 15524
rect 18693 15521 18705 15524
rect 18739 15552 18751 15555
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 18739 15524 19257 15552
rect 18739 15521 18751 15524
rect 18693 15515 18751 15521
rect 19245 15521 19257 15524
rect 19291 15521 19303 15555
rect 19245 15515 19303 15521
rect 25777 15555 25835 15561
rect 25777 15521 25789 15555
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 29178 15512 29184 15564
rect 29236 15552 29242 15564
rect 31941 15555 31999 15561
rect 31941 15552 31953 15555
rect 29236 15524 31953 15552
rect 29236 15512 29242 15524
rect 11103 15456 12434 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 19501 15487 19559 15493
rect 19501 15484 19513 15487
rect 18564 15456 19513 15484
rect 18564 15444 18570 15456
rect 19501 15453 19513 15456
rect 19547 15453 19559 15487
rect 19501 15447 19559 15453
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 30484 15493 30512 15524
rect 31941 15521 31953 15524
rect 31987 15552 31999 15555
rect 35360 15552 35388 15648
rect 31987 15524 35388 15552
rect 31987 15521 31999 15524
rect 31941 15515 31999 15521
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 20404 15456 29745 15484
rect 20404 15444 20410 15456
rect 29733 15453 29745 15456
rect 29779 15484 29791 15487
rect 30285 15487 30343 15493
rect 30285 15484 30297 15487
rect 29779 15456 30297 15484
rect 29779 15453 29791 15456
rect 29733 15447 29791 15453
rect 30285 15453 30297 15456
rect 30331 15453 30343 15487
rect 30285 15447 30343 15453
rect 30469 15487 30527 15493
rect 30469 15453 30481 15487
rect 30515 15453 30527 15487
rect 30469 15447 30527 15453
rect 34790 15444 34796 15496
rect 34848 15484 34854 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34848 15456 34897 15484
rect 34848 15444 34854 15456
rect 34885 15453 34897 15456
rect 34931 15484 34943 15487
rect 35345 15487 35403 15493
rect 35345 15484 35357 15487
rect 34931 15456 35357 15484
rect 34931 15453 34943 15456
rect 34885 15447 34943 15453
rect 35345 15453 35357 15456
rect 35391 15453 35403 15487
rect 35345 15447 35403 15453
rect 36541 15487 36599 15493
rect 36541 15453 36553 15487
rect 36587 15484 36599 15487
rect 37182 15484 37188 15496
rect 36587 15456 37188 15484
rect 36587 15453 36599 15456
rect 36541 15447 36599 15453
rect 37182 15444 37188 15456
rect 37240 15444 37246 15496
rect 38010 15484 38016 15496
rect 37971 15456 38016 15484
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 11324 15419 11382 15425
rect 11324 15385 11336 15419
rect 11370 15416 11382 15419
rect 12066 15416 12072 15428
rect 11370 15388 12072 15416
rect 11370 15385 11382 15388
rect 11324 15379 11382 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 26044 15419 26102 15425
rect 26044 15385 26056 15419
rect 26090 15416 26102 15419
rect 26234 15416 26240 15428
rect 26090 15388 26240 15416
rect 26090 15385 26102 15388
rect 26044 15379 26102 15385
rect 26234 15376 26240 15388
rect 26292 15376 26298 15428
rect 36630 15376 36636 15428
rect 36688 15416 36694 15428
rect 37001 15419 37059 15425
rect 37001 15416 37013 15419
rect 36688 15388 37013 15416
rect 36688 15376 36694 15388
rect 37001 15385 37013 15388
rect 37047 15385 37059 15419
rect 37001 15379 37059 15385
rect 3786 15348 3792 15360
rect 3747 15320 3792 15348
rect 3786 15308 3792 15320
rect 3844 15308 3850 15360
rect 31478 15348 31484 15360
rect 31439 15320 31484 15348
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 7285 15147 7343 15153
rect 7285 15113 7297 15147
rect 7331 15144 7343 15147
rect 7558 15144 7564 15156
rect 7331 15116 7564 15144
rect 7331 15113 7343 15116
rect 7285 15107 7343 15113
rect 7558 15104 7564 15116
rect 7616 15104 7622 15156
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 11514 15144 11520 15156
rect 10652 15116 11520 15144
rect 10652 15104 10658 15116
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 17126 15144 17132 15156
rect 17087 15116 17132 15144
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 22922 15104 22928 15156
rect 22980 15144 22986 15156
rect 23201 15147 23259 15153
rect 23201 15144 23213 15147
rect 22980 15116 23213 15144
rect 22980 15104 22986 15116
rect 23201 15113 23213 15116
rect 23247 15113 23259 15147
rect 23201 15107 23259 15113
rect 28261 15147 28319 15153
rect 28261 15113 28273 15147
rect 28307 15144 28319 15147
rect 28994 15144 29000 15156
rect 28307 15116 29000 15144
rect 28307 15113 28319 15116
rect 28261 15107 28319 15113
rect 28994 15104 29000 15116
rect 29052 15104 29058 15156
rect 29641 15147 29699 15153
rect 29641 15113 29653 15147
rect 29687 15144 29699 15147
rect 30558 15144 30564 15156
rect 29687 15116 30564 15144
rect 29687 15113 29699 15116
rect 29641 15107 29699 15113
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 36538 15104 36544 15156
rect 36596 15144 36602 15156
rect 36633 15147 36691 15153
rect 36633 15144 36645 15147
rect 36596 15116 36645 15144
rect 36596 15104 36602 15116
rect 36633 15113 36645 15116
rect 36679 15113 36691 15147
rect 36633 15107 36691 15113
rect 37366 15104 37372 15156
rect 37424 15144 37430 15156
rect 37461 15147 37519 15153
rect 37461 15144 37473 15147
rect 37424 15116 37473 15144
rect 37424 15104 37430 15116
rect 37461 15113 37473 15116
rect 37507 15113 37519 15147
rect 38010 15144 38016 15156
rect 37971 15116 38016 15144
rect 37461 15107 37519 15113
rect 38010 15104 38016 15116
rect 38068 15104 38074 15156
rect 22002 15036 22008 15088
rect 22060 15076 22066 15088
rect 22373 15079 22431 15085
rect 22373 15076 22385 15079
rect 22060 15048 22385 15076
rect 22060 15036 22066 15048
rect 22373 15045 22385 15048
rect 22419 15045 22431 15079
rect 22373 15039 22431 15045
rect 28721 15079 28779 15085
rect 28721 15045 28733 15079
rect 28767 15076 28779 15079
rect 29178 15076 29184 15088
rect 28767 15048 29184 15076
rect 28767 15045 28779 15048
rect 28721 15039 28779 15045
rect 29178 15036 29184 15048
rect 29236 15036 29242 15088
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 7190 15008 7196 15020
rect 4120 14980 7196 15008
rect 4120 14968 4126 14980
rect 7190 14968 7196 14980
rect 7248 15008 7254 15020
rect 7469 15011 7527 15017
rect 7469 15008 7481 15011
rect 7248 14980 7481 15008
rect 7248 14968 7254 14980
rect 7469 14977 7481 14980
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17678 15008 17684 15020
rect 17267 14980 17684 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17678 14968 17684 14980
rect 17736 14968 17742 15020
rect 22554 15008 22560 15020
rect 22515 14980 22560 15008
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 24486 14968 24492 15020
rect 24544 15008 24550 15020
rect 35989 15011 36047 15017
rect 35989 15008 36001 15011
rect 24544 14980 36001 15008
rect 24544 14968 24550 14980
rect 35989 14977 36001 14980
rect 36035 15008 36047 15011
rect 36541 15011 36599 15017
rect 36541 15008 36553 15011
rect 36035 14980 36553 15008
rect 36035 14977 36047 14980
rect 35989 14971 36047 14977
rect 36541 14977 36553 14980
rect 36587 14977 36599 15011
rect 36541 14971 36599 14977
rect 37277 15011 37335 15017
rect 37277 14977 37289 15011
rect 37323 15008 37335 15011
rect 38470 15008 38476 15020
rect 37323 14980 38476 15008
rect 37323 14977 37335 14980
rect 37277 14971 37335 14977
rect 38470 14968 38476 14980
rect 38528 14968 38534 15020
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7742 14940 7748 14952
rect 7699 14912 7748 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 24394 14940 24400 14952
rect 11664 14912 24400 14940
rect 11664 14900 11670 14912
rect 24394 14900 24400 14912
rect 24452 14900 24458 14952
rect 24504 14912 28488 14940
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 24504 14872 24532 14912
rect 28353 14875 28411 14881
rect 28353 14872 28365 14875
rect 18012 14844 24532 14872
rect 27724 14844 28365 14872
rect 18012 14832 18018 14844
rect 14642 14804 14648 14816
rect 14603 14776 14648 14804
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 23750 14804 23756 14816
rect 23711 14776 23756 14804
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 27724 14813 27752 14844
rect 28353 14841 28365 14844
rect 28399 14841 28411 14875
rect 28460 14872 28488 14912
rect 29454 14872 29460 14884
rect 28460 14844 29460 14872
rect 28353 14835 28411 14841
rect 29454 14832 29460 14844
rect 29512 14832 29518 14884
rect 27709 14807 27767 14813
rect 27709 14804 27721 14807
rect 23992 14776 27721 14804
rect 23992 14764 23998 14776
rect 27709 14773 27721 14776
rect 27755 14773 27767 14807
rect 27709 14767 27767 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 13630 14560 13636 14612
rect 13688 14600 13694 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 13688 14572 14289 14600
rect 13688 14560 13694 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14976 14572 15117 14600
rect 14976 14560 14982 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 23934 14600 23940 14612
rect 19392 14572 23940 14600
rect 19392 14560 19398 14572
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 24394 14600 24400 14612
rect 24355 14572 24400 14600
rect 24394 14560 24400 14572
rect 24452 14560 24458 14612
rect 29454 14560 29460 14612
rect 29512 14600 29518 14612
rect 29549 14603 29607 14609
rect 29549 14600 29561 14603
rect 29512 14572 29561 14600
rect 29512 14560 29518 14572
rect 29549 14569 29561 14572
rect 29595 14569 29607 14603
rect 29549 14563 29607 14569
rect 10778 14492 10784 14544
rect 10836 14532 10842 14544
rect 23750 14532 23756 14544
rect 10836 14504 23756 14532
rect 10836 14492 10842 14504
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 15749 14467 15807 14473
rect 6880 14436 7604 14464
rect 6880 14424 6886 14436
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7576 14405 7604 14436
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 20806 14464 20812 14476
rect 15795 14436 20812 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7742 14396 7748 14408
rect 7703 14368 7748 14396
rect 7561 14359 7619 14365
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15764 14396 15792 14427
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 22922 14424 22928 14476
rect 22980 14464 22986 14476
rect 23109 14467 23167 14473
rect 23109 14464 23121 14467
rect 22980 14436 23121 14464
rect 22980 14424 22986 14436
rect 23109 14433 23121 14436
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 15059 14368 15792 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 23676 14405 23704 14504
rect 23750 14492 23756 14504
rect 23808 14492 23814 14544
rect 23845 14535 23903 14541
rect 23845 14501 23857 14535
rect 23891 14532 23903 14535
rect 24854 14532 24860 14544
rect 23891 14504 24860 14532
rect 23891 14501 23903 14504
rect 23845 14495 23903 14501
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22796 14368 22845 14396
rect 22796 14356 22802 14368
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 36817 14399 36875 14405
rect 36817 14365 36829 14399
rect 36863 14396 36875 14399
rect 37274 14396 37280 14408
rect 36863 14368 37280 14396
rect 36863 14365 36875 14368
rect 36817 14359 36875 14365
rect 37274 14356 37280 14368
rect 37332 14356 37338 14408
rect 37550 14396 37556 14408
rect 37511 14368 37556 14396
rect 37550 14356 37556 14368
rect 37608 14356 37614 14408
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 14829 14331 14887 14337
rect 14829 14328 14841 14331
rect 14700 14300 14841 14328
rect 14700 14288 14706 14300
rect 14829 14297 14841 14300
rect 14875 14297 14887 14331
rect 14829 14291 14887 14297
rect 16206 14288 16212 14340
rect 16264 14328 16270 14340
rect 25314 14328 25320 14340
rect 16264 14300 25320 14328
rect 16264 14288 16270 14300
rect 25314 14288 25320 14300
rect 25372 14288 25378 14340
rect 7101 14263 7159 14269
rect 7101 14229 7113 14263
rect 7147 14260 7159 14263
rect 7190 14260 7196 14272
rect 7147 14232 7196 14260
rect 7147 14229 7159 14232
rect 7101 14223 7159 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 31389 14059 31447 14065
rect 31389 14056 31401 14059
rect 15620 14028 22094 14056
rect 15620 14016 15626 14028
rect 4525 13991 4583 13997
rect 4525 13988 4537 13991
rect 2700 13960 4537 13988
rect 2700 13929 2728 13960
rect 4525 13957 4537 13960
rect 4571 13988 4583 13991
rect 6914 13988 6920 14000
rect 4571 13960 6920 13988
rect 4571 13957 4583 13960
rect 4525 13951 4583 13957
rect 6914 13948 6920 13960
rect 6972 13988 6978 14000
rect 9950 13988 9956 14000
rect 6972 13960 9956 13988
rect 6972 13948 6978 13960
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 14182 13988 14188 14000
rect 14143 13960 14188 13988
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 16114 13948 16120 14000
rect 16172 13988 16178 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16172 13960 17049 13988
rect 16172 13948 16178 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2952 13923 3010 13929
rect 2952 13889 2964 13923
rect 2998 13920 3010 13923
rect 3786 13920 3792 13932
rect 2998 13892 3792 13920
rect 2998 13889 3010 13892
rect 2952 13883 3010 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 14458 13920 14464 13932
rect 14047 13892 14464 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 17218 13920 17224 13932
rect 17179 13892 17224 13920
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 22066 13920 22094 14028
rect 25608 14028 31401 14056
rect 24305 13991 24363 13997
rect 24305 13957 24317 13991
rect 24351 13988 24363 13991
rect 24394 13988 24400 14000
rect 24351 13960 24400 13988
rect 24351 13957 24363 13960
rect 24305 13951 24363 13957
rect 24394 13948 24400 13960
rect 24452 13948 24458 14000
rect 24489 13991 24547 13997
rect 24489 13957 24501 13991
rect 24535 13988 24547 13991
rect 25406 13988 25412 14000
rect 24535 13960 25412 13988
rect 24535 13957 24547 13960
rect 24489 13951 24547 13957
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 23477 13923 23535 13929
rect 23477 13920 23489 13923
rect 22066 13892 23489 13920
rect 23477 13889 23489 13892
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 23658 13880 23664 13932
rect 23716 13920 23722 13932
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 23716 13892 23765 13920
rect 23716 13880 23722 13892
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 25314 13880 25320 13932
rect 25372 13920 25378 13932
rect 25501 13923 25559 13929
rect 25501 13920 25513 13923
rect 25372 13892 25513 13920
rect 25372 13880 25378 13892
rect 25501 13889 25513 13892
rect 25547 13889 25559 13923
rect 25501 13883 25559 13889
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 13446 13852 13452 13864
rect 11848 13824 13452 13852
rect 11848 13812 11854 13824
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 14642 13852 14648 13864
rect 14603 13824 14648 13852
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 17862 13852 17868 13864
rect 15151 13824 17868 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 18506 13812 18512 13864
rect 18564 13852 18570 13864
rect 25608 13852 25636 14028
rect 31389 14025 31401 14028
rect 31435 14025 31447 14059
rect 31389 14019 31447 14025
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 37734 14056 37740 14068
rect 37332 14028 37740 14056
rect 37332 14016 37338 14028
rect 37734 14016 37740 14028
rect 37792 14016 37798 14068
rect 25685 13991 25743 13997
rect 25685 13957 25697 13991
rect 25731 13988 25743 13991
rect 26237 13991 26295 13997
rect 26237 13988 26249 13991
rect 25731 13960 26249 13988
rect 25731 13957 25743 13960
rect 25685 13951 25743 13957
rect 26237 13957 26249 13960
rect 26283 13988 26295 13991
rect 26326 13988 26332 14000
rect 26283 13960 26332 13988
rect 26283 13957 26295 13960
rect 26237 13951 26295 13957
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 31478 13988 31484 14000
rect 31439 13960 31484 13988
rect 31478 13948 31484 13960
rect 31536 13948 31542 14000
rect 37921 13991 37979 13997
rect 37921 13957 37933 13991
rect 37967 13988 37979 13991
rect 38654 13988 38660 14000
rect 37967 13960 38660 13988
rect 37967 13957 37979 13960
rect 37921 13951 37979 13957
rect 38654 13948 38660 13960
rect 38712 13948 38718 14000
rect 37734 13920 37740 13932
rect 37695 13892 37740 13920
rect 37734 13880 37740 13892
rect 37792 13880 37798 13932
rect 18564 13824 25636 13852
rect 18564 13812 18570 13824
rect 13630 13744 13636 13796
rect 13688 13784 13694 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 13688 13756 14933 13784
rect 13688 13744 13694 13756
rect 14921 13753 14933 13756
rect 14967 13753 14979 13787
rect 14921 13747 14979 13753
rect 14090 13676 14096 13728
rect 14148 13716 14154 13728
rect 15746 13716 15752 13728
rect 14148 13688 15752 13716
rect 14148 13676 14154 13688
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22612 13484 22845 13512
rect 22612 13472 22618 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 23716 13484 24409 13512
rect 23716 13472 23722 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 23750 13376 23756 13388
rect 23523 13348 23756 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13308 23351 13311
rect 37550 13308 37556 13320
rect 23339 13280 37556 13308
rect 23339 13277 23351 13280
rect 23293 13271 23351 13277
rect 37550 13268 37556 13280
rect 37608 13268 37614 13320
rect 24118 13200 24124 13252
rect 24176 13240 24182 13252
rect 37461 13243 37519 13249
rect 37461 13240 37473 13243
rect 24176 13212 37473 13240
rect 24176 13200 24182 13212
rect 37461 13209 37473 13212
rect 37507 13240 37519 13243
rect 37734 13240 37740 13252
rect 37507 13212 37740 13240
rect 37507 13209 37519 13212
rect 37461 13203 37519 13209
rect 37734 13200 37740 13212
rect 37792 13200 37798 13252
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 13136 13144 14473 13172
rect 13136 13132 13142 13144
rect 14461 13141 14473 13144
rect 14507 13172 14519 13175
rect 14642 13172 14648 13184
rect 14507 13144 14648 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 22278 13172 22284 13184
rect 22239 13144 22284 13172
rect 22278 13132 22284 13144
rect 22336 13172 22342 13184
rect 23201 13175 23259 13181
rect 23201 13172 23213 13175
rect 22336 13144 23213 13172
rect 22336 13132 22342 13144
rect 23201 13141 23213 13144
rect 23247 13141 23259 13175
rect 23201 13135 23259 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7800 12940 8309 12968
rect 7800 12928 7806 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 22278 12968 22284 12980
rect 8297 12931 8355 12937
rect 17236 12940 22284 12968
rect 8757 12903 8815 12909
rect 8757 12900 8769 12903
rect 6932 12872 8769 12900
rect 6932 12844 6960 12872
rect 8757 12869 8769 12872
rect 8803 12869 8815 12903
rect 8757 12863 8815 12869
rect 13265 12903 13323 12909
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 13906 12900 13912 12912
rect 13311 12872 13912 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 6914 12832 6920 12844
rect 6875 12804 6920 12832
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7190 12841 7196 12844
rect 7184 12832 7196 12841
rect 7151 12804 7196 12832
rect 7184 12795 7196 12804
rect 7190 12792 7196 12795
rect 7248 12792 7254 12844
rect 12158 12792 12164 12844
rect 12216 12832 12222 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12216 12804 13093 12832
rect 12216 12792 12222 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 17236 12764 17264 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 25774 12968 25780 12980
rect 25735 12940 25780 12968
rect 25774 12928 25780 12940
rect 25832 12928 25838 12980
rect 17862 12860 17868 12912
rect 17920 12900 17926 12912
rect 17920 12872 33456 12900
rect 17920 12860 17926 12872
rect 25961 12835 26019 12841
rect 25961 12801 25973 12835
rect 26007 12832 26019 12835
rect 28902 12832 28908 12844
rect 26007 12804 28908 12832
rect 26007 12801 26019 12804
rect 25961 12795 26019 12801
rect 28902 12792 28908 12804
rect 28960 12792 28966 12844
rect 33428 12841 33456 12872
rect 32125 12835 32183 12841
rect 32125 12801 32137 12835
rect 32171 12832 32183 12835
rect 33413 12835 33471 12841
rect 32171 12804 32812 12832
rect 32171 12801 32183 12804
rect 32125 12795 32183 12801
rect 32398 12764 32404 12776
rect 10744 12736 17264 12764
rect 32359 12736 32404 12764
rect 10744 12724 10750 12736
rect 32398 12724 32404 12736
rect 32456 12724 32462 12776
rect 32784 12764 32812 12804
rect 33413 12801 33425 12835
rect 33459 12832 33471 12835
rect 34057 12835 34115 12841
rect 34057 12832 34069 12835
rect 33459 12804 34069 12832
rect 33459 12801 33471 12804
rect 33413 12795 33471 12801
rect 34057 12801 34069 12804
rect 34103 12801 34115 12835
rect 34057 12795 34115 12801
rect 33778 12764 33784 12776
rect 32784 12736 33784 12764
rect 33778 12724 33784 12736
rect 33836 12724 33842 12776
rect 19794 12628 19800 12640
rect 19755 12600 19800 12628
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 23750 12628 23756 12640
rect 23711 12600 23756 12628
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 33597 12631 33655 12637
rect 33597 12597 33609 12631
rect 33643 12628 33655 12631
rect 33870 12628 33876 12640
rect 33643 12600 33876 12628
rect 33643 12597 33655 12600
rect 33597 12591 33655 12597
rect 33870 12588 33876 12600
rect 33928 12588 33934 12640
rect 38102 12628 38108 12640
rect 38063 12600 38108 12628
rect 38102 12588 38108 12600
rect 38160 12588 38166 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 10226 12424 10232 12436
rect 10187 12396 10232 12424
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 20714 12424 20720 12436
rect 19567 12396 20720 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 31018 12384 31024 12436
rect 31076 12424 31082 12436
rect 31113 12427 31171 12433
rect 31113 12424 31125 12427
rect 31076 12396 31125 12424
rect 31076 12384 31082 12396
rect 31113 12393 31125 12396
rect 31159 12393 31171 12427
rect 31113 12387 31171 12393
rect 4433 12359 4491 12365
rect 4433 12325 4445 12359
rect 4479 12356 4491 12359
rect 4706 12356 4712 12368
rect 4479 12328 4712 12356
rect 4479 12325 4491 12328
rect 4433 12319 4491 12325
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 20625 12359 20683 12365
rect 20625 12325 20637 12359
rect 20671 12356 20683 12359
rect 21818 12356 21824 12368
rect 20671 12328 21824 12356
rect 20671 12325 20683 12328
rect 20625 12319 20683 12325
rect 21818 12316 21824 12328
rect 21876 12356 21882 12368
rect 21913 12359 21971 12365
rect 21913 12356 21925 12359
rect 21876 12328 21925 12356
rect 21876 12316 21882 12328
rect 21913 12325 21925 12328
rect 21959 12325 21971 12359
rect 21913 12319 21971 12325
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 10226 12220 10232 12232
rect 9539 12192 10232 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 4249 12155 4307 12161
rect 4249 12121 4261 12155
rect 4295 12152 4307 12155
rect 4614 12152 4620 12164
rect 4295 12124 4620 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 18601 12155 18659 12161
rect 18601 12152 18613 12155
rect 10376 12124 18613 12152
rect 10376 12112 10382 12124
rect 18601 12121 18613 12124
rect 18647 12152 18659 12155
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 18647 12124 19257 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 19426 12112 19432 12164
rect 19484 12152 19490 12164
rect 19794 12152 19800 12164
rect 19484 12124 19800 12152
rect 19484 12112 19490 12124
rect 19794 12112 19800 12124
rect 19852 12152 19858 12164
rect 20901 12155 20959 12161
rect 20901 12152 20913 12155
rect 19852 12124 20913 12152
rect 19852 12112 19858 12124
rect 20901 12121 20913 12124
rect 20947 12121 20959 12155
rect 23750 12152 23756 12164
rect 20901 12115 20959 12121
rect 22066 12124 23756 12152
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 11330 12084 11336 12096
rect 9723 12056 11336 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 20438 12084 20444 12096
rect 20399 12056 20444 12084
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20916 12084 20944 12115
rect 21453 12087 21511 12093
rect 21453 12084 21465 12087
rect 20916 12056 21465 12084
rect 21453 12053 21465 12056
rect 21499 12084 21511 12087
rect 22066 12084 22094 12124
rect 23750 12112 23756 12124
rect 23808 12152 23814 12164
rect 23808 12124 28488 12152
rect 23808 12112 23814 12124
rect 27982 12084 27988 12096
rect 21499 12056 22094 12084
rect 27895 12056 27988 12084
rect 21499 12053 21511 12056
rect 21453 12047 21511 12053
rect 27982 12044 27988 12056
rect 28040 12084 28046 12096
rect 28350 12084 28356 12096
rect 28040 12056 28356 12084
rect 28040 12044 28046 12056
rect 28350 12044 28356 12056
rect 28408 12044 28414 12096
rect 28460 12084 28488 12124
rect 31110 12112 31116 12164
rect 31168 12152 31174 12164
rect 31389 12155 31447 12161
rect 31389 12152 31401 12155
rect 31168 12124 31401 12152
rect 31168 12112 31174 12124
rect 31389 12121 31401 12124
rect 31435 12121 31447 12155
rect 31389 12115 31447 12121
rect 37918 12084 37924 12096
rect 28460 12056 37924 12084
rect 37918 12044 37924 12056
rect 37976 12044 37982 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2832 11852 2881 11880
rect 2832 11840 2838 11852
rect 2869 11849 2881 11852
rect 2915 11849 2927 11883
rect 2869 11843 2927 11849
rect 10321 11883 10379 11889
rect 10321 11849 10333 11883
rect 10367 11880 10379 11883
rect 12434 11880 12440 11892
rect 10367 11852 12440 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 16632 11852 17693 11880
rect 16632 11840 16638 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 17681 11843 17739 11849
rect 19061 11883 19119 11889
rect 19061 11849 19073 11883
rect 19107 11880 19119 11883
rect 20070 11880 20076 11892
rect 19107 11852 20076 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 28902 11840 28908 11892
rect 28960 11880 28966 11892
rect 30193 11883 30251 11889
rect 30193 11880 30205 11883
rect 28960 11852 30205 11880
rect 28960 11840 28966 11852
rect 30193 11849 30205 11852
rect 30239 11849 30251 11883
rect 31110 11880 31116 11892
rect 31071 11852 31116 11880
rect 30193 11843 30251 11849
rect 31110 11840 31116 11852
rect 31168 11840 31174 11892
rect 3697 11815 3755 11821
rect 3697 11781 3709 11815
rect 3743 11812 3755 11815
rect 4798 11812 4804 11824
rect 3743 11784 4804 11812
rect 3743 11781 3755 11784
rect 3697 11775 3755 11781
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 18141 11815 18199 11821
rect 18141 11781 18153 11815
rect 18187 11812 18199 11815
rect 18601 11815 18659 11821
rect 18601 11812 18613 11815
rect 18187 11784 18613 11812
rect 18187 11781 18199 11784
rect 18141 11775 18199 11781
rect 18601 11781 18613 11784
rect 18647 11812 18659 11815
rect 19426 11812 19432 11824
rect 18647 11784 19432 11812
rect 18647 11781 18659 11784
rect 18601 11775 18659 11781
rect 19426 11772 19432 11784
rect 19484 11812 19490 11824
rect 19521 11815 19579 11821
rect 19521 11812 19533 11815
rect 19484 11784 19533 11812
rect 19484 11772 19490 11784
rect 19521 11781 19533 11784
rect 19567 11781 19579 11815
rect 22462 11812 22468 11824
rect 22423 11784 22468 11812
rect 19521 11775 19579 11781
rect 22462 11772 22468 11784
rect 22520 11772 22526 11824
rect 27617 11815 27675 11821
rect 27617 11781 27629 11815
rect 27663 11812 27675 11815
rect 27982 11812 27988 11824
rect 27663 11784 27988 11812
rect 27663 11781 27675 11784
rect 27617 11775 27675 11781
rect 27982 11772 27988 11784
rect 28040 11812 28046 11824
rect 28077 11815 28135 11821
rect 28077 11812 28089 11815
rect 28040 11784 28089 11812
rect 28040 11772 28046 11784
rect 28077 11781 28089 11784
rect 28123 11812 28135 11815
rect 30653 11815 30711 11821
rect 30653 11812 30665 11815
rect 28123 11784 30665 11812
rect 28123 11781 28135 11784
rect 28077 11775 28135 11781
rect 30653 11781 30665 11784
rect 30699 11812 30711 11815
rect 31573 11815 31631 11821
rect 31573 11812 31585 11815
rect 30699 11784 31585 11812
rect 30699 11781 30711 11784
rect 30653 11775 30711 11781
rect 31573 11781 31585 11784
rect 31619 11812 31631 11815
rect 32398 11812 32404 11824
rect 31619 11784 32404 11812
rect 31619 11781 31631 11784
rect 31573 11775 31631 11781
rect 32398 11772 32404 11784
rect 32456 11772 32462 11824
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2464 11716 2789 11744
rect 2464 11704 2470 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 3510 11744 3516 11756
rect 3471 11716 3516 11744
rect 2777 11707 2835 11713
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11744 10195 11747
rect 20438 11744 20444 11756
rect 10183 11716 20444 11744
rect 10183 11713 10195 11716
rect 10137 11707 10195 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22281 11747 22339 11753
rect 22281 11744 22293 11747
rect 22060 11716 22293 11744
rect 22060 11704 22066 11716
rect 22281 11713 22293 11716
rect 22327 11713 22339 11747
rect 22281 11707 22339 11713
rect 11974 11636 11980 11688
rect 12032 11676 12038 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 12032 11648 12081 11676
rect 12032 11636 12038 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 24578 11676 24584 11688
rect 12069 11639 12127 11645
rect 12176 11648 17908 11676
rect 10870 11568 10876 11620
rect 10928 11608 10934 11620
rect 12176 11608 12204 11648
rect 10928 11580 12204 11608
rect 12437 11611 12495 11617
rect 10928 11568 10934 11580
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 12483 11580 13124 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 12526 11540 12532 11552
rect 12487 11512 12532 11540
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13096 11549 13124 11580
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 17773 11611 17831 11617
rect 17773 11608 17785 11611
rect 15068 11580 17785 11608
rect 15068 11568 15074 11580
rect 17773 11577 17785 11580
rect 17819 11577 17831 11611
rect 17880 11608 17908 11648
rect 18984 11648 24584 11676
rect 18877 11611 18935 11617
rect 18877 11608 18889 11611
rect 17880 11580 18889 11608
rect 17773 11571 17831 11577
rect 18877 11577 18889 11580
rect 18923 11577 18935 11611
rect 18877 11571 18935 11577
rect 13081 11543 13139 11549
rect 13081 11509 13093 11543
rect 13127 11540 13139 11543
rect 18984 11540 19012 11648
rect 24578 11636 24584 11648
rect 24636 11636 24642 11688
rect 31036 11648 31340 11676
rect 26786 11568 26792 11620
rect 26844 11608 26850 11620
rect 27249 11611 27307 11617
rect 27249 11608 27261 11611
rect 26844 11580 27261 11608
rect 26844 11568 26850 11580
rect 27249 11577 27261 11580
rect 27295 11577 27307 11611
rect 28350 11608 28356 11620
rect 28311 11580 28356 11608
rect 27249 11571 27307 11577
rect 28350 11568 28356 11580
rect 28408 11568 28414 11620
rect 30377 11611 30435 11617
rect 30377 11577 30389 11611
rect 30423 11608 30435 11611
rect 31036 11608 31064 11648
rect 31202 11608 31208 11620
rect 30423 11580 31064 11608
rect 31163 11580 31208 11608
rect 30423 11577 30435 11580
rect 30377 11571 30435 11577
rect 31202 11568 31208 11580
rect 31260 11568 31266 11620
rect 27154 11540 27160 11552
rect 13127 11512 19012 11540
rect 27115 11512 27160 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 27154 11500 27160 11512
rect 27212 11500 27218 11552
rect 28534 11540 28540 11552
rect 28495 11512 28540 11540
rect 28534 11500 28540 11512
rect 28592 11500 28598 11552
rect 31312 11540 31340 11648
rect 32030 11540 32036 11552
rect 31312 11512 32036 11540
rect 32030 11500 32036 11512
rect 32088 11500 32094 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 12713 11339 12771 11345
rect 12713 11305 12725 11339
rect 12759 11336 12771 11339
rect 13722 11336 13728 11348
rect 12759 11308 13728 11336
rect 12759 11305 12771 11308
rect 12713 11299 12771 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 18325 11339 18383 11345
rect 18325 11305 18337 11339
rect 18371 11336 18383 11339
rect 19426 11336 19432 11348
rect 18371 11308 19432 11336
rect 18371 11305 18383 11308
rect 18325 11299 18383 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 26786 11296 26792 11348
rect 26844 11336 26850 11348
rect 26973 11339 27031 11345
rect 26973 11336 26985 11339
rect 26844 11308 26985 11336
rect 26844 11296 26850 11308
rect 26973 11305 26985 11308
rect 27019 11305 27031 11339
rect 37918 11336 37924 11348
rect 37879 11308 37924 11336
rect 26973 11299 27031 11305
rect 37918 11296 37924 11308
rect 37976 11296 37982 11348
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 15010 11268 15016 11280
rect 8812 11240 15016 11268
rect 8812 11228 8818 11240
rect 15010 11228 15016 11240
rect 15068 11228 15074 11280
rect 27798 11228 27804 11280
rect 27856 11268 27862 11280
rect 28261 11271 28319 11277
rect 28261 11268 28273 11271
rect 27856 11240 28273 11268
rect 27856 11228 27862 11240
rect 28261 11237 28273 11240
rect 28307 11237 28319 11271
rect 28261 11231 28319 11237
rect 33321 11271 33379 11277
rect 33321 11237 33333 11271
rect 33367 11268 33379 11271
rect 33594 11268 33600 11280
rect 33367 11240 33600 11268
rect 33367 11237 33379 11240
rect 33321 11231 33379 11237
rect 33594 11228 33600 11240
rect 33652 11228 33658 11280
rect 27982 11200 27988 11212
rect 27943 11172 27988 11200
rect 27982 11160 27988 11172
rect 28040 11160 28046 11212
rect 28442 11200 28448 11212
rect 28403 11172 28448 11200
rect 28442 11160 28448 11172
rect 28500 11160 28506 11212
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2096 11104 2697 11132
rect 2096 11092 2102 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11974 11132 11980 11144
rect 11204 11104 11980 11132
rect 11204 11092 11210 11104
rect 11974 11092 11980 11104
rect 12032 11132 12038 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12032 11104 12817 11132
rect 12032 11092 12038 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 37369 11135 37427 11141
rect 37369 11101 37381 11135
rect 37415 11132 37427 11135
rect 38102 11132 38108 11144
rect 37415 11104 38108 11132
rect 37415 11101 37427 11104
rect 37369 11095 37427 11101
rect 38102 11092 38108 11104
rect 38160 11092 38166 11144
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 10410 11064 10416 11076
rect 2915 11036 10416 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13538 11064 13544 11076
rect 13035 11036 13544 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 20990 11024 20996 11076
rect 21048 11064 21054 11076
rect 22002 11064 22008 11076
rect 21048 11036 22008 11064
rect 21048 11024 21054 11036
rect 22002 11024 22008 11036
rect 22060 11064 22066 11076
rect 22097 11067 22155 11073
rect 22097 11064 22109 11067
rect 22060 11036 22109 11064
rect 22060 11024 22066 11036
rect 22097 11033 22109 11036
rect 22143 11033 22155 11067
rect 22097 11027 22155 11033
rect 26878 11024 26884 11076
rect 26936 11064 26942 11076
rect 33137 11067 33195 11073
rect 33137 11064 33149 11067
rect 26936 11036 33149 11064
rect 26936 11024 26942 11036
rect 33137 11033 33149 11036
rect 33183 11033 33195 11067
rect 33137 11027 33195 11033
rect 35342 11024 35348 11076
rect 35400 11064 35406 11076
rect 37274 11064 37280 11076
rect 35400 11036 37280 11064
rect 35400 11024 35406 11036
rect 37274 11024 37280 11036
rect 37332 11024 37338 11076
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 27798 10792 27804 10804
rect 27759 10764 27804 10792
rect 27798 10752 27804 10764
rect 27856 10752 27862 10804
rect 35986 10792 35992 10804
rect 35947 10764 35992 10792
rect 35986 10752 35992 10764
rect 36044 10752 36050 10804
rect 37366 10752 37372 10804
rect 37424 10792 37430 10804
rect 37461 10795 37519 10801
rect 37461 10792 37473 10795
rect 37424 10764 37473 10792
rect 37424 10752 37430 10764
rect 37461 10761 37473 10764
rect 37507 10761 37519 10795
rect 37461 10755 37519 10761
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 5534 10724 5540 10736
rect 5123 10696 5540 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12526 10656 12532 10668
rect 12207 10628 12532 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 36004 10656 36032 10752
rect 36541 10659 36599 10665
rect 36541 10656 36553 10659
rect 36004 10628 36553 10656
rect 36541 10625 36553 10628
rect 36587 10625 36599 10659
rect 37274 10656 37280 10668
rect 37235 10628 37280 10656
rect 36541 10619 36599 10625
rect 37274 10616 37280 10628
rect 37332 10616 37338 10668
rect 12345 10455 12403 10461
rect 12345 10421 12357 10455
rect 12391 10452 12403 10455
rect 12986 10452 12992 10464
rect 12391 10424 12992 10452
rect 12391 10421 12403 10424
rect 12345 10415 12403 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 36722 10452 36728 10464
rect 36683 10424 36728 10452
rect 36722 10412 36728 10424
rect 36780 10412 36786 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2866 10248 2872 10260
rect 2827 10220 2872 10248
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 15286 10248 15292 10260
rect 14844 10220 15292 10248
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 7098 10180 7104 10192
rect 6227 10152 7104 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 14844 10189 14872 10220
rect 15286 10208 15292 10220
rect 15344 10248 15350 10260
rect 15381 10251 15439 10257
rect 15381 10248 15393 10251
rect 15344 10220 15393 10248
rect 15344 10208 15350 10220
rect 15381 10217 15393 10220
rect 15427 10217 15439 10251
rect 15381 10211 15439 10217
rect 17681 10251 17739 10257
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 17770 10248 17776 10260
rect 17727 10220 17776 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 14829 10183 14887 10189
rect 14829 10149 14841 10183
rect 14875 10149 14887 10183
rect 14829 10143 14887 10149
rect 17037 10183 17095 10189
rect 17037 10149 17049 10183
rect 17083 10180 17095 10183
rect 17402 10180 17408 10192
rect 17083 10152 17408 10180
rect 17083 10149 17095 10152
rect 17037 10143 17095 10149
rect 17402 10140 17408 10152
rect 17460 10140 17466 10192
rect 27154 10004 27160 10056
rect 27212 10044 27218 10056
rect 28445 10047 28503 10053
rect 28445 10044 28457 10047
rect 27212 10016 28457 10044
rect 27212 10004 27218 10016
rect 28445 10013 28457 10016
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 5994 9976 6000 9988
rect 2832 9948 2877 9976
rect 5955 9948 6000 9976
rect 2832 9936 2838 9948
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 14274 9936 14280 9988
rect 14332 9976 14338 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 14332 9948 14473 9976
rect 14332 9936 14338 9948
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 14461 9939 14519 9945
rect 16209 9979 16267 9985
rect 16209 9945 16221 9979
rect 16255 9976 16267 9979
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 16255 9948 16681 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 16669 9945 16681 9948
rect 16715 9976 16727 9979
rect 17034 9976 17040 9988
rect 16715 9948 17040 9976
rect 16715 9945 16727 9948
rect 16669 9939 16727 9945
rect 17034 9936 17040 9948
rect 17092 9976 17098 9988
rect 17494 9976 17500 9988
rect 17092 9948 17500 9976
rect 17092 9936 17098 9948
rect 17494 9936 17500 9948
rect 17552 9976 17558 9988
rect 17773 9979 17831 9985
rect 17773 9976 17785 9979
rect 17552 9948 17785 9976
rect 17552 9936 17558 9948
rect 17773 9945 17785 9948
rect 17819 9945 17831 9979
rect 17773 9939 17831 9945
rect 17957 9979 18015 9985
rect 17957 9945 17969 9979
rect 18003 9976 18015 9979
rect 18509 9979 18567 9985
rect 18509 9976 18521 9979
rect 18003 9948 18521 9976
rect 18003 9945 18015 9948
rect 17957 9939 18015 9945
rect 18509 9945 18521 9948
rect 18555 9976 18567 9979
rect 36998 9976 37004 9988
rect 18555 9948 37004 9976
rect 18555 9945 18567 9948
rect 18509 9939 18567 9945
rect 36998 9936 37004 9948
rect 37056 9936 37062 9988
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 13872 9880 14933 9908
rect 13872 9868 13878 9880
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 17126 9908 17132 9920
rect 17087 9880 17132 9908
rect 14921 9871 14979 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 28629 9911 28687 9917
rect 28629 9877 28641 9911
rect 28675 9908 28687 9911
rect 30742 9908 30748 9920
rect 28675 9880 30748 9908
rect 28675 9877 28687 9880
rect 28629 9871 28687 9877
rect 30742 9868 30748 9880
rect 30800 9868 30806 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 33042 9704 33048 9716
rect 17184 9676 33048 9704
rect 17184 9664 17190 9676
rect 33042 9664 33048 9676
rect 33100 9664 33106 9716
rect 9766 9636 9772 9648
rect 9727 9608 9772 9636
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 14090 9636 14096 9648
rect 14051 9608 14096 9636
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14274 9636 14280 9648
rect 14235 9608 14280 9636
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 17313 9639 17371 9645
rect 17313 9605 17325 9639
rect 17359 9636 17371 9639
rect 17402 9636 17408 9648
rect 17359 9608 17408 9636
rect 17359 9605 17371 9608
rect 17313 9599 17371 9605
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 24210 9596 24216 9648
rect 24268 9636 24274 9648
rect 24397 9639 24455 9645
rect 24397 9636 24409 9639
rect 24268 9608 24409 9636
rect 24268 9596 24274 9608
rect 24397 9605 24409 9608
rect 24443 9605 24455 9639
rect 24397 9599 24455 9605
rect 28442 9596 28448 9648
rect 28500 9636 28506 9648
rect 28500 9608 30052 9636
rect 28500 9596 28506 9608
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13814 9568 13820 9580
rect 13495 9540 13820 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 14461 9571 14519 9577
rect 14461 9568 14473 9571
rect 14424 9540 14473 9568
rect 14424 9528 14430 9540
rect 14461 9537 14473 9540
rect 14507 9537 14519 9571
rect 24765 9571 24823 9577
rect 14461 9531 14519 9537
rect 22066 9540 24716 9568
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 22066 9432 22094 9540
rect 24305 9503 24363 9509
rect 24305 9469 24317 9503
rect 24351 9469 24363 9503
rect 24688 9500 24716 9540
rect 24765 9537 24777 9571
rect 24811 9568 24823 9571
rect 25130 9568 25136 9580
rect 24811 9540 25136 9568
rect 24811 9537 24823 9540
rect 24765 9531 24823 9537
rect 25130 9528 25136 9540
rect 25188 9528 25194 9580
rect 28534 9528 28540 9580
rect 28592 9568 28598 9580
rect 30024 9577 30052 9608
rect 28997 9571 29055 9577
rect 28997 9568 29009 9571
rect 28592 9540 29009 9568
rect 28592 9528 28598 9540
rect 28997 9537 29009 9540
rect 29043 9537 29055 9571
rect 28997 9531 29055 9537
rect 30009 9571 30067 9577
rect 30009 9537 30021 9571
rect 30055 9537 30067 9571
rect 37734 9568 37740 9580
rect 37695 9540 37740 9568
rect 30009 9531 30067 9537
rect 37734 9528 37740 9540
rect 37792 9528 37798 9580
rect 27982 9500 27988 9512
rect 24688 9472 27988 9500
rect 24305 9463 24363 9469
rect 7340 9404 22094 9432
rect 7340 9392 7346 9404
rect 13633 9367 13691 9373
rect 13633 9333 13645 9367
rect 13679 9364 13691 9367
rect 13722 9364 13728 9376
rect 13679 9336 13728 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 24320 9364 24348 9463
rect 27982 9460 27988 9472
rect 28040 9460 28046 9512
rect 29181 9435 29239 9441
rect 29181 9401 29193 9435
rect 29227 9432 29239 9435
rect 31018 9432 31024 9444
rect 29227 9404 31024 9432
rect 29227 9401 29239 9404
rect 29181 9395 29239 9401
rect 31018 9392 31024 9404
rect 31076 9392 31082 9444
rect 24854 9364 24860 9376
rect 24320 9336 24860 9364
rect 24854 9324 24860 9336
rect 24912 9364 24918 9376
rect 25317 9367 25375 9373
rect 25317 9364 25329 9367
rect 24912 9336 25329 9364
rect 24912 9324 24918 9336
rect 25317 9333 25329 9336
rect 25363 9333 25375 9367
rect 25317 9327 25375 9333
rect 30193 9367 30251 9373
rect 30193 9333 30205 9367
rect 30239 9364 30251 9367
rect 31938 9364 31944 9376
rect 30239 9336 31944 9364
rect 30239 9333 30251 9336
rect 30193 9327 30251 9333
rect 31938 9324 31944 9336
rect 31996 9324 32002 9376
rect 37458 9324 37464 9376
rect 37516 9364 37522 9376
rect 37829 9367 37887 9373
rect 37829 9364 37841 9367
rect 37516 9336 37841 9364
rect 37516 9324 37522 9336
rect 37829 9333 37841 9336
rect 37875 9333 37887 9367
rect 37829 9327 37887 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3694 9160 3700 9172
rect 2884 9132 3700 9160
rect 2884 9101 2912 9132
rect 3694 9120 3700 9132
rect 3752 9160 3758 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 3752 9132 3801 9160
rect 3752 9120 3758 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 3789 9123 3847 9129
rect 4985 9163 5043 9169
rect 4985 9129 4997 9163
rect 5031 9160 5043 9163
rect 5350 9160 5356 9172
rect 5031 9132 5356 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 5350 9120 5356 9132
rect 5408 9160 5414 9172
rect 5905 9163 5963 9169
rect 5408 9132 5764 9160
rect 5408 9120 5414 9132
rect 5736 9101 5764 9132
rect 5905 9129 5917 9163
rect 5951 9160 5963 9163
rect 26142 9160 26148 9172
rect 5951 9132 26148 9160
rect 5951 9129 5963 9132
rect 5905 9123 5963 9129
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 34514 9120 34520 9172
rect 34572 9160 34578 9172
rect 34793 9163 34851 9169
rect 34793 9160 34805 9163
rect 34572 9132 34805 9160
rect 34572 9120 34578 9132
rect 34793 9129 34805 9132
rect 34839 9129 34851 9163
rect 34793 9123 34851 9129
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9061 2927 9095
rect 2869 9055 2927 9061
rect 5721 9095 5779 9101
rect 5721 9061 5733 9095
rect 5767 9061 5779 9095
rect 5721 9055 5779 9061
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 9766 9092 9772 9104
rect 9631 9064 9772 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 10505 9095 10563 9101
rect 10505 9061 10517 9095
rect 10551 9092 10563 9095
rect 10594 9092 10600 9104
rect 10551 9064 10600 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 20993 9095 21051 9101
rect 20993 9061 21005 9095
rect 21039 9092 21051 9095
rect 21542 9092 21548 9104
rect 21039 9064 21548 9092
rect 21039 9061 21051 9064
rect 20993 9055 21051 9061
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 25038 9024 25044 9036
rect 9232 8996 10364 9024
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 2866 8888 2872 8900
rect 2547 8860 2872 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 5224 8860 5457 8888
rect 5224 8848 5230 8860
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 5445 8851 5503 8857
rect 9122 8848 9128 8900
rect 9180 8888 9186 8900
rect 9232 8897 9260 8996
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 9180 8860 9229 8888
rect 9180 8848 9186 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 9217 8851 9275 8857
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 10336 8897 10364 8996
rect 22066 8996 25044 9024
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 22066 8956 22094 8996
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 25590 9024 25596 9036
rect 25551 8996 25596 9024
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 10468 8928 22094 8956
rect 10468 8916 10474 8928
rect 24026 8916 24032 8968
rect 24084 8956 24090 8968
rect 24489 8959 24547 8965
rect 24489 8956 24501 8959
rect 24084 8928 24501 8956
rect 24084 8916 24090 8928
rect 24489 8925 24501 8928
rect 24535 8925 24547 8959
rect 24489 8919 24547 8925
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 9640 8860 10149 8888
rect 9640 8848 9646 8860
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8857 10379 8891
rect 10321 8851 10379 8857
rect 20073 8891 20131 8897
rect 20073 8857 20085 8891
rect 20119 8888 20131 8891
rect 20622 8888 20628 8900
rect 20119 8860 20628 8888
rect 20119 8857 20131 8860
rect 20073 8851 20131 8857
rect 20622 8848 20628 8860
rect 20680 8848 20686 8900
rect 24854 8848 24860 8900
rect 24912 8888 24918 8900
rect 24949 8891 25007 8897
rect 24949 8888 24961 8891
rect 24912 8860 24961 8888
rect 24912 8848 24918 8860
rect 24949 8857 24961 8860
rect 24995 8888 25007 8891
rect 25884 8888 25912 8919
rect 33042 8916 33048 8968
rect 33100 8956 33106 8968
rect 35897 8959 35955 8965
rect 35897 8956 35909 8959
rect 33100 8928 35909 8956
rect 33100 8916 33106 8928
rect 35897 8925 35909 8928
rect 35943 8956 35955 8959
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 35943 8928 36553 8956
rect 35943 8925 35955 8928
rect 35897 8919 35955 8925
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 36541 8919 36599 8925
rect 37461 8959 37519 8965
rect 37461 8925 37473 8959
rect 37507 8956 37519 8959
rect 38102 8956 38108 8968
rect 37507 8928 38108 8956
rect 37507 8925 37519 8928
rect 37461 8919 37519 8925
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 24995 8860 25912 8888
rect 24995 8857 25007 8860
rect 24949 8851 25007 8857
rect 2958 8820 2964 8832
rect 2919 8792 2964 8820
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9766 8820 9772 8832
rect 9723 8792 9772 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 21085 8823 21143 8829
rect 21085 8820 21097 8823
rect 20220 8792 21097 8820
rect 20220 8780 20226 8792
rect 21085 8789 21097 8792
rect 21131 8789 21143 8823
rect 24670 8820 24676 8832
rect 24631 8792 24676 8820
rect 21085 8783 21143 8789
rect 24670 8780 24676 8792
rect 24728 8780 24734 8832
rect 25884 8820 25912 8860
rect 26053 8891 26111 8897
rect 26053 8857 26065 8891
rect 26099 8888 26111 8891
rect 26970 8888 26976 8900
rect 26099 8860 26976 8888
rect 26099 8857 26111 8860
rect 26053 8851 26111 8857
rect 26970 8848 26976 8860
rect 27028 8848 27034 8900
rect 34790 8848 34796 8900
rect 34848 8888 34854 8900
rect 35069 8891 35127 8897
rect 35069 8888 35081 8891
rect 34848 8860 35081 8888
rect 34848 8848 34854 8860
rect 35069 8857 35081 8860
rect 35115 8857 35127 8891
rect 35069 8851 35127 8857
rect 35345 8891 35403 8897
rect 35345 8857 35357 8891
rect 35391 8888 35403 8891
rect 35802 8888 35808 8900
rect 35391 8860 35808 8888
rect 35391 8857 35403 8860
rect 35345 8851 35403 8857
rect 35802 8848 35808 8860
rect 35860 8848 35866 8900
rect 36004 8860 37964 8888
rect 26605 8823 26663 8829
rect 26605 8820 26617 8823
rect 25884 8792 26617 8820
rect 26605 8789 26617 8792
rect 26651 8820 26663 8823
rect 27430 8820 27436 8832
rect 26651 8792 27436 8820
rect 26651 8789 26663 8792
rect 26605 8783 26663 8789
rect 27430 8780 27436 8792
rect 27488 8780 27494 8832
rect 35253 8823 35311 8829
rect 35253 8789 35265 8823
rect 35299 8820 35311 8823
rect 36004 8820 36032 8860
rect 35299 8792 36032 8820
rect 36081 8823 36139 8829
rect 35299 8789 35311 8792
rect 35253 8783 35311 8789
rect 36081 8789 36093 8823
rect 36127 8820 36139 8823
rect 36446 8820 36452 8832
rect 36127 8792 36452 8820
rect 36127 8789 36139 8792
rect 36081 8783 36139 8789
rect 36446 8780 36452 8792
rect 36504 8780 36510 8832
rect 37936 8829 37964 8860
rect 37921 8823 37979 8829
rect 37921 8789 37933 8823
rect 37967 8789 37979 8823
rect 37921 8783 37979 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8616 2743 8619
rect 2774 8616 2780 8628
rect 2731 8588 2780 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 23477 8619 23535 8625
rect 4203 8588 20852 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 2958 8508 2964 8560
rect 3016 8548 3022 8560
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 3016 8520 4077 8548
rect 3016 8508 3022 8520
rect 4065 8517 4077 8520
rect 4111 8517 4123 8551
rect 4065 8511 4123 8517
rect 6365 8551 6423 8557
rect 6365 8517 6377 8551
rect 6411 8548 6423 8551
rect 6454 8548 6460 8560
rect 6411 8520 6460 8548
rect 6411 8517 6423 8520
rect 6365 8511 6423 8517
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 7282 8548 7288 8560
rect 6779 8520 7288 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 12529 8551 12587 8557
rect 12529 8548 12541 8551
rect 12406 8520 12541 8548
rect 2866 8480 2872 8492
rect 2779 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5224 8452 6561 8480
rect 5224 8440 5230 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 6549 8443 6607 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 2884 8412 2912 8440
rect 2958 8412 2964 8424
rect 2884 8384 2964 8412
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11020 8384 11529 8412
rect 11020 8372 11026 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 12250 8412 12256 8424
rect 11517 8375 11575 8381
rect 11808 8384 12256 8412
rect 9953 8347 10011 8353
rect 9953 8313 9965 8347
rect 9999 8344 10011 8347
rect 11808 8344 11836 8384
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 9999 8316 11836 8344
rect 11885 8347 11943 8353
rect 9999 8313 10011 8316
rect 9953 8307 10011 8313
rect 11885 8313 11897 8347
rect 11931 8344 11943 8347
rect 12406 8344 12434 8520
rect 12529 8517 12541 8520
rect 12575 8548 12587 8551
rect 12894 8548 12900 8560
rect 12575 8520 12900 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20162 8480 20168 8492
rect 19935 8452 20168 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 18782 8372 18788 8424
rect 18840 8412 18846 8424
rect 20346 8412 20352 8424
rect 18840 8384 20352 8412
rect 18840 8372 18846 8384
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 11931 8316 12434 8344
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 17494 8304 17500 8356
rect 17552 8344 17558 8356
rect 19334 8344 19340 8356
rect 17552 8316 19340 8344
rect 17552 8304 17558 8316
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 20073 8347 20131 8353
rect 20073 8313 20085 8347
rect 20119 8344 20131 8347
rect 20254 8344 20260 8356
rect 20119 8316 20260 8344
rect 20119 8313 20131 8316
rect 20073 8307 20131 8313
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 20548 8344 20576 8443
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20717 8483 20775 8489
rect 20717 8480 20729 8483
rect 20680 8452 20729 8480
rect 20680 8440 20686 8452
rect 20717 8449 20729 8452
rect 20763 8449 20775 8483
rect 20824 8480 20852 8588
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23566 8616 23572 8628
rect 23523 8588 23572 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24854 8576 24860 8588
rect 24912 8616 24918 8628
rect 25409 8619 25467 8625
rect 25409 8616 25421 8619
rect 24912 8588 25421 8616
rect 24912 8576 24918 8588
rect 25409 8585 25421 8588
rect 25455 8585 25467 8619
rect 25409 8579 25467 8585
rect 38105 8619 38163 8625
rect 38105 8585 38117 8619
rect 38151 8616 38163 8619
rect 38286 8616 38292 8628
rect 38151 8588 38292 8616
rect 38151 8585 38163 8588
rect 38105 8579 38163 8585
rect 38286 8576 38292 8588
rect 38344 8576 38350 8628
rect 20901 8551 20959 8557
rect 20901 8517 20913 8551
rect 20947 8548 20959 8551
rect 26878 8548 26884 8560
rect 20947 8520 26884 8548
rect 20947 8517 20959 8520
rect 20901 8511 20959 8517
rect 26878 8508 26884 8520
rect 26936 8508 26942 8560
rect 32122 8508 32128 8560
rect 32180 8548 32186 8560
rect 32309 8551 32367 8557
rect 32309 8548 32321 8551
rect 32180 8520 32321 8548
rect 32180 8508 32186 8520
rect 32309 8517 32321 8520
rect 32355 8517 32367 8551
rect 32309 8511 32367 8517
rect 33229 8551 33287 8557
rect 33229 8517 33241 8551
rect 33275 8548 33287 8551
rect 33318 8548 33324 8560
rect 33275 8520 33324 8548
rect 33275 8517 33287 8520
rect 33229 8511 33287 8517
rect 33318 8508 33324 8520
rect 33376 8508 33382 8560
rect 33413 8551 33471 8557
rect 33413 8517 33425 8551
rect 33459 8548 33471 8551
rect 35802 8548 35808 8560
rect 33459 8520 35808 8548
rect 33459 8517 33471 8520
rect 33413 8511 33471 8517
rect 26694 8480 26700 8492
rect 20824 8452 26700 8480
rect 20717 8443 20775 8449
rect 26694 8440 26700 8452
rect 26752 8440 26758 8492
rect 32674 8480 32680 8492
rect 32635 8452 32680 8480
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8412 24455 8415
rect 24854 8412 24860 8424
rect 24443 8384 24860 8412
rect 24443 8381 24455 8384
rect 24397 8375 24455 8381
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 32122 8372 32128 8424
rect 32180 8412 32186 8424
rect 32217 8415 32275 8421
rect 32217 8412 32229 8415
rect 32180 8384 32229 8412
rect 32180 8372 32186 8384
rect 32217 8381 32229 8384
rect 32263 8412 32275 8415
rect 33428 8412 33456 8511
rect 35802 8508 35808 8520
rect 35860 8508 35866 8560
rect 33594 8480 33600 8492
rect 33555 8452 33600 8480
rect 33594 8440 33600 8452
rect 33652 8440 33658 8492
rect 32263 8384 33456 8412
rect 35713 8415 35771 8421
rect 32263 8381 32275 8384
rect 32217 8375 32275 8381
rect 35713 8381 35725 8415
rect 35759 8412 35771 8415
rect 37918 8412 37924 8424
rect 35759 8384 37924 8412
rect 35759 8381 35771 8384
rect 35713 8375 35771 8381
rect 37918 8372 37924 8384
rect 37976 8372 37982 8424
rect 20714 8344 20720 8356
rect 20548 8316 20720 8344
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 23566 8304 23572 8356
rect 23624 8344 23630 8356
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23624 8316 24041 8344
rect 23624 8304 23630 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 36262 8344 36268 8356
rect 36223 8316 36268 8344
rect 24029 8307 24087 8313
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 37458 8344 37464 8356
rect 37419 8316 37464 8344
rect 37458 8304 37464 8316
rect 37516 8304 37522 8356
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 11977 8279 12035 8285
rect 11977 8276 11989 8279
rect 11572 8248 11989 8276
rect 11572 8236 11578 8248
rect 11977 8245 11989 8248
rect 12023 8245 12035 8279
rect 23934 8276 23940 8288
rect 23895 8248 23940 8276
rect 11977 8239 12035 8245
rect 23934 8236 23940 8248
rect 23992 8236 23998 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 30098 8072 30104 8084
rect 30059 8044 30104 8072
rect 30098 8032 30104 8044
rect 30156 8032 30162 8084
rect 36170 8032 36176 8084
rect 36228 8072 36234 8084
rect 37185 8075 37243 8081
rect 37185 8072 37197 8075
rect 36228 8044 37197 8072
rect 36228 8032 36234 8044
rect 37185 8041 37197 8044
rect 37231 8041 37243 8075
rect 37185 8035 37243 8041
rect 11790 8004 11796 8016
rect 11751 7976 11796 8004
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 32033 7939 32091 7945
rect 32033 7905 32045 7939
rect 32079 7936 32091 7939
rect 32214 7936 32220 7948
rect 32079 7908 32220 7936
rect 32079 7905 32091 7908
rect 32033 7899 32091 7905
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10962 7868 10968 7880
rect 9916 7840 10968 7868
rect 9916 7828 9922 7840
rect 10962 7828 10968 7840
rect 11020 7868 11026 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11020 7840 11621 7868
rect 11020 7828 11026 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 23992 7840 24869 7868
rect 23992 7828 23998 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 32398 7868 32404 7880
rect 32359 7840 32404 7868
rect 24857 7831 24915 7837
rect 32398 7828 32404 7840
rect 32456 7828 32462 7880
rect 35069 7871 35127 7877
rect 35069 7837 35081 7871
rect 35115 7868 35127 7871
rect 35710 7868 35716 7880
rect 35115 7840 35716 7868
rect 35115 7837 35127 7840
rect 35069 7831 35127 7837
rect 35710 7828 35716 7840
rect 35768 7828 35774 7880
rect 38102 7868 38108 7880
rect 38063 7840 38108 7868
rect 38102 7828 38108 7840
rect 38160 7828 38166 7880
rect 11422 7800 11428 7812
rect 11383 7772 11428 7800
rect 11422 7760 11428 7772
rect 11480 7760 11486 7812
rect 23198 7760 23204 7812
rect 23256 7800 23262 7812
rect 28994 7800 29000 7812
rect 23256 7772 29000 7800
rect 23256 7760 23262 7772
rect 28994 7760 29000 7772
rect 29052 7760 29058 7812
rect 30006 7800 30012 7812
rect 29967 7772 30012 7800
rect 30006 7760 30012 7772
rect 30064 7760 30070 7812
rect 31941 7803 31999 7809
rect 31941 7769 31953 7803
rect 31987 7800 31999 7803
rect 32122 7800 32128 7812
rect 31987 7772 32128 7800
rect 31987 7769 31999 7772
rect 31941 7763 31999 7769
rect 32122 7760 32128 7772
rect 32180 7760 32186 7812
rect 37093 7803 37151 7809
rect 37093 7800 37105 7803
rect 34440 7772 37105 7800
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 3108 7704 3249 7732
rect 3108 7692 3114 7704
rect 3237 7701 3249 7704
rect 3283 7732 3295 7735
rect 15010 7732 15016 7744
rect 3283 7704 15016 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 20441 7735 20499 7741
rect 20441 7701 20453 7735
rect 20487 7732 20499 7735
rect 20622 7732 20628 7744
rect 20487 7704 20628 7732
rect 20487 7701 20499 7704
rect 20441 7695 20499 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 25041 7735 25099 7741
rect 25041 7701 25053 7735
rect 25087 7732 25099 7735
rect 25958 7732 25964 7744
rect 25087 7704 25964 7732
rect 25087 7701 25099 7704
rect 25041 7695 25099 7701
rect 25958 7692 25964 7704
rect 26016 7692 26022 7744
rect 28350 7692 28356 7744
rect 28408 7732 28414 7744
rect 34440 7732 34468 7772
rect 37093 7769 37105 7772
rect 37139 7769 37151 7803
rect 37093 7763 37151 7769
rect 35526 7732 35532 7744
rect 28408 7704 34468 7732
rect 35487 7704 35532 7732
rect 28408 7692 28414 7704
rect 35526 7692 35532 7704
rect 35584 7692 35590 7744
rect 36538 7732 36544 7744
rect 36499 7704 36544 7732
rect 36538 7692 36544 7704
rect 36596 7692 36602 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 7650 7488 7656 7540
rect 7708 7488 7714 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 18414 7528 18420 7540
rect 14783 7500 18420 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 26329 7531 26387 7537
rect 26329 7528 26341 7531
rect 26200 7500 26341 7528
rect 26200 7488 26206 7500
rect 26329 7497 26341 7500
rect 26375 7497 26387 7531
rect 28626 7528 28632 7540
rect 26329 7491 26387 7497
rect 28092 7500 28632 7528
rect 7469 7463 7527 7469
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 7668 7460 7696 7488
rect 28092 7469 28120 7500
rect 28626 7488 28632 7500
rect 28684 7488 28690 7540
rect 7515 7432 7696 7460
rect 7837 7463 7895 7469
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 7837 7429 7849 7463
rect 7883 7460 7895 7463
rect 8389 7463 8447 7469
rect 8389 7460 8401 7463
rect 7883 7432 8401 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8389 7429 8401 7432
rect 8435 7460 8447 7463
rect 28077 7463 28135 7469
rect 8435 7432 28028 7460
rect 8435 7429 8447 7432
rect 8389 7423 8447 7429
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 6564 7364 7665 7392
rect 6564 7336 6592 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 11514 7392 11520 7404
rect 11475 7364 11520 7392
rect 7653 7355 7711 7361
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 15194 7392 15200 7404
rect 15155 7364 15200 7392
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16114 7392 16120 7404
rect 15611 7364 16120 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 6546 7324 6552 7336
rect 6507 7296 6552 7324
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 7055 7296 13952 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 6825 7259 6883 7265
rect 6825 7256 6837 7259
rect 6696 7228 6837 7256
rect 6696 7216 6702 7228
rect 6825 7225 6837 7228
rect 6871 7225 6883 7259
rect 6825 7219 6883 7225
rect 11701 7191 11759 7197
rect 11701 7157 11713 7191
rect 11747 7188 11759 7191
rect 12618 7188 12624 7200
rect 11747 7160 12624 7188
rect 11747 7157 11759 7160
rect 11701 7151 11759 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 13924 7188 13952 7296
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 14240 7296 14289 7324
rect 14240 7284 14246 7296
rect 14277 7293 14289 7296
rect 14323 7324 14335 7327
rect 15396 7324 15424 7355
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 26142 7352 26148 7404
rect 26200 7392 26206 7404
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26200 7364 26985 7392
rect 26200 7352 26206 7364
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 14323 7296 15424 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 20162 7284 20168 7336
rect 20220 7324 20226 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 20220 7296 20361 7324
rect 20220 7284 20226 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 27893 7327 27951 7333
rect 27893 7324 27905 7327
rect 26292 7296 27905 7324
rect 26292 7284 26298 7296
rect 27893 7293 27905 7296
rect 27939 7293 27951 7327
rect 28000 7324 28028 7432
rect 28077 7429 28089 7463
rect 28123 7429 28135 7463
rect 28077 7423 28135 7429
rect 37829 7463 37887 7469
rect 37829 7429 37841 7463
rect 37875 7460 37887 7463
rect 38286 7460 38292 7472
rect 37875 7432 38292 7460
rect 37875 7429 37887 7432
rect 37829 7423 37887 7429
rect 38286 7420 38292 7432
rect 38344 7420 38350 7472
rect 34057 7395 34115 7401
rect 34057 7361 34069 7395
rect 34103 7392 34115 7395
rect 37182 7392 37188 7404
rect 34103 7364 37188 7392
rect 34103 7361 34115 7364
rect 34057 7355 34115 7361
rect 37182 7352 37188 7364
rect 37240 7352 37246 7404
rect 29362 7324 29368 7336
rect 28000 7296 29368 7324
rect 27893 7287 27951 7293
rect 29362 7284 29368 7296
rect 29420 7284 29426 7336
rect 35621 7327 35679 7333
rect 35621 7293 35633 7327
rect 35667 7324 35679 7327
rect 36170 7324 36176 7336
rect 35667 7296 36176 7324
rect 35667 7293 35679 7296
rect 35621 7287 35679 7293
rect 36170 7284 36176 7296
rect 36228 7284 36234 7336
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 14056 7228 14565 7256
rect 14056 7216 14062 7228
rect 14553 7225 14565 7228
rect 14599 7256 14611 7259
rect 14826 7256 14832 7268
rect 14599 7228 14832 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 19334 7256 19340 7268
rect 14936 7228 19340 7256
rect 14936 7188 14964 7228
rect 19334 7216 19340 7228
rect 19392 7216 19398 7268
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 20588 7228 20637 7256
rect 20588 7216 20594 7228
rect 20625 7225 20637 7228
rect 20671 7256 20683 7259
rect 21082 7256 21088 7268
rect 20671 7228 21088 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 21082 7216 21088 7228
rect 21140 7216 21146 7268
rect 26786 7216 26792 7268
rect 26844 7256 26850 7268
rect 26844 7228 28764 7256
rect 26844 7216 26850 7228
rect 16114 7188 16120 7200
rect 13924 7160 14964 7188
rect 16075 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 27157 7191 27215 7197
rect 27157 7157 27169 7191
rect 27203 7188 27215 7191
rect 27798 7188 27804 7200
rect 27203 7160 27804 7188
rect 27203 7157 27215 7160
rect 27157 7151 27215 7157
rect 27798 7148 27804 7160
rect 27856 7148 27862 7200
rect 28736 7188 28764 7228
rect 28994 7216 29000 7268
rect 29052 7256 29058 7268
rect 37645 7259 37703 7265
rect 37645 7256 37657 7259
rect 29052 7228 37657 7256
rect 29052 7216 29058 7228
rect 37645 7225 37657 7228
rect 37691 7225 37703 7259
rect 37645 7219 37703 7225
rect 34330 7188 34336 7200
rect 28736 7160 34336 7188
rect 34330 7148 34336 7160
rect 34388 7148 34394 7200
rect 34606 7188 34612 7200
rect 34567 7160 34612 7188
rect 34606 7148 34612 7160
rect 34664 7148 34670 7200
rect 35894 7148 35900 7200
rect 35952 7188 35958 7200
rect 36081 7191 36139 7197
rect 36081 7188 36093 7191
rect 35952 7160 36093 7188
rect 35952 7148 35958 7160
rect 36081 7157 36093 7160
rect 36127 7157 36139 7191
rect 36081 7151 36139 7157
rect 36725 7191 36783 7197
rect 36725 7157 36737 7191
rect 36771 7188 36783 7191
rect 38102 7188 38108 7200
rect 36771 7160 38108 7188
rect 36771 7157 36783 7160
rect 36725 7151 36783 7157
rect 38102 7148 38108 7160
rect 38160 7148 38166 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 14826 6984 14832 6996
rect 14787 6956 14832 6984
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 16114 6944 16120 6996
rect 16172 6984 16178 6996
rect 26786 6984 26792 6996
rect 16172 6956 26792 6984
rect 16172 6944 16178 6956
rect 26786 6944 26792 6956
rect 26844 6944 26850 6996
rect 33778 6984 33784 6996
rect 26896 6956 33784 6984
rect 16853 6919 16911 6925
rect 16853 6885 16865 6919
rect 16899 6885 16911 6919
rect 16853 6879 16911 6885
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6696 6820 7113 6848
rect 6696 6808 6702 6820
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 16022 6848 16028 6860
rect 15983 6820 16028 6848
rect 7101 6811 7159 6817
rect 16022 6808 16028 6820
rect 16080 6848 16086 6860
rect 16868 6848 16896 6879
rect 18414 6876 18420 6928
rect 18472 6916 18478 6928
rect 26896 6916 26924 6956
rect 33778 6944 33784 6956
rect 33836 6944 33842 6996
rect 18472 6888 26924 6916
rect 31757 6919 31815 6925
rect 18472 6876 18478 6888
rect 31757 6885 31769 6919
rect 31803 6885 31815 6919
rect 31757 6879 31815 6885
rect 16080 6820 16896 6848
rect 20349 6851 20407 6857
rect 16080 6808 16086 6820
rect 20349 6817 20361 6851
rect 20395 6848 20407 6851
rect 20395 6820 22094 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 20806 6780 20812 6792
rect 19567 6752 20812 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6780 21051 6783
rect 21082 6780 21088 6792
rect 21039 6752 21088 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 22066 6780 22094 6820
rect 24946 6808 24952 6860
rect 25004 6848 25010 6860
rect 25041 6851 25099 6857
rect 25041 6848 25053 6851
rect 25004 6820 25053 6848
rect 25004 6808 25010 6820
rect 25041 6817 25053 6820
rect 25087 6817 25099 6851
rect 30006 6848 30012 6860
rect 25041 6811 25099 6817
rect 25240 6820 30012 6848
rect 25240 6780 25268 6820
rect 30006 6808 30012 6820
rect 30064 6808 30070 6860
rect 31205 6851 31263 6857
rect 31205 6817 31217 6851
rect 31251 6848 31263 6851
rect 31570 6848 31576 6860
rect 31251 6820 31576 6848
rect 31251 6817 31263 6820
rect 31205 6811 31263 6817
rect 31570 6808 31576 6820
rect 31628 6848 31634 6860
rect 31772 6848 31800 6879
rect 32122 6848 32128 6860
rect 31628 6820 31800 6848
rect 32083 6820 32128 6848
rect 31628 6808 31634 6820
rect 32122 6808 32128 6820
rect 32180 6808 32186 6860
rect 36722 6808 36728 6860
rect 36780 6848 36786 6860
rect 36780 6820 37872 6848
rect 36780 6808 36786 6820
rect 27614 6780 27620 6792
rect 22066 6752 25268 6780
rect 27575 6752 27620 6780
rect 27614 6740 27620 6752
rect 27672 6780 27678 6792
rect 28261 6783 28319 6789
rect 28261 6780 28273 6783
rect 27672 6752 28273 6780
rect 27672 6740 27678 6752
rect 28261 6749 28273 6752
rect 28307 6749 28319 6783
rect 35253 6783 35311 6789
rect 35253 6780 35265 6783
rect 28261 6743 28319 6749
rect 31726 6752 35265 6780
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 16577 6715 16635 6721
rect 16577 6712 16589 6715
rect 16540 6684 16589 6712
rect 16540 6672 16546 6684
rect 16577 6681 16589 6684
rect 16623 6681 16635 6715
rect 19978 6712 19984 6724
rect 16577 6675 16635 6681
rect 17052 6684 19564 6712
rect 19939 6684 19984 6712
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5350 6644 5356 6656
rect 5307 6616 5356 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 17052 6653 17080 6684
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 19426 6644 19432 6656
rect 19383 6616 19432 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 19536 6644 19564 6684
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 20162 6712 20168 6724
rect 20123 6684 20168 6712
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 24854 6712 24860 6724
rect 24815 6684 24860 6712
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 31726 6712 31754 6752
rect 35253 6749 35265 6752
rect 35299 6780 35311 6783
rect 35434 6780 35440 6792
rect 35299 6752 35440 6780
rect 35299 6749 35311 6752
rect 35253 6743 35311 6749
rect 35434 6740 35440 6752
rect 35492 6740 35498 6792
rect 36633 6783 36691 6789
rect 36633 6749 36645 6783
rect 36679 6780 36691 6783
rect 37185 6783 37243 6789
rect 37185 6780 37197 6783
rect 36679 6752 37197 6780
rect 36679 6749 36691 6752
rect 36633 6743 36691 6749
rect 37185 6749 37197 6752
rect 37231 6780 37243 6783
rect 37366 6780 37372 6792
rect 37231 6752 37372 6780
rect 37231 6749 37243 6752
rect 37185 6743 37243 6749
rect 37366 6740 37372 6752
rect 37424 6740 37430 6792
rect 37844 6789 37872 6820
rect 37829 6783 37887 6789
rect 37829 6749 37841 6783
rect 37875 6749 37887 6783
rect 37829 6743 37887 6749
rect 38470 6740 38476 6792
rect 38528 6740 38534 6792
rect 38488 6712 38516 6740
rect 26896 6684 31754 6712
rect 37384 6684 38516 6712
rect 26896 6644 26924 6684
rect 19536 6616 26924 6644
rect 27801 6647 27859 6653
rect 27801 6613 27813 6647
rect 27847 6644 27859 6647
rect 28166 6644 28172 6656
rect 27847 6616 28172 6644
rect 27847 6613 27859 6616
rect 27801 6607 27859 6613
rect 28166 6604 28172 6616
rect 28224 6604 28230 6656
rect 29917 6647 29975 6653
rect 29917 6613 29929 6647
rect 29963 6644 29975 6647
rect 30006 6644 30012 6656
rect 29963 6616 30012 6644
rect 29963 6613 29975 6616
rect 29917 6607 29975 6613
rect 30006 6604 30012 6616
rect 30064 6604 30070 6656
rect 30558 6644 30564 6656
rect 30519 6616 30564 6644
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 31665 6647 31723 6653
rect 31665 6613 31677 6647
rect 31711 6644 31723 6647
rect 32214 6644 32220 6656
rect 31711 6616 32220 6644
rect 31711 6613 31723 6616
rect 31665 6607 31723 6613
rect 32214 6604 32220 6616
rect 32272 6604 32278 6656
rect 32582 6644 32588 6656
rect 32543 6616 32588 6644
rect 32582 6604 32588 6616
rect 32640 6604 32646 6656
rect 33229 6647 33287 6653
rect 33229 6613 33241 6647
rect 33275 6644 33287 6647
rect 33318 6644 33324 6656
rect 33275 6616 33324 6644
rect 33275 6613 33287 6616
rect 33229 6607 33287 6613
rect 33318 6604 33324 6616
rect 33376 6604 33382 6656
rect 33781 6647 33839 6653
rect 33781 6613 33793 6647
rect 33827 6644 33839 6647
rect 33962 6644 33968 6656
rect 33827 6616 33968 6644
rect 33827 6613 33839 6616
rect 33781 6607 33839 6613
rect 33962 6604 33968 6616
rect 34020 6604 34026 6656
rect 34514 6604 34520 6656
rect 34572 6644 34578 6656
rect 34701 6647 34759 6653
rect 34701 6644 34713 6647
rect 34572 6616 34713 6644
rect 34572 6604 34578 6616
rect 34701 6613 34713 6616
rect 34747 6613 34759 6647
rect 34701 6607 34759 6613
rect 35802 6604 35808 6656
rect 35860 6644 35866 6656
rect 37384 6653 37412 6684
rect 36081 6647 36139 6653
rect 36081 6644 36093 6647
rect 35860 6616 36093 6644
rect 35860 6604 35866 6616
rect 36081 6613 36093 6616
rect 36127 6613 36139 6647
rect 36081 6607 36139 6613
rect 37369 6647 37427 6653
rect 37369 6613 37381 6647
rect 37415 6613 37427 6647
rect 37369 6607 37427 6613
rect 38013 6647 38071 6653
rect 38013 6613 38025 6647
rect 38059 6644 38071 6647
rect 38470 6644 38476 6656
rect 38059 6616 38476 6644
rect 38059 6613 38071 6616
rect 38013 6607 38071 6613
rect 38470 6604 38476 6616
rect 38528 6604 38534 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 25682 6440 25688 6452
rect 3835 6412 25688 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 25682 6400 25688 6412
rect 25740 6400 25746 6452
rect 36725 6443 36783 6449
rect 36725 6409 36737 6443
rect 36771 6440 36783 6443
rect 37734 6440 37740 6452
rect 36771 6412 37740 6440
rect 36771 6409 36783 6412
rect 36725 6403 36783 6409
rect 37734 6400 37740 6412
rect 37792 6400 37798 6452
rect 4341 6375 4399 6381
rect 4341 6341 4353 6375
rect 4387 6372 4399 6375
rect 5258 6372 5264 6384
rect 4387 6344 5264 6372
rect 4387 6341 4399 6344
rect 4341 6335 4399 6341
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 3016 6208 3341 6236
rect 3016 6196 3022 6208
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 3329 6199 3387 6205
rect 3697 6171 3755 6177
rect 3697 6137 3709 6171
rect 3743 6168 3755 6171
rect 4356 6168 4384 6335
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 15562 6372 15568 6384
rect 15523 6344 15568 6372
rect 15562 6332 15568 6344
rect 15620 6332 15626 6384
rect 16669 6375 16727 6381
rect 16669 6341 16681 6375
rect 16715 6372 16727 6375
rect 16758 6372 16764 6384
rect 16715 6344 16764 6372
rect 16715 6341 16727 6344
rect 16669 6335 16727 6341
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 16960 6344 17724 6372
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 16482 6304 16488 6316
rect 15896 6276 16488 6304
rect 15896 6264 15902 6276
rect 16482 6264 16488 6276
rect 16540 6304 16546 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16540 6276 16865 6304
rect 16540 6264 16546 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 15010 6196 15016 6248
rect 15068 6236 15074 6248
rect 16960 6236 16988 6344
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17083 6276 17632 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 15068 6208 16988 6236
rect 15068 6196 15074 6208
rect 3743 6140 4384 6168
rect 3743 6137 3755 6140
rect 3697 6131 3755 6137
rect 1489 6103 1547 6109
rect 1489 6069 1501 6103
rect 1535 6100 1547 6103
rect 1578 6100 1584 6112
rect 1535 6072 1584 6100
rect 1535 6069 1547 6072
rect 1489 6063 1547 6069
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2498 6100 2504 6112
rect 2459 6072 2504 6100
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5442 6100 5448 6112
rect 5403 6072 5448 6100
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 15010 6100 15016 6112
rect 14971 6072 15016 6100
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 17604 6109 17632 6276
rect 17696 6168 17724 6344
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 27614 6372 27620 6384
rect 19392 6344 27620 6372
rect 19392 6332 19398 6344
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 35526 6372 35532 6384
rect 35268 6344 35532 6372
rect 35268 6313 35296 6344
rect 35526 6332 35532 6344
rect 35584 6372 35590 6384
rect 37826 6372 37832 6384
rect 35584 6344 36860 6372
rect 37787 6344 37832 6372
rect 35584 6332 35590 6344
rect 35253 6307 35311 6313
rect 35253 6273 35265 6307
rect 35299 6273 35311 6307
rect 35253 6267 35311 6273
rect 35618 6264 35624 6316
rect 35676 6304 35682 6316
rect 36081 6307 36139 6313
rect 36081 6304 36093 6307
rect 35676 6276 36093 6304
rect 35676 6264 35682 6276
rect 36081 6273 36093 6276
rect 36127 6273 36139 6307
rect 36081 6267 36139 6273
rect 36170 6264 36176 6316
rect 36228 6304 36234 6316
rect 36541 6307 36599 6313
rect 36541 6304 36553 6307
rect 36228 6276 36553 6304
rect 36228 6264 36234 6276
rect 36541 6273 36553 6276
rect 36587 6304 36599 6307
rect 36722 6304 36728 6316
rect 36587 6276 36728 6304
rect 36587 6273 36599 6276
rect 36541 6267 36599 6273
rect 36722 6264 36728 6276
rect 36780 6264 36786 6316
rect 19150 6196 19156 6248
rect 19208 6236 19214 6248
rect 29822 6236 29828 6248
rect 19208 6208 29828 6236
rect 19208 6196 19214 6208
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 34793 6239 34851 6245
rect 34793 6205 34805 6239
rect 34839 6236 34851 6239
rect 35636 6236 35664 6264
rect 34839 6208 35664 6236
rect 36832 6236 36860 6344
rect 37826 6332 37832 6344
rect 37884 6332 37890 6384
rect 37366 6264 37372 6316
rect 37424 6304 37430 6316
rect 39574 6304 39580 6316
rect 37424 6276 39580 6304
rect 37424 6264 37430 6276
rect 39574 6264 39580 6276
rect 39632 6264 39638 6316
rect 39850 6236 39856 6248
rect 36832 6208 39856 6236
rect 34839 6205 34851 6208
rect 34793 6199 34851 6205
rect 39850 6196 39856 6208
rect 39908 6196 39914 6248
rect 27246 6168 27252 6180
rect 17696 6140 27252 6168
rect 27246 6128 27252 6140
rect 27304 6128 27310 6180
rect 30098 6128 30104 6180
rect 30156 6168 30162 6180
rect 31481 6171 31539 6177
rect 31481 6168 31493 6171
rect 30156 6140 31493 6168
rect 30156 6128 30162 6140
rect 31481 6137 31493 6140
rect 31527 6137 31539 6171
rect 31481 6131 31539 6137
rect 35437 6171 35495 6177
rect 35437 6137 35449 6171
rect 35483 6168 35495 6171
rect 37274 6168 37280 6180
rect 35483 6140 37280 6168
rect 35483 6137 35495 6140
rect 35437 6131 35495 6137
rect 37274 6128 37280 6140
rect 37332 6128 37338 6180
rect 17589 6103 17647 6109
rect 17589 6069 17601 6103
rect 17635 6100 17647 6103
rect 18690 6100 18696 6112
rect 17635 6072 18696 6100
rect 17635 6069 17647 6072
rect 17589 6063 17647 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 29638 6100 29644 6112
rect 29599 6072 29644 6100
rect 29638 6060 29644 6072
rect 29696 6060 29702 6112
rect 30466 6100 30472 6112
rect 30427 6072 30472 6100
rect 30466 6060 30472 6072
rect 30524 6060 30530 6112
rect 30926 6100 30932 6112
rect 30887 6072 30932 6100
rect 30926 6060 30932 6072
rect 30984 6060 30990 6112
rect 31386 6060 31392 6112
rect 31444 6100 31450 6112
rect 32125 6103 32183 6109
rect 32125 6100 32137 6103
rect 31444 6072 32137 6100
rect 31444 6060 31450 6072
rect 32125 6069 32137 6072
rect 32171 6069 32183 6103
rect 32858 6100 32864 6112
rect 32819 6072 32864 6100
rect 32125 6063 32183 6069
rect 32858 6060 32864 6072
rect 32916 6060 32922 6112
rect 33502 6060 33508 6112
rect 33560 6100 33566 6112
rect 33597 6103 33655 6109
rect 33597 6100 33609 6103
rect 33560 6072 33609 6100
rect 33560 6060 33566 6072
rect 33597 6069 33609 6072
rect 33643 6069 33655 6103
rect 33597 6063 33655 6069
rect 34054 6060 34060 6112
rect 34112 6100 34118 6112
rect 34149 6103 34207 6109
rect 34149 6100 34161 6103
rect 34112 6072 34161 6100
rect 34112 6060 34118 6072
rect 34149 6069 34161 6072
rect 34195 6069 34207 6103
rect 34149 6063 34207 6069
rect 35897 6103 35955 6109
rect 35897 6069 35909 6103
rect 35943 6100 35955 6103
rect 35986 6100 35992 6112
rect 35943 6072 35992 6100
rect 35943 6069 35955 6072
rect 35897 6063 35955 6069
rect 35986 6060 35992 6072
rect 36044 6060 36050 6112
rect 37734 6100 37740 6112
rect 37695 6072 37740 6100
rect 37734 6060 37740 6072
rect 37792 6060 37798 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 4614 5896 4620 5908
rect 3835 5868 4620 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 16206 5896 16212 5908
rect 16167 5868 16212 5896
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 18690 5856 18696 5908
rect 18748 5896 18754 5908
rect 18748 5868 22094 5896
rect 18748 5856 18754 5868
rect 22066 5828 22094 5868
rect 25038 5856 25044 5908
rect 25096 5896 25102 5908
rect 25133 5899 25191 5905
rect 25133 5896 25145 5899
rect 25096 5868 25145 5896
rect 25096 5856 25102 5868
rect 25133 5865 25145 5868
rect 25179 5896 25191 5899
rect 25406 5896 25412 5908
rect 25179 5868 25412 5896
rect 25179 5865 25191 5868
rect 25133 5859 25191 5865
rect 25406 5856 25412 5868
rect 25464 5856 25470 5908
rect 26510 5856 26516 5908
rect 26568 5896 26574 5908
rect 26694 5896 26700 5908
rect 26568 5868 26700 5896
rect 26568 5856 26574 5868
rect 26694 5856 26700 5868
rect 26752 5896 26758 5908
rect 26881 5899 26939 5905
rect 26881 5896 26893 5899
rect 26752 5868 26893 5896
rect 26752 5856 26758 5868
rect 26881 5865 26893 5868
rect 26927 5865 26939 5899
rect 26881 5859 26939 5865
rect 29822 5856 29828 5908
rect 29880 5896 29886 5908
rect 30009 5899 30067 5905
rect 30009 5896 30021 5899
rect 29880 5868 30021 5896
rect 29880 5856 29886 5868
rect 30009 5865 30021 5868
rect 30055 5865 30067 5899
rect 30650 5896 30656 5908
rect 30611 5868 30656 5896
rect 30009 5859 30067 5865
rect 30650 5856 30656 5868
rect 30708 5856 30714 5908
rect 31297 5899 31355 5905
rect 31297 5865 31309 5899
rect 31343 5896 31355 5899
rect 31662 5896 31668 5908
rect 31343 5868 31668 5896
rect 31343 5865 31355 5868
rect 31297 5859 31355 5865
rect 31662 5856 31668 5868
rect 31720 5856 31726 5908
rect 32674 5856 32680 5908
rect 32732 5896 32738 5908
rect 33321 5899 33379 5905
rect 33321 5896 33333 5899
rect 32732 5868 33333 5896
rect 32732 5856 32738 5868
rect 33321 5865 33333 5868
rect 33367 5865 33379 5899
rect 33321 5859 33379 5865
rect 33778 5856 33784 5908
rect 33836 5896 33842 5908
rect 33965 5899 34023 5905
rect 33965 5896 33977 5899
rect 33836 5868 33977 5896
rect 33836 5856 33842 5868
rect 33965 5865 33977 5868
rect 34011 5865 34023 5899
rect 33965 5859 34023 5865
rect 34790 5856 34796 5908
rect 34848 5896 34854 5908
rect 34885 5899 34943 5905
rect 34885 5896 34897 5899
rect 34848 5868 34897 5896
rect 34848 5856 34854 5868
rect 34885 5865 34897 5868
rect 34931 5865 34943 5899
rect 34885 5859 34943 5865
rect 36078 5856 36084 5908
rect 36136 5896 36142 5908
rect 37921 5899 37979 5905
rect 37921 5896 37933 5899
rect 36136 5868 37933 5896
rect 36136 5856 36142 5868
rect 37921 5865 37933 5868
rect 37967 5865 37979 5899
rect 37921 5859 37979 5865
rect 35526 5828 35532 5840
rect 22066 5800 35532 5828
rect 35526 5788 35532 5800
rect 35584 5788 35590 5840
rect 36449 5831 36507 5837
rect 36449 5797 36461 5831
rect 36495 5828 36507 5831
rect 39298 5828 39304 5840
rect 36495 5800 39304 5828
rect 36495 5797 36507 5800
rect 36449 5791 36507 5797
rect 39298 5788 39304 5800
rect 39356 5788 39362 5840
rect 10962 5720 10968 5772
rect 11020 5760 11026 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 11020 5732 12541 5760
rect 11020 5720 11026 5732
rect 12529 5729 12541 5732
rect 12575 5760 12587 5763
rect 14274 5760 14280 5772
rect 12575 5732 14280 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 24762 5720 24768 5772
rect 24820 5760 24826 5772
rect 37734 5760 37740 5772
rect 24820 5732 37740 5760
rect 24820 5720 24826 5732
rect 37734 5720 37740 5732
rect 37792 5720 37798 5772
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4203 5664 4721 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4709 5661 4721 5664
rect 4755 5692 4767 5695
rect 18874 5692 18880 5704
rect 4755 5664 18880 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 25682 5692 25688 5704
rect 25643 5664 25688 5692
rect 25682 5652 25688 5664
rect 25740 5692 25746 5704
rect 26329 5695 26387 5701
rect 26329 5692 26341 5695
rect 25740 5664 26341 5692
rect 25740 5652 25746 5664
rect 26329 5661 26341 5664
rect 26375 5661 26387 5695
rect 26329 5655 26387 5661
rect 30101 5695 30159 5701
rect 30101 5661 30113 5695
rect 30147 5692 30159 5695
rect 30650 5692 30656 5704
rect 30147 5664 30656 5692
rect 30147 5661 30159 5664
rect 30101 5655 30159 5661
rect 30650 5652 30656 5664
rect 30708 5652 30714 5704
rect 33505 5695 33563 5701
rect 33505 5692 33517 5695
rect 33244 5664 33517 5692
rect 1762 5584 1768 5636
rect 1820 5624 1826 5636
rect 2501 5627 2559 5633
rect 2501 5624 2513 5627
rect 1820 5596 2513 5624
rect 1820 5584 1826 5596
rect 2501 5593 2513 5596
rect 2547 5593 2559 5627
rect 2501 5587 2559 5593
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 3973 5627 4031 5633
rect 3973 5624 3985 5627
rect 3016 5596 3985 5624
rect 3016 5584 3022 5596
rect 3973 5593 3985 5596
rect 4019 5593 4031 5627
rect 3973 5587 4031 5593
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 12621 5627 12679 5633
rect 12621 5624 12633 5627
rect 7064 5596 12633 5624
rect 7064 5584 7070 5596
rect 12621 5593 12633 5596
rect 12667 5593 12679 5627
rect 24854 5624 24860 5636
rect 12621 5587 12679 5593
rect 13096 5596 24860 5624
rect 1394 5556 1400 5568
rect 1355 5528 1400 5556
rect 1394 5516 1400 5528
rect 1452 5516 1458 5568
rect 1670 5516 1676 5568
rect 1728 5556 1734 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1728 5528 1961 5556
rect 1728 5516 1734 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 1949 5519 2007 5525
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3694 5556 3700 5568
rect 3283 5528 3700 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 4120 5528 5181 5556
rect 4120 5516 4126 5528
rect 5169 5525 5181 5528
rect 5215 5525 5227 5559
rect 5718 5556 5724 5568
rect 5679 5528 5724 5556
rect 5169 5519 5227 5525
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6362 5556 6368 5568
rect 6323 5528 6368 5556
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 8018 5556 8024 5568
rect 7979 5528 8024 5556
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11054 5556 11060 5568
rect 11015 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13096 5565 13124 5596
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 33244 5568 33272 5664
rect 33505 5661 33517 5664
rect 33551 5661 33563 5695
rect 33505 5655 33563 5661
rect 34054 5652 34060 5704
rect 34112 5692 34118 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 34112 5664 34713 5692
rect 34112 5652 34118 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 35434 5692 35440 5704
rect 35395 5664 35440 5692
rect 34701 5655 34759 5661
rect 35434 5652 35440 5664
rect 35492 5652 35498 5704
rect 36630 5692 36636 5704
rect 36591 5664 36636 5692
rect 36630 5652 36636 5664
rect 36688 5652 36694 5704
rect 37090 5692 37096 5704
rect 37051 5664 37096 5692
rect 37090 5652 37096 5664
rect 37148 5652 37154 5704
rect 35802 5584 35808 5636
rect 35860 5624 35866 5636
rect 38010 5624 38016 5636
rect 35860 5596 38016 5624
rect 35860 5584 35866 5596
rect 38010 5584 38016 5596
rect 38068 5584 38074 5636
rect 13081 5559 13139 5565
rect 13081 5525 13093 5559
rect 13127 5525 13139 5559
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 13081 5519 13139 5525
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15654 5556 15660 5568
rect 15615 5528 15660 5556
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 20349 5559 20407 5565
rect 20349 5556 20361 5559
rect 20128 5528 20361 5556
rect 20128 5516 20134 5528
rect 20349 5525 20361 5528
rect 20395 5525 20407 5559
rect 20349 5519 20407 5525
rect 20898 5516 20904 5568
rect 20956 5556 20962 5568
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 20956 5528 21189 5556
rect 20956 5516 20962 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 21177 5519 21235 5525
rect 22097 5559 22155 5565
rect 22097 5525 22109 5559
rect 22143 5556 22155 5559
rect 22186 5556 22192 5568
rect 22143 5528 22192 5556
rect 22143 5525 22155 5528
rect 22097 5519 22155 5525
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 24578 5556 24584 5568
rect 24539 5528 24584 5556
rect 24578 5516 24584 5528
rect 24636 5516 24642 5568
rect 25869 5559 25927 5565
rect 25869 5525 25881 5559
rect 25915 5556 25927 5559
rect 26786 5556 26792 5568
rect 25915 5528 26792 5556
rect 25915 5525 25927 5528
rect 25869 5519 25927 5525
rect 26786 5516 26792 5528
rect 26844 5516 26850 5568
rect 28997 5559 29055 5565
rect 28997 5525 29009 5559
rect 29043 5556 29055 5559
rect 29730 5556 29736 5568
rect 29043 5528 29736 5556
rect 29043 5525 29055 5528
rect 28997 5519 29055 5525
rect 29730 5516 29736 5528
rect 29788 5516 29794 5568
rect 30650 5516 30656 5568
rect 30708 5556 30714 5568
rect 30926 5556 30932 5568
rect 30708 5528 30932 5556
rect 30708 5516 30714 5528
rect 30926 5516 30932 5528
rect 30984 5516 30990 5568
rect 31110 5516 31116 5568
rect 31168 5556 31174 5568
rect 31846 5556 31852 5568
rect 31168 5528 31852 5556
rect 31168 5516 31174 5528
rect 31846 5516 31852 5528
rect 31904 5556 31910 5568
rect 31941 5559 31999 5565
rect 31941 5556 31953 5559
rect 31904 5528 31953 5556
rect 31904 5516 31910 5528
rect 31941 5525 31953 5528
rect 31987 5525 31999 5559
rect 31941 5519 31999 5525
rect 32861 5559 32919 5565
rect 32861 5525 32873 5559
rect 32907 5556 32919 5559
rect 33226 5556 33232 5568
rect 32907 5528 33232 5556
rect 32907 5525 32919 5528
rect 32861 5519 32919 5525
rect 33226 5516 33232 5528
rect 33284 5516 33290 5568
rect 35621 5559 35679 5565
rect 35621 5525 35633 5559
rect 35667 5556 35679 5559
rect 36078 5556 36084 5568
rect 35667 5528 36084 5556
rect 35667 5525 35679 5528
rect 35621 5519 35679 5525
rect 36078 5516 36084 5528
rect 36136 5516 36142 5568
rect 37277 5559 37335 5565
rect 37277 5525 37289 5559
rect 37323 5556 37335 5559
rect 37550 5556 37556 5568
rect 37323 5528 37556 5556
rect 37323 5525 37335 5528
rect 37277 5519 37335 5525
rect 37550 5516 37556 5528
rect 37608 5516 37614 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 26050 5312 26056 5364
rect 26108 5352 26114 5364
rect 26329 5355 26387 5361
rect 26329 5352 26341 5355
rect 26108 5324 26341 5352
rect 26108 5312 26114 5324
rect 26329 5321 26341 5324
rect 26375 5352 26387 5355
rect 26602 5352 26608 5364
rect 26375 5324 26608 5352
rect 26375 5321 26387 5324
rect 26329 5315 26387 5321
rect 26602 5312 26608 5324
rect 26660 5312 26666 5364
rect 29270 5352 29276 5364
rect 29231 5324 29276 5352
rect 29270 5312 29276 5324
rect 29328 5312 29334 5364
rect 30009 5355 30067 5361
rect 30009 5321 30021 5355
rect 30055 5352 30067 5355
rect 30926 5352 30932 5364
rect 30055 5324 30932 5352
rect 30055 5321 30067 5324
rect 30009 5315 30067 5321
rect 30926 5312 30932 5324
rect 30984 5312 30990 5364
rect 32030 5312 32036 5364
rect 32088 5352 32094 5364
rect 32125 5355 32183 5361
rect 32125 5352 32137 5355
rect 32088 5324 32137 5352
rect 32088 5312 32094 5324
rect 32125 5321 32137 5324
rect 32171 5321 32183 5355
rect 32125 5315 32183 5321
rect 32398 5312 32404 5364
rect 32456 5352 32462 5364
rect 33045 5355 33103 5361
rect 33045 5352 33057 5355
rect 32456 5324 33057 5352
rect 32456 5312 32462 5324
rect 33045 5321 33057 5324
rect 33091 5321 33103 5355
rect 33045 5315 33103 5321
rect 33594 5312 33600 5364
rect 33652 5352 33658 5364
rect 33873 5355 33931 5361
rect 33873 5352 33885 5355
rect 33652 5324 33885 5352
rect 33652 5312 33658 5324
rect 33873 5321 33885 5324
rect 33919 5321 33931 5355
rect 33873 5315 33931 5321
rect 34422 5312 34428 5364
rect 34480 5352 34486 5364
rect 34885 5355 34943 5361
rect 34885 5352 34897 5355
rect 34480 5324 34897 5352
rect 34480 5312 34486 5324
rect 34885 5321 34897 5324
rect 34931 5321 34943 5355
rect 34885 5315 34943 5321
rect 37369 5355 37427 5361
rect 37369 5321 37381 5355
rect 37415 5352 37427 5355
rect 37826 5352 37832 5364
rect 37415 5324 37832 5352
rect 37415 5321 37427 5324
rect 37369 5315 37427 5321
rect 37826 5312 37832 5324
rect 37884 5312 37890 5364
rect 21634 5244 21640 5296
rect 21692 5284 21698 5296
rect 26878 5284 26884 5296
rect 21692 5256 26884 5284
rect 21692 5244 21698 5256
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 27430 5244 27436 5296
rect 27488 5284 27494 5296
rect 31478 5284 31484 5296
rect 27488 5256 31484 5284
rect 27488 5244 27494 5256
rect 31478 5244 31484 5256
rect 31536 5244 31542 5296
rect 32766 5244 32772 5296
rect 32824 5284 32830 5296
rect 34793 5287 34851 5293
rect 34793 5284 34805 5287
rect 32824 5256 34805 5284
rect 32824 5244 32830 5256
rect 34793 5253 34805 5256
rect 34839 5253 34851 5287
rect 35434 5284 35440 5296
rect 35395 5256 35440 5284
rect 34793 5247 34851 5253
rect 35434 5244 35440 5256
rect 35492 5244 35498 5296
rect 29270 5176 29276 5228
rect 29328 5216 29334 5228
rect 29825 5219 29883 5225
rect 29825 5216 29837 5219
rect 29328 5188 29837 5216
rect 29328 5176 29334 5188
rect 29825 5185 29837 5188
rect 29871 5185 29883 5219
rect 29825 5179 29883 5185
rect 31389 5219 31447 5225
rect 31389 5185 31401 5219
rect 31435 5216 31447 5219
rect 31662 5216 31668 5228
rect 31435 5188 31668 5216
rect 31435 5185 31447 5188
rect 31389 5179 31447 5185
rect 31662 5176 31668 5188
rect 31720 5176 31726 5228
rect 31846 5176 31852 5228
rect 31904 5216 31910 5228
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31904 5188 32321 5216
rect 31904 5176 31910 5188
rect 32309 5185 32321 5188
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 32858 5176 32864 5228
rect 32916 5216 32922 5228
rect 33229 5219 33287 5225
rect 33229 5216 33241 5219
rect 32916 5188 33241 5216
rect 32916 5176 32922 5188
rect 33229 5185 33241 5188
rect 33275 5185 33287 5219
rect 33229 5179 33287 5185
rect 33962 5176 33968 5228
rect 34020 5216 34026 5228
rect 34057 5219 34115 5225
rect 34057 5216 34069 5219
rect 34020 5188 34069 5216
rect 34020 5176 34026 5188
rect 34057 5185 34069 5188
rect 34103 5185 34115 5219
rect 34057 5179 34115 5185
rect 35621 5219 35679 5225
rect 35621 5185 35633 5219
rect 35667 5185 35679 5219
rect 36446 5216 36452 5228
rect 36407 5188 36452 5216
rect 35621 5179 35679 5185
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 22278 5148 22284 5160
rect 8352 5120 22284 5148
rect 8352 5108 8358 5120
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 30374 5108 30380 5160
rect 30432 5148 30438 5160
rect 30469 5151 30527 5157
rect 30469 5148 30481 5151
rect 30432 5120 30481 5148
rect 30432 5108 30438 5120
rect 30469 5117 30481 5120
rect 30515 5117 30527 5151
rect 35636 5148 35664 5179
rect 36446 5176 36452 5188
rect 36504 5176 36510 5228
rect 38102 5216 38108 5228
rect 38063 5188 38108 5216
rect 38102 5176 38108 5188
rect 38160 5176 38166 5228
rect 30469 5111 30527 5117
rect 30576 5120 35664 5148
rect 4525 5083 4583 5089
rect 4525 5049 4537 5083
rect 4571 5080 4583 5083
rect 4706 5080 4712 5092
rect 4571 5052 4712 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 23382 5080 23388 5092
rect 6144 5052 23388 5080
rect 6144 5040 6150 5052
rect 23382 5040 23388 5052
rect 23440 5040 23446 5092
rect 24854 5040 24860 5092
rect 24912 5080 24918 5092
rect 30576 5080 30604 5120
rect 33502 5080 33508 5092
rect 24912 5052 30604 5080
rect 31036 5052 33508 5080
rect 24912 5040 24918 5052
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 2593 5015 2651 5021
rect 2593 4981 2605 5015
rect 2639 5012 2651 5015
rect 2774 5012 2780 5024
rect 2639 4984 2780 5012
rect 2639 4981 2651 4984
rect 2593 4975 2651 4981
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 3234 5012 3240 5024
rect 3191 4984 3240 5012
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3786 5012 3792 5024
rect 3747 4984 3792 5012
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4672 4984 4997 5012
rect 4672 4972 4678 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5684 4984 5733 5012
rect 5684 4972 5690 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 6454 5012 6460 5024
rect 6415 4984 6460 5012
rect 5721 4975 5779 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 7190 5012 7196 5024
rect 7151 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 7929 5015 7987 5021
rect 7929 5012 7941 5015
rect 7800 4984 7941 5012
rect 7800 4972 7806 4984
rect 7929 4981 7941 4984
rect 7975 4981 7987 5015
rect 8478 5012 8484 5024
rect 8439 4984 8484 5012
rect 7929 4975 7987 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 9030 5012 9036 5024
rect 8991 4984 9036 5012
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 9272 4984 9597 5012
rect 9272 4972 9278 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 9732 4984 10149 5012
rect 9732 4972 9738 4984
rect 10137 4981 10149 4984
rect 10183 4981 10195 5015
rect 10137 4975 10195 4981
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 10689 5015 10747 5021
rect 10689 5012 10701 5015
rect 10652 4984 10701 5012
rect 10652 4972 10658 4984
rect 10689 4981 10701 4984
rect 10735 4981 10747 5015
rect 10689 4975 10747 4981
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11572 4984 11713 5012
rect 11572 4972 11578 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11940 4984 12265 5012
rect 11940 4972 11946 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12584 4984 12817 5012
rect 12584 4972 12590 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 13354 5012 13360 5024
rect 13315 4984 13360 5012
rect 12805 4975 12863 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13998 5012 14004 5024
rect 13959 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14826 5012 14832 5024
rect 14787 4984 14832 5012
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 15746 5012 15752 5024
rect 15707 4984 15752 5012
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 16666 5012 16672 5024
rect 16627 4984 16672 5012
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 17218 5012 17224 5024
rect 17179 4984 17224 5012
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 18322 5012 18328 5024
rect 18283 4984 18328 5012
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 18966 5012 18972 5024
rect 18927 4984 18972 5012
rect 18966 4972 18972 4984
rect 19024 4972 19030 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 19392 4984 19441 5012
rect 19392 4972 19398 4984
rect 19429 4981 19441 4984
rect 19475 4981 19487 5015
rect 20438 5012 20444 5024
rect 20399 4984 20444 5012
rect 19429 4975 19487 4981
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 21085 5015 21143 5021
rect 21085 4981 21097 5015
rect 21131 5012 21143 5015
rect 21174 5012 21180 5024
rect 21131 4984 21180 5012
rect 21131 4981 21143 4984
rect 21085 4975 21143 4981
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 21450 4972 21456 5024
rect 21508 5012 21514 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21508 4984 21833 5012
rect 21508 4972 21514 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 22462 5012 22468 5024
rect 22423 4984 22468 5012
rect 21821 4975 21879 4981
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 22646 4972 22652 5024
rect 22704 5012 22710 5024
rect 22925 5015 22983 5021
rect 22925 5012 22937 5015
rect 22704 4984 22937 5012
rect 22704 4972 22710 4984
rect 22925 4981 22937 4984
rect 22971 4981 22983 5015
rect 23750 5012 23756 5024
rect 23711 4984 23756 5012
rect 22925 4975 22983 4981
rect 23750 4972 23756 4984
rect 23808 4972 23814 5024
rect 24305 5015 24363 5021
rect 24305 4981 24317 5015
rect 24351 5012 24363 5015
rect 24394 5012 24400 5024
rect 24351 4984 24400 5012
rect 24351 4981 24363 4984
rect 24305 4975 24363 4981
rect 24394 4972 24400 4984
rect 24452 4972 24458 5024
rect 25038 5012 25044 5024
rect 24999 4984 25044 5012
rect 25038 4972 25044 4984
rect 25096 4972 25102 5024
rect 25777 5015 25835 5021
rect 25777 4981 25789 5015
rect 25823 5012 25835 5015
rect 26602 5012 26608 5024
rect 25823 4984 26608 5012
rect 25823 4981 25835 4984
rect 25777 4975 25835 4981
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 27522 5012 27528 5024
rect 27483 4984 27528 5012
rect 27522 4972 27528 4984
rect 27580 4972 27586 5024
rect 27982 5012 27988 5024
rect 27943 4984 27988 5012
rect 27982 4972 27988 4984
rect 28040 4972 28046 5024
rect 28718 5012 28724 5024
rect 28679 4984 28724 5012
rect 28718 4972 28724 4984
rect 28776 4972 28782 5024
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 31036 5012 31064 5052
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 33778 5040 33784 5092
rect 33836 5080 33842 5092
rect 37921 5083 37979 5089
rect 37921 5080 37933 5083
rect 33836 5052 37933 5080
rect 33836 5040 33842 5052
rect 37921 5049 37933 5052
rect 37967 5049 37979 5083
rect 37921 5043 37979 5049
rect 28868 4984 31064 5012
rect 31573 5015 31631 5021
rect 28868 4972 28874 4984
rect 31573 4981 31585 5015
rect 31619 5012 31631 5015
rect 31938 5012 31944 5024
rect 31619 4984 31944 5012
rect 31619 4981 31631 4984
rect 31573 4975 31631 4981
rect 31938 4972 31944 4984
rect 31996 4972 32002 5024
rect 36633 5015 36691 5021
rect 36633 4981 36645 5015
rect 36679 5012 36691 5015
rect 36814 5012 36820 5024
rect 36679 4984 36820 5012
rect 36679 4981 36691 4984
rect 36633 4975 36691 4981
rect 36814 4972 36820 4984
rect 36872 4972 36878 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 6086 4808 6092 4820
rect 5316 4780 6092 4808
rect 5316 4768 5322 4780
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 8294 4808 8300 4820
rect 8255 4780 8300 4808
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 12768 4780 14105 4808
rect 12768 4768 12774 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 20990 4808 20996 4820
rect 14093 4771 14151 4777
rect 15672 4780 20996 4808
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 2866 4740 2872 4752
rect 1627 4712 2872 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 3878 4740 3884 4752
rect 3791 4712 3884 4740
rect 3878 4700 3884 4712
rect 3936 4740 3942 4752
rect 8846 4740 8852 4752
rect 3936 4712 8852 4740
rect 3936 4700 3942 4712
rect 8846 4700 8852 4712
rect 8904 4700 8910 4752
rect 9585 4743 9643 4749
rect 9585 4709 9597 4743
rect 9631 4740 9643 4743
rect 15672 4740 15700 4780
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 25130 4808 25136 4820
rect 25091 4780 25136 4808
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 27430 4808 27436 4820
rect 26436 4780 27436 4808
rect 26234 4740 26240 4752
rect 9631 4712 15700 4740
rect 15764 4712 26240 4740
rect 9631 4709 9643 4712
rect 9585 4703 9643 4709
rect 8294 4672 8300 4684
rect 2884 4644 8300 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1578 4604 1584 4616
rect 1443 4576 1584 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 1820 4576 2053 4604
rect 1820 4564 1826 4576
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2685 4607 2743 4613
rect 2685 4604 2697 4607
rect 2556 4576 2697 4604
rect 2556 4564 2562 4576
rect 2685 4573 2697 4576
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2222 4468 2228 4480
rect 2183 4440 2228 4468
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 2884 4477 2912 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 13078 4672 13084 4684
rect 12452 4644 13084 4672
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6972 4576 7113 4604
rect 6972 4564 6978 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9122 4604 9128 4616
rect 9079 4576 9128 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11112 4576 11345 4604
rect 11112 4564 11118 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 12452 4600 12480 4644
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 11333 4567 11391 4573
rect 12406 4572 12480 4600
rect 7650 4536 7656 4548
rect 5552 4508 7656 4536
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4437 2927 4471
rect 2869 4431 2927 4437
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 5552 4477 5580 4508
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8205 4539 8263 4545
rect 8205 4536 8217 4539
rect 7800 4508 8217 4536
rect 7800 4496 7806 4508
rect 8205 4505 8217 4508
rect 8251 4505 8263 4539
rect 8205 4499 8263 4505
rect 9309 4539 9367 4545
rect 9309 4505 9321 4539
rect 9355 4536 9367 4539
rect 12253 4539 12311 4545
rect 9355 4508 11192 4536
rect 9355 4505 9367 4508
rect 9309 4499 9367 4505
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 4028 4440 4353 4468
rect 4028 4428 4034 4440
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 4341 4431 4399 4437
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4437 5595 4471
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 5537 4431 5595 4437
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7282 4468 7288 4480
rect 7243 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 8444 4440 9137 4468
rect 8444 4428 8450 4440
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 10134 4468 10140 4480
rect 10095 4440 10140 4468
rect 9125 4431 9183 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 11164 4477 11192 4508
rect 12253 4505 12265 4539
rect 12299 4536 12311 4539
rect 12406 4536 12434 4572
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 12860 4576 13001 4604
rect 12860 4564 12866 4576
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 13354 4604 13360 4616
rect 13035 4576 13360 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13446 4564 13452 4616
rect 13504 4604 13510 4616
rect 14090 4604 14096 4616
rect 13504 4576 14096 4604
rect 13504 4564 13510 4576
rect 14090 4564 14096 4576
rect 14148 4604 14154 4616
rect 15764 4613 15792 4712
rect 26234 4700 26240 4712
rect 26292 4700 26298 4752
rect 22738 4672 22744 4684
rect 16592 4644 22744 4672
rect 16592 4613 16620 4644
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 25866 4632 25872 4684
rect 25924 4672 25930 4684
rect 25961 4675 26019 4681
rect 25961 4672 25973 4675
rect 25924 4644 25973 4672
rect 25924 4632 25930 4644
rect 25961 4641 25973 4644
rect 26007 4641 26019 4675
rect 25961 4635 26019 4641
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 14148 4576 14289 4604
rect 14148 4564 14154 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 16577 4567 16635 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 21508 4576 21557 4604
rect 21508 4564 21514 4576
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 22186 4604 22192 4616
rect 22147 4576 22192 4604
rect 21545 4567 21603 4573
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 25038 4564 25044 4616
rect 25096 4604 25102 4616
rect 26436 4613 26464 4780
rect 27430 4768 27436 4780
rect 27488 4768 27494 4820
rect 30561 4811 30619 4817
rect 30561 4777 30573 4811
rect 30607 4808 30619 4811
rect 31202 4808 31208 4820
rect 30607 4780 31208 4808
rect 30607 4777 30619 4780
rect 30561 4771 30619 4777
rect 31202 4768 31208 4780
rect 31260 4768 31266 4820
rect 32306 4808 32312 4820
rect 32267 4780 32312 4808
rect 32306 4768 32312 4780
rect 32364 4768 32370 4820
rect 33410 4808 33416 4820
rect 33371 4780 33416 4808
rect 33410 4768 33416 4780
rect 33468 4768 33474 4820
rect 33502 4768 33508 4820
rect 33560 4808 33566 4820
rect 35253 4811 35311 4817
rect 35253 4808 35265 4811
rect 33560 4780 35265 4808
rect 33560 4768 33566 4780
rect 35253 4777 35265 4780
rect 35299 4777 35311 4811
rect 35253 4771 35311 4777
rect 35986 4740 35992 4752
rect 26620 4712 35992 4740
rect 26620 4613 26648 4712
rect 35986 4700 35992 4712
rect 36044 4700 36050 4752
rect 36998 4700 37004 4752
rect 37056 4740 37062 4752
rect 37185 4743 37243 4749
rect 37185 4740 37197 4743
rect 37056 4712 37197 4740
rect 37056 4700 37062 4712
rect 37185 4709 37197 4712
rect 37231 4709 37243 4743
rect 37185 4703 37243 4709
rect 26878 4632 26884 4684
rect 26936 4672 26942 4684
rect 26936 4644 33272 4672
rect 26936 4632 26942 4644
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 25096 4576 25329 4604
rect 25096 4564 25102 4576
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 26421 4607 26479 4613
rect 26421 4573 26433 4607
rect 26467 4573 26479 4607
rect 26421 4567 26479 4573
rect 26605 4607 26663 4613
rect 26605 4573 26617 4607
rect 26651 4573 26663 4607
rect 26605 4567 26663 4573
rect 26694 4564 26700 4616
rect 26752 4604 26758 4616
rect 28626 4604 28632 4616
rect 26752 4576 26797 4604
rect 26896 4576 28632 4604
rect 26752 4564 26758 4576
rect 26896 4536 26924 4576
rect 28626 4564 28632 4576
rect 28684 4564 28690 4616
rect 30377 4607 30435 4613
rect 30377 4573 30389 4607
rect 30423 4573 30435 4607
rect 31018 4604 31024 4616
rect 30979 4576 31024 4604
rect 30377 4567 30435 4573
rect 12299 4508 12434 4536
rect 22066 4508 26924 4536
rect 12299 4505 12311 4508
rect 12253 4499 12311 4505
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 12805 4471 12863 4477
rect 12805 4468 12817 4471
rect 11296 4440 12817 4468
rect 11296 4428 11302 4440
rect 12805 4437 12817 4440
rect 12851 4437 12863 4471
rect 12805 4431 12863 4437
rect 13354 4428 13360 4480
rect 13412 4468 13418 4480
rect 13449 4471 13507 4477
rect 13449 4468 13461 4471
rect 13412 4440 13461 4468
rect 13412 4428 13418 4440
rect 13449 4437 13461 4440
rect 13495 4437 13507 4471
rect 14918 4468 14924 4480
rect 14879 4440 14924 4468
rect 13449 4431 13507 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 15528 4440 15577 4468
rect 15528 4428 15534 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 15565 4431 15623 4437
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16264 4440 16405 4468
rect 16264 4428 16270 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 17034 4468 17040 4480
rect 16995 4440 17040 4468
rect 16393 4431 16451 4437
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 17586 4468 17592 4480
rect 17547 4440 17592 4468
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 18141 4471 18199 4477
rect 18141 4468 18153 4471
rect 18104 4440 18153 4468
rect 18104 4428 18110 4440
rect 18141 4437 18153 4440
rect 18187 4437 18199 4471
rect 18141 4431 18199 4437
rect 19613 4471 19671 4477
rect 19613 4437 19625 4471
rect 19659 4468 19671 4471
rect 20162 4468 20168 4480
rect 19659 4440 20168 4468
rect 19659 4437 19671 4440
rect 19613 4431 19671 4437
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 20530 4468 20536 4480
rect 20303 4440 20536 4468
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21542 4468 21548 4480
rect 21131 4440 21548 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 21729 4471 21787 4477
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 22066 4468 22094 4508
rect 27338 4496 27344 4548
rect 27396 4536 27402 4548
rect 27985 4539 28043 4545
rect 27985 4536 27997 4539
rect 27396 4508 27997 4536
rect 27396 4496 27402 4508
rect 27985 4505 27997 4508
rect 28031 4505 28043 4539
rect 30392 4536 30420 4567
rect 31018 4564 31024 4576
rect 31076 4564 31082 4616
rect 31110 4564 31116 4616
rect 31168 4604 31174 4616
rect 33244 4613 33272 4644
rect 32125 4607 32183 4613
rect 32125 4604 32137 4607
rect 31168 4576 32137 4604
rect 31168 4564 31174 4576
rect 32125 4573 32137 4576
rect 32171 4573 32183 4607
rect 32125 4567 32183 4573
rect 33229 4607 33287 4613
rect 33229 4573 33241 4607
rect 33275 4573 33287 4607
rect 33229 4567 33287 4573
rect 33686 4564 33692 4616
rect 33744 4604 33750 4616
rect 33965 4607 34023 4613
rect 33965 4604 33977 4607
rect 33744 4576 33977 4604
rect 33744 4564 33750 4576
rect 33965 4573 33977 4576
rect 34011 4573 34023 4607
rect 36078 4604 36084 4616
rect 36039 4576 36084 4604
rect 33965 4567 34023 4573
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 37182 4564 37188 4616
rect 37240 4604 37246 4616
rect 38105 4607 38163 4613
rect 38105 4604 38117 4607
rect 37240 4576 38117 4604
rect 37240 4564 37246 4576
rect 38105 4573 38117 4576
rect 38151 4573 38163 4607
rect 38105 4567 38163 4573
rect 30558 4536 30564 4548
rect 30392 4508 30564 4536
rect 27985 4499 28043 4505
rect 30558 4496 30564 4508
rect 30616 4536 30622 4548
rect 31570 4536 31576 4548
rect 30616 4508 31576 4536
rect 30616 4496 30622 4508
rect 31570 4496 31576 4508
rect 31628 4496 31634 4548
rect 35158 4536 35164 4548
rect 35119 4508 35164 4536
rect 35158 4496 35164 4508
rect 35216 4496 35222 4548
rect 37366 4536 37372 4548
rect 37279 4508 37372 4536
rect 37366 4496 37372 4508
rect 37424 4536 37430 4548
rect 37918 4536 37924 4548
rect 37424 4508 37924 4536
rect 37424 4496 37430 4508
rect 37918 4496 37924 4508
rect 37976 4496 37982 4548
rect 22370 4468 22376 4480
rect 21775 4440 22094 4468
rect 22331 4440 22376 4468
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 22370 4428 22376 4440
rect 22428 4428 22434 4480
rect 22925 4471 22983 4477
rect 22925 4437 22937 4471
rect 22971 4468 22983 4471
rect 23014 4468 23020 4480
rect 22971 4440 23020 4468
rect 22971 4437 22983 4440
rect 22925 4431 22983 4437
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 23842 4468 23848 4480
rect 23803 4440 23848 4468
rect 23842 4428 23848 4440
rect 23900 4428 23906 4480
rect 24670 4468 24676 4480
rect 24631 4440 24676 4468
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 28258 4428 28264 4480
rect 28316 4468 28322 4480
rect 28537 4471 28595 4477
rect 28537 4468 28549 4471
rect 28316 4440 28549 4468
rect 28316 4428 28322 4440
rect 28537 4437 28549 4440
rect 28583 4437 28595 4471
rect 28537 4431 28595 4437
rect 29270 4428 29276 4480
rect 29328 4468 29334 4480
rect 29549 4471 29607 4477
rect 29549 4468 29561 4471
rect 29328 4440 29561 4468
rect 29328 4428 29334 4440
rect 29549 4437 29561 4440
rect 29595 4437 29607 4471
rect 29549 4431 29607 4437
rect 30374 4428 30380 4480
rect 30432 4468 30438 4480
rect 31205 4471 31263 4477
rect 31205 4468 31217 4471
rect 30432 4440 31217 4468
rect 30432 4428 30438 4440
rect 31205 4437 31217 4440
rect 31251 4437 31263 4471
rect 31205 4431 31263 4437
rect 31478 4428 31484 4480
rect 31536 4468 31542 4480
rect 33778 4468 33784 4480
rect 31536 4440 33784 4468
rect 31536 4428 31542 4440
rect 33778 4428 33784 4440
rect 33836 4428 33842 4480
rect 34146 4468 34152 4480
rect 34107 4440 34152 4468
rect 34146 4428 34152 4440
rect 34204 4428 34210 4480
rect 35986 4428 35992 4480
rect 36044 4468 36050 4480
rect 36265 4471 36323 4477
rect 36265 4468 36277 4471
rect 36044 4440 36277 4468
rect 36044 4428 36050 4440
rect 36265 4437 36277 4440
rect 36311 4437 36323 4471
rect 36265 4431 36323 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2777 4267 2835 4273
rect 2777 4233 2789 4267
rect 2823 4264 2835 4267
rect 3878 4264 3884 4276
rect 2823 4236 3884 4264
rect 2823 4233 2835 4236
rect 2777 4227 2835 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4433 4267 4491 4273
rect 4433 4233 4445 4267
rect 4479 4264 4491 4267
rect 5534 4264 5540 4276
rect 4479 4236 5540 4264
rect 4479 4233 4491 4236
rect 4433 4227 4491 4233
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 7340 4236 19257 4264
rect 7340 4224 7346 4236
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 20530 4264 20536 4276
rect 20491 4236 20536 4264
rect 19245 4227 19303 4233
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4264 20959 4267
rect 21634 4264 21640 4276
rect 20947 4236 21640 4264
rect 20947 4233 20959 4236
rect 20901 4227 20959 4233
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 22278 4224 22284 4276
rect 22336 4264 22342 4276
rect 24489 4267 24547 4273
rect 24489 4264 24501 4267
rect 22336 4236 24501 4264
rect 22336 4224 22342 4236
rect 24489 4233 24501 4236
rect 24535 4264 24547 4267
rect 24670 4264 24676 4276
rect 24535 4236 24676 4264
rect 24535 4233 24547 4236
rect 24489 4227 24547 4233
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 28994 4224 29000 4276
rect 29052 4264 29058 4276
rect 32398 4264 32404 4276
rect 29052 4236 32404 4264
rect 29052 4224 29058 4236
rect 32398 4224 32404 4236
rect 32456 4224 32462 4276
rect 4798 4156 4804 4208
rect 4856 4156 4862 4208
rect 5368 4168 5672 4196
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 624 4100 1409 4128
rect 624 4088 630 4100
rect 1397 4097 1409 4100
rect 1443 4128 1455 4131
rect 1946 4128 1952 4140
rect 1443 4100 1952 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 2924 4100 2969 4128
rect 2924 4088 2930 4100
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 3200 4100 3617 4128
rect 3200 4088 3206 4100
rect 3605 4097 3617 4100
rect 3651 4128 3663 4131
rect 4062 4128 4068 4140
rect 3651 4100 4068 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4816 4128 4844 4156
rect 4295 4100 4844 4128
rect 4893 4131 4951 4137
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4893 4097 4905 4131
rect 4939 4128 4951 4131
rect 4982 4128 4988 4140
rect 4939 4100 4988 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 290 4020 296 4072
rect 348 4060 354 4072
rect 1578 4060 1584 4072
rect 348 4032 1584 4060
rect 348 4020 354 4032
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 3050 4060 3056 4072
rect 3011 4032 3056 4060
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 4264 4060 4292 4091
rect 4982 4088 4988 4100
rect 5040 4128 5046 4140
rect 5368 4128 5396 4168
rect 5040 4100 5396 4128
rect 5040 4088 5046 4100
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5500 4100 5549 4128
rect 5500 4088 5506 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5644 4128 5672 4168
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 7469 4199 7527 4205
rect 7469 4196 7481 4199
rect 7248 4168 7481 4196
rect 7248 4156 7254 4168
rect 7469 4165 7481 4168
rect 7515 4165 7527 4199
rect 7469 4159 7527 4165
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 10137 4199 10195 4205
rect 10137 4196 10149 4199
rect 7708 4168 10149 4196
rect 7708 4156 7714 4168
rect 10137 4165 10149 4168
rect 10183 4165 10195 4199
rect 19794 4196 19800 4208
rect 10137 4159 10195 4165
rect 14660 4168 14872 4196
rect 5718 4128 5724 4140
rect 5644 4100 5724 4128
rect 5537 4091 5595 4097
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 6420 4100 6469 4128
rect 6420 4088 6426 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8628 4100 8677 4128
rect 8628 4088 8634 4100
rect 8665 4097 8677 4100
rect 8711 4128 8723 4131
rect 9030 4128 9036 4140
rect 8711 4100 9036 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 11882 4128 11888 4140
rect 10152 4100 10364 4128
rect 11843 4100 11888 4128
rect 3620 4032 4292 4060
rect 3620 4004 3648 4032
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5460 4060 5488 4088
rect 8386 4060 8392 4072
rect 4856 4032 5488 4060
rect 5736 4032 8392 4060
rect 4856 4020 4862 4032
rect 2406 3992 2412 4004
rect 2367 3964 2412 3992
rect 2406 3952 2412 3964
rect 2464 3952 2470 4004
rect 3602 3952 3608 4004
rect 3660 3952 3666 4004
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 5074 3992 5080 4004
rect 3835 3964 4936 3992
rect 5035 3964 5080 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2866 3924 2872 3936
rect 1627 3896 2872 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 4908 3924 4936 3964
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5442 3992 5448 4004
rect 5224 3964 5448 3992
rect 5224 3952 5230 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5736 4001 5764 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8938 4060 8944 4072
rect 8899 4032 8944 4060
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 9916 4032 10057 4060
rect 9916 4020 9922 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 5721 3995 5779 4001
rect 5721 3961 5733 3995
rect 5767 3961 5779 3995
rect 7558 3992 7564 4004
rect 5721 3955 5779 3961
rect 6564 3964 7564 3992
rect 6564 3924 6592 3964
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 7653 3995 7711 4001
rect 7653 3961 7665 3995
rect 7699 3992 7711 3995
rect 10152 3992 10180 4100
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4029 10287 4063
rect 10336 4060 10364 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12526 4128 12532 4140
rect 12032 4100 12532 4128
rect 12032 4088 12038 4100
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13722 4128 13728 4140
rect 13683 4100 13728 4128
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14660 4060 14688 4168
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14844 4128 14872 4168
rect 15396 4168 16252 4196
rect 15396 4128 15424 4168
rect 14844 4100 15424 4128
rect 15473 4131 15531 4137
rect 14737 4091 14795 4097
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 16114 4128 16120 4140
rect 15519 4100 16120 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 10336 4032 14688 4060
rect 14752 4060 14780 4091
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 16224 4128 16252 4168
rect 17328 4168 19800 4196
rect 17328 4128 17356 4168
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 31110 4196 31116 4208
rect 20916 4168 31116 4196
rect 16224 4100 17356 4128
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4128 17463 4131
rect 19150 4128 19156 4140
rect 17451 4100 19156 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 19334 4128 19340 4140
rect 19295 4100 19340 4128
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 20916 4128 20944 4168
rect 31110 4156 31116 4168
rect 31168 4156 31174 4208
rect 31864 4168 32076 4196
rect 19720 4100 20944 4128
rect 15562 4060 15568 4072
rect 14752 4032 15568 4060
rect 10229 4023 10287 4029
rect 7699 3964 10180 3992
rect 10244 3992 10272 4023
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 17770 4060 17776 4072
rect 17092 4032 17776 4060
rect 17092 4020 17098 4032
rect 12345 3995 12403 4001
rect 12345 3992 12357 3995
rect 10244 3964 12357 3992
rect 7699 3961 7711 3964
rect 7653 3955 7711 3961
rect 12345 3961 12357 3964
rect 12391 3961 12403 3995
rect 12345 3955 12403 3961
rect 12986 3952 12992 4004
rect 13044 3992 13050 4004
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 13044 3964 13921 3992
rect 13044 3952 13050 3964
rect 13909 3961 13921 3964
rect 13955 3961 13967 3995
rect 13909 3955 13967 3961
rect 14090 3952 14096 4004
rect 14148 3992 14154 4004
rect 17236 3992 17264 4032
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 19058 4060 19064 4072
rect 19019 4032 19064 4060
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 14148 3964 17264 3992
rect 14148 3952 14154 3964
rect 17310 3952 17316 4004
rect 17368 3992 17374 4004
rect 19720 4001 19748 4100
rect 21726 4088 21732 4140
rect 21784 4128 21790 4140
rect 22186 4128 22192 4140
rect 21784 4100 22192 4128
rect 21784 4088 21790 4100
rect 22186 4088 22192 4100
rect 22244 4088 22250 4140
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 22373 4091 22431 4097
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19852 4032 20269 4060
rect 19852 4020 19858 4032
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20257 4023 20315 4029
rect 17957 3995 18015 4001
rect 17957 3992 17969 3995
rect 17368 3964 17969 3992
rect 17368 3952 17374 3964
rect 17957 3961 17969 3964
rect 18003 3992 18015 3995
rect 19705 3995 19763 4001
rect 18003 3964 19104 3992
rect 18003 3961 18015 3964
rect 17957 3955 18015 3961
rect 4908 3896 6592 3924
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 7006 3924 7012 3936
rect 6687 3896 7012 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 10778 3924 10784 3936
rect 10643 3896 10784 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11480 3896 11713 3924
rect 11480 3884 11486 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12216 3896 13185 3924
rect 12216 3884 12222 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 13173 3887 13231 3893
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 13780 3896 14565 3924
rect 13780 3884 13786 3896
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14553 3887 14611 3893
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 14792 3896 15301 3924
rect 14792 3884 14798 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 15289 3887 15347 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 17092 3896 17233 3924
rect 17092 3884 17098 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18196 3896 18429 3924
rect 18196 3884 18202 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 19076 3924 19104 3964
rect 19705 3961 19717 3995
rect 19751 3961 19763 3995
rect 20272 3992 20300 4023
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 20404 4032 20453 4060
rect 20404 4020 20410 4032
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 22388 4060 22416 4091
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 24029 4131 24087 4137
rect 24029 4097 24041 4131
rect 24075 4128 24087 4131
rect 24762 4128 24768 4140
rect 24075 4100 24768 4128
rect 24075 4097 24087 4100
rect 24029 4091 24087 4097
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 25225 4131 25283 4137
rect 25225 4097 25237 4131
rect 25271 4128 25283 4131
rect 27157 4131 27215 4137
rect 27157 4128 27169 4131
rect 25271 4100 26188 4128
rect 25271 4097 25283 4100
rect 25225 4091 25283 4097
rect 25590 4060 25596 4072
rect 22388 4032 25596 4060
rect 20441 4023 20499 4029
rect 25590 4020 25596 4032
rect 25648 4020 25654 4072
rect 26160 4069 26188 4100
rect 26620 4100 27169 4128
rect 25685 4063 25743 4069
rect 25685 4029 25697 4063
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 26145 4063 26203 4069
rect 26145 4029 26157 4063
rect 26191 4029 26203 4063
rect 26145 4023 26203 4029
rect 20622 3992 20628 4004
rect 20272 3964 20628 3992
rect 19705 3955 19763 3961
rect 20622 3952 20628 3964
rect 20680 3952 20686 4004
rect 22922 3952 22928 4004
rect 22980 3992 22986 4004
rect 25041 3995 25099 4001
rect 25041 3992 25053 3995
rect 22980 3964 25053 3992
rect 22980 3952 22986 3964
rect 25041 3961 25053 3964
rect 25087 3961 25099 3995
rect 25700 3992 25728 4023
rect 26050 3992 26056 4004
rect 25041 3955 25099 3961
rect 25608 3964 25728 3992
rect 26011 3964 26056 3992
rect 20530 3924 20536 3936
rect 19076 3896 20536 3924
rect 18417 3887 18475 3893
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22189 3927 22247 3933
rect 22189 3924 22201 3927
rect 22060 3896 22201 3924
rect 22060 3884 22066 3896
rect 22189 3893 22201 3896
rect 22235 3893 22247 3927
rect 22189 3887 22247 3893
rect 22830 3884 22836 3936
rect 22888 3924 22894 3936
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22888 3896 23029 3924
rect 22888 3884 22894 3896
rect 23017 3893 23029 3896
rect 23063 3893 23075 3927
rect 23017 3887 23075 3893
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 23716 3896 23857 3924
rect 23716 3884 23722 3896
rect 23845 3893 23857 3896
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 24670 3884 24676 3936
rect 24728 3924 24734 3936
rect 25314 3924 25320 3936
rect 24728 3896 25320 3924
rect 24728 3884 24734 3896
rect 25314 3884 25320 3896
rect 25372 3924 25378 3936
rect 25608 3924 25636 3964
rect 26050 3952 26056 3964
rect 26108 3952 26114 4004
rect 25372 3896 25636 3924
rect 25372 3884 25378 3896
rect 25682 3884 25688 3936
rect 25740 3924 25746 3936
rect 26620 3924 26648 4100
rect 27157 4097 27169 4100
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27522 4088 27528 4140
rect 27580 4128 27586 4140
rect 27801 4131 27859 4137
rect 27801 4128 27813 4131
rect 27580 4100 27813 4128
rect 27580 4088 27586 4100
rect 27801 4097 27813 4100
rect 27847 4097 27859 4131
rect 27801 4091 27859 4097
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 28629 4131 28687 4137
rect 28629 4128 28641 4131
rect 28224 4100 28641 4128
rect 28224 4088 28230 4100
rect 28629 4097 28641 4100
rect 28675 4097 28687 4131
rect 28629 4091 28687 4097
rect 28810 4088 28816 4140
rect 28868 4128 28874 4140
rect 30282 4128 30288 4140
rect 28868 4100 29960 4128
rect 30243 4100 30288 4128
rect 28868 4088 28874 4100
rect 28074 4020 28080 4072
rect 28132 4060 28138 4072
rect 28132 4032 29224 4060
rect 28132 4020 28138 4032
rect 29196 4004 29224 4032
rect 29270 4020 29276 4072
rect 29328 4060 29334 4072
rect 29825 4063 29883 4069
rect 29825 4060 29837 4063
rect 29328 4032 29837 4060
rect 29328 4020 29334 4032
rect 29825 4029 29837 4032
rect 29871 4029 29883 4063
rect 29932 4060 29960 4100
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 30469 4131 30527 4137
rect 30469 4097 30481 4131
rect 30515 4128 30527 4131
rect 30558 4128 30564 4140
rect 30515 4100 30564 4128
rect 30515 4097 30527 4100
rect 30469 4091 30527 4097
rect 30558 4088 30564 4100
rect 30616 4088 30622 4140
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 31021 4131 31079 4137
rect 31021 4128 31033 4131
rect 30800 4100 31033 4128
rect 30800 4088 30806 4100
rect 31021 4097 31033 4100
rect 31067 4097 31079 4131
rect 31021 4091 31079 4097
rect 31864 4060 31892 4168
rect 29932 4032 31892 4060
rect 32048 4060 32076 4168
rect 32214 4156 32220 4208
rect 32272 4196 32278 4208
rect 32766 4196 32772 4208
rect 32272 4168 32772 4196
rect 32272 4156 32278 4168
rect 32766 4156 32772 4168
rect 32824 4156 32830 4208
rect 36262 4156 36268 4208
rect 36320 4196 36326 4208
rect 36541 4199 36599 4205
rect 36541 4196 36553 4199
rect 36320 4168 36553 4196
rect 36320 4156 36326 4168
rect 36541 4165 36553 4168
rect 36587 4165 36599 4199
rect 36541 4159 36599 4165
rect 32122 4088 32128 4140
rect 32180 4128 32186 4140
rect 32180 4100 32225 4128
rect 32180 4088 32186 4100
rect 32306 4088 32312 4140
rect 32364 4128 32370 4140
rect 32861 4131 32919 4137
rect 32861 4128 32873 4131
rect 32364 4100 32873 4128
rect 32364 4088 32370 4100
rect 32861 4097 32873 4100
rect 32907 4097 32919 4131
rect 32861 4091 32919 4097
rect 33965 4131 34023 4137
rect 33965 4097 33977 4131
rect 34011 4097 34023 4131
rect 33965 4091 34023 4097
rect 33980 4060 34008 4091
rect 34146 4088 34152 4140
rect 34204 4128 34210 4140
rect 35253 4131 35311 4137
rect 35253 4128 35265 4131
rect 34204 4100 35265 4128
rect 34204 4088 34210 4100
rect 35253 4097 35265 4100
rect 35299 4097 35311 4131
rect 35253 4091 35311 4097
rect 35526 4088 35532 4140
rect 35584 4128 35590 4140
rect 36357 4131 36415 4137
rect 36357 4128 36369 4131
rect 35584 4100 36369 4128
rect 35584 4088 35590 4100
rect 36357 4097 36369 4100
rect 36403 4097 36415 4131
rect 36357 4091 36415 4097
rect 37277 4131 37335 4137
rect 37277 4097 37289 4131
rect 37323 4097 37335 4131
rect 37277 4091 37335 4097
rect 38105 4131 38163 4137
rect 38105 4097 38117 4131
rect 38151 4128 38163 4131
rect 38378 4128 38384 4140
rect 38151 4100 38384 4128
rect 38151 4097 38163 4100
rect 38105 4091 38163 4097
rect 32048 4032 34008 4060
rect 29825 4023 29883 4029
rect 34422 4020 34428 4072
rect 34480 4060 34486 4072
rect 37292 4060 37320 4091
rect 38378 4088 38384 4100
rect 38436 4088 38442 4140
rect 34480 4032 37320 4060
rect 34480 4020 34486 4032
rect 26694 3952 26700 4004
rect 26752 3992 26758 4004
rect 27617 3995 27675 4001
rect 27617 3992 27629 3995
rect 26752 3964 27629 3992
rect 26752 3952 26758 3964
rect 27617 3961 27629 3964
rect 27663 3961 27675 3995
rect 27617 3955 27675 3961
rect 28166 3952 28172 4004
rect 28224 3992 28230 4004
rect 28350 3992 28356 4004
rect 28224 3964 28356 3992
rect 28224 3952 28230 3964
rect 28350 3952 28356 3964
rect 28408 3952 28414 4004
rect 29178 3992 29184 4004
rect 29091 3964 29184 3992
rect 29178 3952 29184 3964
rect 29236 3992 29242 4004
rect 29457 3995 29515 4001
rect 29457 3992 29469 3995
rect 29236 3964 29469 3992
rect 29236 3952 29242 3964
rect 29457 3961 29469 3964
rect 29503 3961 29515 3995
rect 29457 3955 29515 3961
rect 29546 3952 29552 4004
rect 29604 3992 29610 4004
rect 32214 3992 32220 4004
rect 29604 3964 32220 3992
rect 29604 3952 29610 3964
rect 32214 3952 32220 3964
rect 32272 3952 32278 4004
rect 32398 3952 32404 4004
rect 32456 3992 32462 4004
rect 34149 3995 34207 4001
rect 34149 3992 34161 3995
rect 32456 3964 34161 3992
rect 32456 3952 32462 3964
rect 34149 3961 34161 3964
rect 34195 3961 34207 3995
rect 34149 3955 34207 3961
rect 34330 3952 34336 4004
rect 34388 3992 34394 4004
rect 35618 3992 35624 4004
rect 34388 3964 35624 3992
rect 34388 3952 34394 3964
rect 35618 3952 35624 3964
rect 35676 3952 35682 4004
rect 37090 3952 37096 4004
rect 37148 3992 37154 4004
rect 37366 3992 37372 4004
rect 37148 3964 37372 3992
rect 37148 3952 37154 3964
rect 37366 3952 37372 3964
rect 37424 3952 37430 4004
rect 37461 3995 37519 4001
rect 37461 3961 37473 3995
rect 37507 3992 37519 3995
rect 38194 3992 38200 4004
rect 37507 3964 38200 3992
rect 37507 3961 37519 3964
rect 37461 3955 37519 3961
rect 38194 3952 38200 3964
rect 38252 3952 38258 4004
rect 26970 3924 26976 3936
rect 25740 3896 26648 3924
rect 26931 3896 26976 3924
rect 25740 3884 25746 3896
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 28534 3884 28540 3936
rect 28592 3924 28598 3936
rect 28813 3927 28871 3933
rect 28813 3924 28825 3927
rect 28592 3896 28825 3924
rect 28592 3884 28598 3896
rect 28813 3893 28825 3896
rect 28859 3893 28871 3927
rect 28813 3887 28871 3893
rect 28994 3884 29000 3936
rect 29052 3924 29058 3936
rect 29365 3927 29423 3933
rect 29365 3924 29377 3927
rect 29052 3896 29377 3924
rect 29052 3884 29058 3896
rect 29365 3893 29377 3896
rect 29411 3893 29423 3927
rect 29365 3887 29423 3893
rect 29822 3884 29828 3936
rect 29880 3924 29886 3936
rect 31205 3927 31263 3933
rect 31205 3924 31217 3927
rect 29880 3896 31217 3924
rect 29880 3884 29886 3896
rect 31205 3893 31217 3896
rect 31251 3893 31263 3927
rect 31205 3887 31263 3893
rect 31846 3884 31852 3936
rect 31904 3924 31910 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 31904 3896 32321 3924
rect 31904 3884 31910 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 32309 3887 32367 3893
rect 33045 3927 33103 3933
rect 33045 3893 33057 3927
rect 33091 3924 33103 3927
rect 33778 3924 33784 3936
rect 33091 3896 33784 3924
rect 33091 3893 33103 3896
rect 33045 3887 33103 3893
rect 33778 3884 33784 3896
rect 33836 3884 33842 3936
rect 34238 3884 34244 3936
rect 34296 3924 34302 3936
rect 34701 3927 34759 3933
rect 34701 3924 34713 3927
rect 34296 3896 34713 3924
rect 34296 3884 34302 3896
rect 34701 3893 34713 3896
rect 34747 3893 34759 3927
rect 34701 3887 34759 3893
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 35437 3927 35495 3933
rect 35437 3924 35449 3927
rect 35400 3896 35449 3924
rect 35400 3884 35406 3896
rect 35437 3893 35449 3896
rect 35483 3893 35495 3927
rect 35437 3887 35495 3893
rect 36722 3884 36728 3936
rect 36780 3924 36786 3936
rect 39022 3924 39028 3936
rect 36780 3896 39028 3924
rect 36780 3884 36786 3896
rect 39022 3884 39028 3896
rect 39080 3884 39086 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4948 3692 4997 3720
rect 4948 3680 4954 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 4985 3683 5043 3689
rect 5184 3692 5764 3720
rect 5184 3652 5212 3692
rect 2056 3624 5212 3652
rect 2056 3593 2084 3624
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2280 3556 5120 3584
rect 2280 3544 2286 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1728 3488 1777 3516
rect 1728 3476 1734 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 3234 3516 3240 3528
rect 1765 3479 1823 3485
rect 1872 3488 3240 3516
rect 842 3408 848 3460
rect 900 3448 906 3460
rect 1872 3448 1900 3488
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3752 3488 3801 3516
rect 3752 3476 3758 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4982 3516 4988 3528
rect 4212 3488 4988 3516
rect 4212 3476 4218 3488
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5092 3516 5120 3556
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5537 3587 5595 3593
rect 5537 3584 5549 3587
rect 5500 3556 5549 3584
rect 5500 3544 5506 3556
rect 5537 3553 5549 3556
rect 5583 3553 5595 3587
rect 5736 3584 5764 3692
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 6052 3692 6193 3720
rect 6052 3680 6058 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 11606 3720 11612 3732
rect 11563 3692 11612 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 12124 3692 13185 3720
rect 12124 3680 12130 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 14458 3720 14464 3732
rect 14139 3692 14464 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 16485 3723 16543 3729
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 17126 3720 17132 3732
rect 16531 3692 17132 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 19334 3720 19340 3732
rect 19295 3692 19340 3720
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 19794 3680 19800 3732
rect 19852 3720 19858 3732
rect 19981 3723 20039 3729
rect 19981 3720 19993 3723
rect 19852 3692 19993 3720
rect 19852 3680 19858 3692
rect 19981 3689 19993 3692
rect 20027 3689 20039 3723
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 19981 3683 20039 3689
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 21361 3723 21419 3729
rect 21361 3689 21373 3723
rect 21407 3720 21419 3723
rect 25593 3723 25651 3729
rect 21407 3692 25268 3720
rect 21407 3689 21419 3692
rect 21361 3683 21419 3689
rect 7745 3655 7803 3661
rect 7745 3621 7757 3655
rect 7791 3652 7803 3655
rect 7926 3652 7932 3664
rect 7791 3624 7932 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8389 3655 8447 3661
rect 8389 3621 8401 3655
rect 8435 3652 8447 3655
rect 20346 3652 20352 3664
rect 8435 3624 20352 3652
rect 8435 3621 8447 3624
rect 8389 3615 8447 3621
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 22554 3652 22560 3664
rect 22515 3624 22560 3652
rect 22554 3612 22560 3624
rect 22612 3612 22618 3664
rect 24486 3612 24492 3664
rect 24544 3652 24550 3664
rect 24765 3655 24823 3661
rect 24765 3652 24777 3655
rect 24544 3624 24777 3652
rect 24544 3612 24550 3624
rect 24765 3621 24777 3624
rect 24811 3621 24823 3655
rect 24765 3615 24823 3621
rect 6546 3584 6552 3596
rect 5736 3556 6552 3584
rect 5537 3547 5595 3553
rect 6546 3544 6552 3556
rect 6604 3584 6610 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 6604 3556 6745 3584
rect 6604 3544 6610 3556
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 6840 3556 8616 3584
rect 5092 3512 5212 3516
rect 5276 3512 5488 3516
rect 5092 3488 5488 3512
rect 5184 3484 5304 3488
rect 900 3420 1900 3448
rect 900 3408 906 3420
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 3712 3448 3740 3476
rect 2004 3420 3740 3448
rect 2004 3408 2010 3420
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 3016 3352 3065 3380
rect 3016 3340 3022 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4430 3380 4436 3392
rect 4019 3352 4436 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4525 3383 4583 3389
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 4890 3380 4896 3392
rect 4571 3352 4896 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 5460 3389 5488 3488
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6840 3516 6868 3556
rect 5776 3488 6868 3516
rect 5776 3476 5782 3488
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7524 3488 8217 3516
rect 7524 3476 7530 3488
rect 8205 3485 8217 3488
rect 8251 3516 8263 3519
rect 8478 3516 8484 3528
rect 8251 3488 8484 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8588 3516 8616 3556
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 9456 3556 9505 3584
rect 9456 3544 9462 3556
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 12529 3587 12587 3593
rect 9493 3547 9551 3553
rect 9600 3556 12434 3584
rect 9600 3516 9628 3556
rect 8588 3488 9628 3516
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 10870 3516 10876 3528
rect 9815 3488 10876 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11238 3516 11244 3528
rect 11199 3488 11244 3516
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 6270 3408 6276 3460
rect 6328 3448 6334 3460
rect 6641 3451 6699 3457
rect 6641 3448 6653 3451
rect 6328 3420 6653 3448
rect 6328 3408 6334 3420
rect 6641 3417 6653 3420
rect 6687 3417 6699 3451
rect 6641 3411 6699 3417
rect 6730 3408 6736 3460
rect 6788 3448 6794 3460
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 6788 3420 7573 3448
rect 6788 3408 6794 3420
rect 7561 3417 7573 3420
rect 7607 3448 7619 3451
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 7607 3420 8953 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 8941 3417 8953 3420
rect 8987 3417 8999 3451
rect 10965 3451 11023 3457
rect 10965 3448 10977 3451
rect 8941 3411 8999 3417
rect 9048 3420 10977 3448
rect 5353 3383 5411 3389
rect 5353 3380 5365 3383
rect 5316 3352 5365 3380
rect 5316 3340 5322 3352
rect 5353 3349 5365 3352
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 5445 3383 5503 3389
rect 5445 3349 5457 3383
rect 5491 3349 5503 3383
rect 5445 3343 5503 3349
rect 6549 3383 6607 3389
rect 6549 3349 6561 3383
rect 6595 3380 6607 3383
rect 7006 3380 7012 3392
rect 6595 3352 7012 3380
rect 6595 3349 6607 3352
rect 6549 3343 6607 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 9048 3380 9076 3420
rect 10965 3417 10977 3420
rect 11011 3448 11023 3451
rect 11146 3448 11152 3460
rect 11011 3420 11152 3448
rect 11011 3417 11023 3420
rect 10965 3411 11023 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 12406 3448 12434 3556
rect 12529 3553 12541 3587
rect 12575 3553 12587 3587
rect 12710 3584 12716 3596
rect 12671 3556 12716 3584
rect 12529 3547 12587 3553
rect 12544 3516 12572 3547
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 14182 3544 14188 3596
rect 14240 3584 14246 3596
rect 14645 3587 14703 3593
rect 14645 3584 14657 3587
rect 14240 3556 14657 3584
rect 14240 3544 14246 3556
rect 14645 3553 14657 3556
rect 14691 3553 14703 3587
rect 15838 3584 15844 3596
rect 14645 3547 14703 3553
rect 15396 3556 15844 3584
rect 13078 3516 13084 3528
rect 12544 3488 13084 3516
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 14090 3476 14096 3528
rect 14148 3476 14154 3528
rect 14458 3516 14464 3528
rect 14371 3488 14464 3516
rect 14458 3476 14464 3488
rect 14516 3516 14522 3528
rect 14918 3516 14924 3528
rect 14516 3488 14924 3516
rect 14516 3476 14522 3488
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 14108 3448 14136 3476
rect 14550 3448 14556 3460
rect 12406 3420 14136 3448
rect 14511 3420 14556 3448
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 7984 3352 9076 3380
rect 7984 3340 7990 3352
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 9364 3352 11069 3380
rect 9364 3340 9370 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11057 3343 11115 3349
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 13630 3380 13636 3392
rect 12851 3352 13636 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 15396 3380 15424 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 17589 3587 17647 3593
rect 16540 3556 17448 3584
rect 16540 3544 16546 3556
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 17310 3516 17316 3528
rect 17271 3488 17316 3516
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17420 3516 17448 3556
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 17770 3584 17776 3596
rect 17635 3556 17776 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 22005 3587 22063 3593
rect 22005 3553 22017 3587
rect 22051 3584 22063 3587
rect 22278 3584 22284 3596
rect 22051 3556 22284 3584
rect 22051 3553 22063 3556
rect 22005 3547 22063 3553
rect 22278 3544 22284 3556
rect 22336 3544 22342 3596
rect 23014 3544 23020 3596
rect 23072 3584 23078 3596
rect 23109 3587 23167 3593
rect 23109 3584 23121 3587
rect 23072 3556 23121 3584
rect 23072 3544 23078 3556
rect 23109 3553 23121 3556
rect 23155 3584 23167 3587
rect 23155 3556 25176 3584
rect 23155 3553 23167 3556
rect 23109 3547 23167 3553
rect 18417 3519 18475 3525
rect 17420 3488 17816 3516
rect 17678 3448 17684 3460
rect 17236 3420 17684 3448
rect 16022 3380 16028 3392
rect 14148 3352 15424 3380
rect 15983 3352 16028 3380
rect 14148 3340 14154 3352
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 16945 3383 17003 3389
rect 16945 3349 16957 3383
rect 16991 3380 17003 3383
rect 17236 3380 17264 3420
rect 17678 3408 17684 3420
rect 17736 3408 17742 3460
rect 17788 3448 17816 3488
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18506 3516 18512 3528
rect 18463 3488 18512 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19242 3516 19248 3528
rect 19024 3488 19248 3516
rect 19024 3476 19030 3488
rect 19242 3476 19248 3488
rect 19300 3516 19306 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19300 3488 19533 3516
rect 19300 3476 19306 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 20438 3476 20444 3528
rect 20496 3516 20502 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20496 3488 20545 3516
rect 20496 3476 20502 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21174 3516 21180 3528
rect 20680 3488 21180 3516
rect 20680 3476 20686 3488
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 21542 3476 21548 3528
rect 21600 3516 21606 3528
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 21600 3488 22201 3516
rect 21600 3476 21606 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 22370 3476 22376 3528
rect 22428 3516 22434 3528
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 22428 3488 23397 3516
rect 22428 3476 22434 3488
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 24210 3516 24216 3528
rect 23808 3488 24216 3516
rect 23808 3476 23814 3488
rect 24210 3476 24216 3488
rect 24268 3516 24274 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24268 3488 24593 3516
rect 24268 3476 24274 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 22097 3451 22155 3457
rect 22097 3448 22109 3451
rect 17788 3420 22109 3448
rect 22097 3417 22109 3420
rect 22143 3417 22155 3451
rect 22097 3411 22155 3417
rect 23293 3451 23351 3457
rect 23293 3417 23305 3451
rect 23339 3417 23351 3451
rect 23293 3411 23351 3417
rect 17402 3380 17408 3392
rect 16991 3352 17264 3380
rect 17363 3352 17408 3380
rect 16991 3349 17003 3352
rect 16945 3343 17003 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17920 3352 18245 3380
rect 17920 3340 17926 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 23308 3380 23336 3411
rect 20772 3352 23336 3380
rect 23753 3383 23811 3389
rect 20772 3340 20778 3352
rect 23753 3349 23765 3383
rect 23799 3380 23811 3383
rect 24854 3380 24860 3392
rect 23799 3352 24860 3380
rect 23799 3349 23811 3352
rect 23753 3343 23811 3349
rect 24854 3340 24860 3352
rect 24912 3340 24918 3392
rect 25148 3380 25176 3556
rect 25240 3525 25268 3692
rect 25593 3689 25605 3723
rect 25639 3689 25651 3723
rect 25593 3683 25651 3689
rect 25608 3652 25636 3683
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 27522 3720 27528 3732
rect 25924 3692 27528 3720
rect 25924 3680 25930 3692
rect 27522 3680 27528 3692
rect 27580 3680 27586 3732
rect 28997 3723 29055 3729
rect 28997 3689 29009 3723
rect 29043 3720 29055 3723
rect 29546 3720 29552 3732
rect 29043 3692 29552 3720
rect 29043 3689 29055 3692
rect 28997 3683 29055 3689
rect 29546 3680 29552 3692
rect 29604 3680 29610 3732
rect 31294 3680 31300 3732
rect 31352 3720 31358 3732
rect 31481 3723 31539 3729
rect 31481 3720 31493 3723
rect 31352 3692 31493 3720
rect 31352 3680 31358 3692
rect 31481 3689 31493 3692
rect 31527 3689 31539 3723
rect 31481 3683 31539 3689
rect 31726 3692 31984 3720
rect 28810 3652 28816 3664
rect 25608 3624 28816 3652
rect 28810 3612 28816 3624
rect 28868 3612 28874 3664
rect 29178 3612 29184 3664
rect 29236 3652 29242 3664
rect 30190 3652 30196 3664
rect 29236 3624 30196 3652
rect 29236 3612 29242 3624
rect 30190 3612 30196 3624
rect 30248 3612 30254 3664
rect 31726 3652 31754 3692
rect 31220 3624 31754 3652
rect 31956 3652 31984 3692
rect 32214 3680 32220 3732
rect 32272 3720 32278 3732
rect 34238 3720 34244 3732
rect 32272 3692 34244 3720
rect 32272 3680 32278 3692
rect 34238 3680 34244 3692
rect 34296 3680 34302 3732
rect 36173 3655 36231 3661
rect 36173 3652 36185 3655
rect 31956 3624 36185 3652
rect 25590 3544 25596 3596
rect 25648 3584 25654 3596
rect 25648 3556 29408 3584
rect 25648 3544 25654 3556
rect 25225 3519 25283 3525
rect 25225 3485 25237 3519
rect 25271 3485 25283 3519
rect 26510 3516 26516 3528
rect 26471 3488 26516 3516
rect 25225 3479 25283 3485
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 26786 3476 26792 3528
rect 26844 3516 26850 3528
rect 26973 3519 27031 3525
rect 26973 3516 26985 3519
rect 26844 3488 26985 3516
rect 26844 3476 26850 3488
rect 26973 3485 26985 3488
rect 27019 3485 27031 3519
rect 27798 3516 27804 3528
rect 27759 3488 27804 3516
rect 26973 3479 27031 3485
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28626 3516 28632 3528
rect 28587 3488 28632 3516
rect 28626 3476 28632 3488
rect 28684 3476 28690 3528
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 25409 3451 25467 3457
rect 25409 3448 25421 3451
rect 25372 3420 25421 3448
rect 25372 3408 25378 3420
rect 25409 3417 25421 3420
rect 25455 3417 25467 3451
rect 28350 3448 28356 3460
rect 25409 3411 25467 3417
rect 26068 3420 28356 3448
rect 26068 3380 26096 3420
rect 28350 3408 28356 3420
rect 28408 3448 28414 3460
rect 28813 3451 28871 3457
rect 28813 3448 28825 3451
rect 28408 3420 28825 3448
rect 28408 3408 28414 3420
rect 28813 3417 28825 3420
rect 28859 3448 28871 3451
rect 29270 3448 29276 3460
rect 28859 3420 29276 3448
rect 28859 3417 28871 3420
rect 28813 3411 28871 3417
rect 29270 3408 29276 3420
rect 29328 3408 29334 3460
rect 29380 3448 29408 3556
rect 29546 3544 29552 3596
rect 29604 3584 29610 3596
rect 29822 3584 29828 3596
rect 29604 3556 29828 3584
rect 29604 3544 29610 3556
rect 29822 3544 29828 3556
rect 29880 3544 29886 3596
rect 30006 3584 30012 3596
rect 29967 3556 30012 3584
rect 30006 3544 30012 3556
rect 30064 3544 30070 3596
rect 31220 3584 31248 3624
rect 36173 3621 36185 3624
rect 36219 3621 36231 3655
rect 36173 3615 36231 3621
rect 30852 3556 31248 3584
rect 29454 3476 29460 3528
rect 29512 3516 29518 3528
rect 30285 3519 30343 3525
rect 30285 3516 30297 3519
rect 29512 3488 30297 3516
rect 29512 3476 29518 3488
rect 30285 3485 30297 3488
rect 30331 3485 30343 3519
rect 30285 3479 30343 3485
rect 30852 3448 30880 3556
rect 31938 3544 31944 3596
rect 31996 3584 32002 3596
rect 31996 3556 32812 3584
rect 31996 3544 32002 3556
rect 30926 3476 30932 3528
rect 30984 3516 30990 3528
rect 32784 3525 32812 3556
rect 37642 3544 37648 3596
rect 37700 3584 37706 3596
rect 37829 3587 37887 3593
rect 37829 3584 37841 3587
rect 37700 3556 37841 3584
rect 37700 3544 37706 3556
rect 37829 3553 37841 3556
rect 37875 3553 37887 3587
rect 37829 3547 37887 3553
rect 32033 3519 32091 3525
rect 30984 3488 31524 3516
rect 30984 3476 30990 3488
rect 31386 3448 31392 3460
rect 29380 3420 30880 3448
rect 30944 3420 31392 3448
rect 25148 3352 26096 3380
rect 26142 3340 26148 3392
rect 26200 3380 26206 3392
rect 26329 3383 26387 3389
rect 26329 3380 26341 3383
rect 26200 3352 26341 3380
rect 26200 3340 26206 3352
rect 26329 3349 26341 3352
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 26878 3340 26884 3392
rect 26936 3380 26942 3392
rect 27157 3383 27215 3389
rect 27157 3380 27169 3383
rect 26936 3352 27169 3380
rect 26936 3340 26942 3352
rect 27157 3349 27169 3352
rect 27203 3349 27215 3383
rect 27157 3343 27215 3349
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 27985 3383 28043 3389
rect 27985 3380 27997 3383
rect 27764 3352 27997 3380
rect 27764 3340 27770 3352
rect 27985 3349 27997 3352
rect 28031 3349 28043 3383
rect 27985 3343 28043 3349
rect 28442 3340 28448 3392
rect 28500 3380 28506 3392
rect 30558 3380 30564 3392
rect 28500 3352 30564 3380
rect 28500 3340 28506 3352
rect 30558 3340 30564 3352
rect 30616 3340 30622 3392
rect 30742 3340 30748 3392
rect 30800 3380 30806 3392
rect 30944 3380 30972 3420
rect 31386 3408 31392 3420
rect 31444 3408 31450 3460
rect 31496 3448 31524 3488
rect 32033 3485 32045 3519
rect 32079 3485 32091 3519
rect 32033 3479 32091 3485
rect 32769 3519 32827 3525
rect 32769 3485 32781 3519
rect 32815 3485 32827 3519
rect 33870 3516 33876 3528
rect 33831 3488 33876 3516
rect 32769 3479 32827 3485
rect 32048 3448 32076 3479
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 34514 3476 34520 3528
rect 34572 3516 34578 3528
rect 34790 3516 34796 3528
rect 34572 3488 34796 3516
rect 34572 3476 34578 3488
rect 34790 3476 34796 3488
rect 34848 3516 34854 3528
rect 35253 3519 35311 3525
rect 35253 3516 35265 3519
rect 34848 3488 35265 3516
rect 34848 3476 34854 3488
rect 35253 3485 35265 3488
rect 35299 3485 35311 3519
rect 35253 3479 35311 3485
rect 36538 3476 36544 3528
rect 36596 3516 36602 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 36596 3488 38117 3516
rect 36596 3476 36602 3488
rect 38105 3485 38117 3488
rect 38151 3516 38163 3519
rect 38194 3516 38200 3528
rect 38151 3488 38200 3516
rect 38151 3485 38163 3488
rect 38105 3479 38163 3485
rect 38194 3476 38200 3488
rect 38252 3476 38258 3528
rect 31496 3420 32076 3448
rect 33042 3408 33048 3460
rect 33100 3448 33106 3460
rect 35069 3451 35127 3457
rect 35069 3448 35081 3451
rect 33100 3420 35081 3448
rect 33100 3408 33106 3420
rect 35069 3417 35081 3420
rect 35115 3417 35127 3451
rect 35069 3411 35127 3417
rect 36357 3451 36415 3457
rect 36357 3417 36369 3451
rect 36403 3448 36415 3451
rect 38378 3448 38384 3460
rect 36403 3420 38384 3448
rect 36403 3417 36415 3420
rect 36357 3411 36415 3417
rect 38378 3408 38384 3420
rect 38436 3408 38442 3460
rect 30800 3352 30972 3380
rect 30800 3340 30806 3352
rect 31018 3340 31024 3392
rect 31076 3380 31082 3392
rect 32217 3383 32275 3389
rect 32217 3380 32229 3383
rect 31076 3352 32229 3380
rect 31076 3340 31082 3352
rect 32217 3349 32229 3352
rect 32263 3349 32275 3383
rect 32217 3343 32275 3349
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 32953 3383 33011 3389
rect 32953 3380 32965 3383
rect 32732 3352 32965 3380
rect 32732 3340 32738 3352
rect 32953 3349 32965 3352
rect 32999 3349 33011 3383
rect 32953 3343 33011 3349
rect 34057 3383 34115 3389
rect 34057 3349 34069 3383
rect 34103 3380 34115 3383
rect 34330 3380 34336 3392
rect 34103 3352 34336 3380
rect 34103 3349 34115 3352
rect 34057 3343 34115 3349
rect 34330 3340 34336 3352
rect 34388 3340 34394 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3510 3176 3516 3188
rect 3467 3148 3516 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 5718 3176 5724 3188
rect 4847 3148 5724 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 9306 3176 9312 3188
rect 5859 3148 9312 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9582 3176 9588 3188
rect 9543 3148 9588 3176
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 10560 3148 12449 3176
rect 10560 3136 10566 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 13596 3148 13737 3176
rect 13596 3136 13602 3148
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 13725 3139 13783 3145
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14424 3148 14565 3176
rect 14424 3136 14430 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 14553 3139 14611 3145
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3145 15991 3179
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 15933 3139 15991 3145
rect 3326 3068 3332 3120
rect 3384 3108 3390 3120
rect 3786 3108 3792 3120
rect 3384 3080 3792 3108
rect 3384 3068 3390 3080
rect 3786 3068 3792 3080
rect 3844 3108 3850 3120
rect 3973 3111 4031 3117
rect 3973 3108 3985 3111
rect 3844 3080 3985 3108
rect 3844 3068 3850 3080
rect 3973 3077 3985 3080
rect 4019 3077 4031 3111
rect 4706 3108 4712 3120
rect 4667 3080 4712 3108
rect 3973 3071 4031 3077
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 6638 3108 6644 3120
rect 5592 3080 6644 3108
rect 5592 3068 5598 3080
rect 6638 3068 6644 3080
rect 6696 3108 6702 3120
rect 6825 3111 6883 3117
rect 6825 3108 6837 3111
rect 6696 3080 6837 3108
rect 6696 3068 6702 3080
rect 6825 3077 6837 3080
rect 6871 3077 6883 3111
rect 6825 3071 6883 3077
rect 7009 3111 7067 3117
rect 7009 3077 7021 3111
rect 7055 3108 7067 3111
rect 7926 3108 7932 3120
rect 7055 3080 7932 3108
rect 7055 3077 7067 3080
rect 7009 3071 7067 3077
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 14090 3108 14096 3120
rect 8220 3080 14096 3108
rect 1118 3000 1124 3052
rect 1176 3040 1182 3052
rect 1394 3040 1400 3052
rect 1176 3012 1400 3040
rect 1176 3000 1182 3012
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 2866 2972 2872 2984
rect 2827 2944 2872 2972
rect 1673 2935 1731 2941
rect 106 2796 112 2848
rect 164 2836 170 2848
rect 1394 2836 1400 2848
rect 164 2808 1400 2836
rect 164 2796 170 2808
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 1688 2836 1716 2935
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3068 2972 3096 3003
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4724 3040 4752 3068
rect 5626 3040 5632 3052
rect 3936 3012 4752 3040
rect 5587 3012 5632 3040
rect 3936 3000 3942 3012
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 8076 3012 8125 3040
rect 8076 3000 8082 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 4890 2972 4896 2984
rect 3068 2944 4896 2972
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 8220 2904 8248 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14274 3068 14280 3120
rect 14332 3108 14338 3120
rect 15948 3108 15976 3139
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 18598 3176 18604 3188
rect 18559 3148 18604 3176
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 20036 3148 20085 3176
rect 20036 3136 20042 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 20588 3148 37596 3176
rect 20588 3136 20594 3148
rect 14332 3080 15976 3108
rect 14332 3068 14338 3080
rect 16390 3068 16396 3120
rect 16448 3108 16454 3120
rect 17402 3108 17408 3120
rect 16448 3080 17408 3108
rect 16448 3068 16454 3080
rect 17402 3068 17408 3080
rect 17460 3068 17466 3120
rect 17954 3108 17960 3120
rect 17915 3080 17960 3108
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18966 3068 18972 3120
rect 19024 3108 19030 3120
rect 20162 3108 20168 3120
rect 19024 3080 20168 3108
rect 19024 3068 19030 3080
rect 8386 3040 8392 3052
rect 8347 3012 8392 3040
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 9674 3040 9680 3052
rect 9447 3012 9680 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 10008 3012 10057 3040
rect 10008 3000 10014 3012
rect 10045 3009 10057 3012
rect 10091 3040 10103 3043
rect 10134 3040 10140 3052
rect 10091 3012 10140 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10318 3040 10324 3052
rect 10279 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 11330 3000 11336 3052
rect 11388 3040 11394 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11388 3012 11529 3040
rect 11388 3000 11394 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 12250 3040 12256 3052
rect 12211 3012 12256 3040
rect 11517 3003 11575 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12676 3012 13001 3040
rect 12676 3000 12682 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 14366 3040 14372 3052
rect 14279 3012 14372 3040
rect 13909 3003 13967 3009
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 9122 2972 9128 2984
rect 8904 2944 9128 2972
rect 8904 2932 8910 2944
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9582 2904 9588 2916
rect 4203 2876 8248 2904
rect 8312 2876 9588 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 5442 2836 5448 2848
rect 1688 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 7561 2839 7619 2845
rect 7561 2836 7573 2839
rect 7064 2808 7573 2836
rect 7064 2796 7070 2808
rect 7561 2805 7573 2808
rect 7607 2836 7619 2839
rect 8312 2836 8340 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 9692 2904 9720 3000
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 13354 2972 13360 2984
rect 12492 2944 13360 2972
rect 12492 2932 12498 2944
rect 13354 2932 13360 2944
rect 13412 2972 13418 2984
rect 13924 2972 13952 3003
rect 14366 3000 14372 3012
rect 14424 3040 14430 3052
rect 14642 3040 14648 3052
rect 14424 3012 14648 3040
rect 14424 3000 14430 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 15068 3012 15209 3040
rect 15068 3000 15074 3012
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15746 3040 15752 3052
rect 15197 3003 15255 3009
rect 15304 3012 15752 3040
rect 13412 2944 13952 2972
rect 13412 2932 13418 2944
rect 10778 2904 10784 2916
rect 9692 2876 10784 2904
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 13173 2907 13231 2913
rect 13173 2904 13185 2907
rect 11388 2876 13185 2904
rect 11388 2864 11394 2876
rect 13173 2873 13185 2876
rect 13219 2873 13231 2907
rect 13173 2867 13231 2873
rect 13262 2864 13268 2916
rect 13320 2904 13326 2916
rect 15304 2904 15332 3012
rect 15746 3000 15752 3012
rect 15804 3040 15810 3052
rect 16117 3043 16175 3049
rect 16117 3040 16129 3043
rect 15804 3012 16129 3040
rect 15804 3000 15810 3012
rect 16117 3009 16129 3012
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 17218 3040 17224 3052
rect 16715 3012 17224 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16684 2972 16712 3003
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 17736 3012 17785 3040
rect 17736 3000 17742 3012
rect 17773 3009 17785 3012
rect 17819 3040 17831 3043
rect 18046 3040 18052 3052
rect 17819 3012 18052 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 18380 3012 18429 3040
rect 18380 3000 18386 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 18417 3003 18475 3009
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 19904 3049 19932 3080
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 22922 3108 22928 3120
rect 21008 3080 22928 3108
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20438 3040 20444 3052
rect 20036 3012 20444 3040
rect 20036 3000 20042 3012
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 21008 3049 21036 3080
rect 22922 3068 22928 3080
rect 22980 3068 22986 3120
rect 23106 3068 23112 3120
rect 23164 3108 23170 3120
rect 23842 3108 23848 3120
rect 23164 3080 23848 3108
rect 23164 3068 23170 3080
rect 23842 3068 23848 3080
rect 23900 3108 23906 3120
rect 24029 3111 24087 3117
rect 24029 3108 24041 3111
rect 23900 3080 24041 3108
rect 23900 3068 23906 3080
rect 24029 3077 24041 3080
rect 24075 3077 24087 3111
rect 24029 3071 24087 3077
rect 24118 3068 24124 3120
rect 24176 3108 24182 3120
rect 24213 3111 24271 3117
rect 24213 3108 24225 3111
rect 24176 3080 24225 3108
rect 24176 3068 24182 3080
rect 24213 3077 24225 3080
rect 24259 3077 24271 3111
rect 24213 3071 24271 3077
rect 24578 3068 24584 3120
rect 24636 3108 24642 3120
rect 24765 3111 24823 3117
rect 24765 3108 24777 3111
rect 24636 3080 24777 3108
rect 24636 3068 24642 3080
rect 24765 3077 24777 3080
rect 24811 3077 24823 3111
rect 24765 3071 24823 3077
rect 24949 3111 25007 3117
rect 24949 3077 24961 3111
rect 24995 3108 25007 3111
rect 25498 3108 25504 3120
rect 24995 3080 25504 3108
rect 24995 3077 25007 3080
rect 24949 3071 25007 3077
rect 25498 3068 25504 3080
rect 25556 3068 25562 3120
rect 27430 3068 27436 3120
rect 27488 3108 27494 3120
rect 27709 3111 27767 3117
rect 27709 3108 27721 3111
rect 27488 3080 27721 3108
rect 27488 3068 27494 3080
rect 27709 3077 27721 3080
rect 27755 3108 27767 3111
rect 27982 3108 27988 3120
rect 27755 3080 27988 3108
rect 27755 3077 27767 3080
rect 27709 3071 27767 3077
rect 27982 3068 27988 3080
rect 28040 3068 28046 3120
rect 28350 3108 28356 3120
rect 28311 3080 28356 3108
rect 28350 3068 28356 3080
rect 28408 3068 28414 3120
rect 28810 3068 28816 3120
rect 28868 3108 28874 3120
rect 29730 3108 29736 3120
rect 28868 3080 29736 3108
rect 28868 3068 28874 3080
rect 29730 3068 29736 3080
rect 29788 3068 29794 3120
rect 34422 3108 34428 3120
rect 31726 3080 34428 3108
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3009 21051 3043
rect 20993 3003 21051 3009
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22646 3040 22652 3052
rect 22152 3012 22197 3040
rect 22607 3012 22652 3040
rect 22152 3000 22158 3012
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 23382 3000 23388 3052
rect 23440 3040 23446 3052
rect 24596 3040 24624 3068
rect 25406 3040 25412 3052
rect 23440 3012 24624 3040
rect 25367 3012 25412 3040
rect 23440 3000 23446 3012
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 25958 3000 25964 3052
rect 26016 3040 26022 3052
rect 26145 3043 26203 3049
rect 26145 3040 26157 3043
rect 26016 3012 26157 3040
rect 26016 3000 26022 3012
rect 26145 3009 26157 3012
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 28074 3000 28080 3052
rect 28132 3040 28138 3052
rect 28718 3040 28724 3052
rect 28132 3012 28724 3040
rect 28132 3000 28138 3012
rect 28718 3000 28724 3012
rect 28776 3040 28782 3052
rect 28997 3043 29055 3049
rect 28997 3040 29009 3043
rect 28776 3012 29009 3040
rect 28776 3000 28782 3012
rect 28997 3009 29009 3012
rect 29043 3009 29055 3043
rect 28997 3003 29055 3009
rect 29362 3000 29368 3052
rect 29420 3040 29426 3052
rect 29549 3043 29607 3049
rect 29549 3040 29561 3043
rect 29420 3012 29561 3040
rect 29420 3000 29426 3012
rect 29549 3009 29561 3012
rect 29595 3009 29607 3043
rect 29549 3003 29607 3009
rect 30466 3000 30472 3052
rect 30524 3040 30530 3052
rect 30561 3043 30619 3049
rect 30561 3040 30573 3043
rect 30524 3012 30573 3040
rect 30524 3000 30530 3012
rect 30561 3009 30573 3012
rect 30607 3009 30619 3043
rect 30834 3040 30840 3052
rect 30795 3012 30840 3040
rect 30561 3003 30619 3009
rect 30834 3000 30840 3012
rect 30892 3000 30898 3052
rect 15988 2944 16712 2972
rect 15988 2932 15994 2944
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 18340 2972 18368 3000
rect 16816 2944 18368 2972
rect 22925 2975 22983 2981
rect 16816 2932 16822 2944
rect 22925 2941 22937 2975
rect 22971 2972 22983 2975
rect 31726 2972 31754 3080
rect 34422 3068 34428 3080
rect 34480 3068 34486 3120
rect 35434 3068 35440 3120
rect 35492 3108 35498 3120
rect 35710 3108 35716 3120
rect 35492 3080 35716 3108
rect 35492 3068 35498 3080
rect 35710 3068 35716 3080
rect 35768 3068 35774 3120
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 32493 3043 32551 3049
rect 32493 3040 32505 3043
rect 32456 3012 32505 3040
rect 32456 3000 32462 3012
rect 32493 3009 32505 3012
rect 32539 3040 32551 3043
rect 32582 3040 32588 3052
rect 32539 3012 32588 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 32582 3000 32588 3012
rect 32640 3000 32646 3052
rect 32769 3043 32827 3049
rect 32769 3009 32781 3043
rect 32815 3040 32827 3043
rect 32950 3040 32956 3052
rect 32815 3012 32956 3040
rect 32815 3009 32827 3012
rect 32769 3003 32827 3009
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 33778 3040 33784 3052
rect 33739 3012 33784 3040
rect 33778 3000 33784 3012
rect 33836 3000 33842 3052
rect 34885 3043 34943 3049
rect 34885 3009 34897 3043
rect 34931 3009 34943 3043
rect 34885 3003 34943 3009
rect 35069 3043 35127 3049
rect 35069 3009 35081 3043
rect 35115 3040 35127 3043
rect 35526 3040 35532 3052
rect 35115 3012 35532 3040
rect 35115 3009 35127 3012
rect 35069 3003 35127 3009
rect 22971 2944 31754 2972
rect 22971 2941 22983 2944
rect 22925 2935 22983 2941
rect 33318 2932 33324 2984
rect 33376 2972 33382 2984
rect 34900 2972 34928 3003
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 36446 3040 36452 3052
rect 36407 3012 36452 3040
rect 36446 3000 36452 3012
rect 36504 3000 36510 3052
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 37458 3040 37464 3052
rect 37323 3012 37464 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 37458 3000 37464 3012
rect 37516 3000 37522 3052
rect 37568 3049 37596 3148
rect 37553 3043 37611 3049
rect 37553 3009 37565 3043
rect 37599 3009 37611 3043
rect 37553 3003 37611 3009
rect 38746 2972 38752 2984
rect 33376 2944 38752 2972
rect 33376 2932 33382 2944
rect 38746 2932 38752 2944
rect 38804 2932 38810 2984
rect 13320 2876 15332 2904
rect 13320 2864 13326 2876
rect 16298 2864 16304 2916
rect 16356 2904 16362 2916
rect 20714 2904 20720 2916
rect 16356 2876 20720 2904
rect 16356 2864 16362 2876
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 24486 2864 24492 2916
rect 24544 2904 24550 2916
rect 24544 2876 24992 2904
rect 24544 2864 24550 2876
rect 7607 2808 8340 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 8996 2808 11713 2836
rect 8996 2796 9002 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 11701 2799 11759 2805
rect 12526 2796 12532 2848
rect 12584 2836 12590 2848
rect 13078 2836 13084 2848
rect 12584 2808 13084 2836
rect 12584 2796 12590 2808
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 13630 2836 13636 2848
rect 13412 2808 13636 2836
rect 13412 2796 13418 2808
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 19245 2839 19303 2845
rect 19245 2836 19257 2839
rect 18748 2808 19257 2836
rect 18748 2796 18754 2808
rect 19245 2805 19257 2808
rect 19291 2805 19303 2839
rect 19245 2799 19303 2805
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20404 2808 20821 2836
rect 20404 2796 20410 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 21913 2839 21971 2845
rect 21913 2836 21925 2839
rect 21232 2808 21925 2836
rect 21232 2796 21238 2808
rect 21913 2805 21925 2808
rect 21959 2805 21971 2839
rect 24964 2836 24992 2876
rect 25314 2864 25320 2916
rect 25372 2904 25378 2916
rect 26329 2907 26387 2913
rect 26329 2904 26341 2907
rect 25372 2876 26341 2904
rect 25372 2864 25378 2876
rect 26329 2873 26341 2876
rect 26375 2873 26387 2907
rect 27522 2904 27528 2916
rect 27483 2876 27528 2904
rect 26329 2867 26387 2873
rect 27522 2864 27528 2876
rect 27580 2864 27586 2916
rect 27890 2864 27896 2916
rect 27948 2904 27954 2916
rect 28813 2907 28871 2913
rect 28813 2904 28825 2907
rect 27948 2876 28825 2904
rect 27948 2864 27954 2876
rect 28813 2873 28825 2876
rect 28859 2873 28871 2907
rect 28813 2867 28871 2873
rect 33594 2864 33600 2916
rect 33652 2904 33658 2916
rect 35710 2904 35716 2916
rect 33652 2876 35716 2904
rect 33652 2864 33658 2876
rect 35710 2864 35716 2876
rect 35768 2864 35774 2916
rect 36354 2864 36360 2916
rect 36412 2904 36418 2916
rect 36633 2907 36691 2913
rect 36633 2904 36645 2907
rect 36412 2876 36645 2904
rect 36412 2864 36418 2876
rect 36633 2873 36645 2876
rect 36679 2873 36691 2907
rect 36633 2867 36691 2873
rect 25593 2839 25651 2845
rect 25593 2836 25605 2839
rect 24964 2808 25605 2836
rect 21913 2799 21971 2805
rect 25593 2805 25605 2808
rect 25639 2805 25651 2839
rect 25593 2799 25651 2805
rect 25682 2796 25688 2848
rect 25740 2836 25746 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 25740 2808 26985 2836
rect 25740 2796 25746 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 26973 2799 27031 2805
rect 33502 2796 33508 2848
rect 33560 2836 33566 2848
rect 33965 2839 34023 2845
rect 33965 2836 33977 2839
rect 33560 2808 33977 2836
rect 33560 2796 33566 2808
rect 33965 2805 33977 2808
rect 34011 2805 34023 2839
rect 35618 2836 35624 2848
rect 35579 2808 35624 2836
rect 33965 2799 34023 2805
rect 35618 2796 35624 2808
rect 35676 2796 35682 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 6595 2635 6653 2641
rect 6595 2601 6607 2635
rect 6641 2632 6653 2635
rect 9858 2632 9864 2644
rect 6641 2604 9864 2632
rect 6641 2601 6653 2604
rect 6595 2595 6653 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10686 2632 10692 2644
rect 10647 2604 10692 2632
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 13354 2632 13360 2644
rect 13315 2604 13360 2632
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 15102 2632 15108 2644
rect 15063 2604 15108 2632
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 16853 2635 16911 2641
rect 16853 2601 16865 2635
rect 16899 2632 16911 2635
rect 16942 2632 16948 2644
rect 16899 2604 16948 2632
rect 16899 2601 16911 2604
rect 16853 2595 16911 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17552 2604 17601 2632
rect 17552 2592 17558 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 21266 2632 21272 2644
rect 17589 2595 17647 2601
rect 18432 2604 21272 2632
rect 4065 2567 4123 2573
rect 4065 2533 4077 2567
rect 4111 2564 4123 2567
rect 8754 2564 8760 2576
rect 4111 2536 8760 2564
rect 4111 2533 4123 2536
rect 4065 2527 4123 2533
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 9180 2536 9352 2564
rect 9180 2524 9186 2536
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 3050 2496 3056 2508
rect 1719 2468 3056 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 4488 2468 4537 2496
rect 4488 2456 4494 2468
rect 4525 2465 4537 2468
rect 4571 2496 4583 2499
rect 4614 2496 4620 2508
rect 4571 2468 4620 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 9030 2496 9036 2508
rect 4847 2468 9036 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9214 2496 9220 2508
rect 9175 2468 9220 2496
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9324 2496 9352 2536
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 9732 2536 12817 2564
rect 9732 2524 9738 2536
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 15933 2567 15991 2573
rect 15933 2533 15945 2567
rect 15979 2564 15991 2567
rect 18432 2564 18460 2604
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 28813 2635 28871 2641
rect 28813 2632 28825 2635
rect 22152 2604 28825 2632
rect 22152 2592 22158 2604
rect 28813 2601 28825 2604
rect 28859 2601 28871 2635
rect 28813 2595 28871 2601
rect 34698 2592 34704 2644
rect 34756 2632 34762 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34756 2604 34897 2632
rect 34756 2592 34762 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 15979 2536 18460 2564
rect 18509 2567 18567 2573
rect 15979 2533 15991 2536
rect 15933 2527 15991 2533
rect 18509 2533 18521 2567
rect 18555 2564 18567 2567
rect 18782 2564 18788 2576
rect 18555 2536 18788 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 18782 2524 18788 2536
rect 18840 2524 18846 2576
rect 19426 2524 19432 2576
rect 19484 2564 19490 2576
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 19484 2536 20545 2564
rect 19484 2524 19490 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 26145 2567 26203 2573
rect 26145 2564 26157 2567
rect 20533 2527 20591 2533
rect 21376 2536 26157 2564
rect 21376 2496 21404 2536
rect 26145 2533 26157 2536
rect 26191 2533 26203 2567
rect 26145 2527 26203 2533
rect 27246 2524 27252 2576
rect 27304 2564 27310 2576
rect 27341 2567 27399 2573
rect 27341 2564 27353 2567
rect 27304 2536 27353 2564
rect 27304 2524 27310 2536
rect 27341 2533 27353 2536
rect 27387 2533 27399 2567
rect 36446 2564 36452 2576
rect 27341 2527 27399 2533
rect 27908 2536 36452 2564
rect 9324 2468 21404 2496
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2496 21971 2499
rect 22278 2496 22284 2508
rect 21959 2468 22284 2496
rect 21959 2465 21971 2468
rect 21913 2459 21971 2465
rect 22278 2456 22284 2468
rect 22336 2456 22342 2508
rect 22373 2499 22431 2505
rect 22373 2465 22385 2499
rect 22419 2496 22431 2499
rect 22462 2496 22468 2508
rect 22419 2468 22468 2496
rect 22419 2465 22431 2468
rect 22373 2459 22431 2465
rect 22462 2456 22468 2468
rect 22520 2456 22526 2508
rect 22649 2499 22707 2505
rect 22649 2465 22661 2499
rect 22695 2496 22707 2499
rect 27908 2496 27936 2536
rect 36446 2524 36452 2536
rect 36504 2524 36510 2576
rect 22695 2468 27936 2496
rect 22695 2465 22707 2468
rect 22649 2459 22707 2465
rect 29638 2456 29644 2508
rect 29696 2496 29702 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29696 2468 29745 2496
rect 29696 2456 29702 2468
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 29733 2459 29791 2465
rect 29914 2456 29920 2508
rect 29972 2496 29978 2508
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 29972 2468 30021 2496
rect 29972 2456 29978 2468
rect 30009 2465 30021 2468
rect 30055 2465 30067 2499
rect 30009 2459 30067 2465
rect 31754 2456 31760 2508
rect 31812 2496 31818 2508
rect 32493 2499 32551 2505
rect 32493 2496 32505 2499
rect 31812 2468 32505 2496
rect 31812 2456 31818 2468
rect 32493 2465 32505 2468
rect 32539 2465 32551 2499
rect 32493 2459 32551 2465
rect 35894 2456 35900 2508
rect 35952 2496 35958 2508
rect 36538 2496 36544 2508
rect 35952 2468 36544 2496
rect 35952 2456 35958 2468
rect 36538 2456 36544 2468
rect 36596 2456 36602 2508
rect 37274 2496 37280 2508
rect 37235 2468 37280 2496
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 37553 2499 37611 2505
rect 37553 2465 37565 2499
rect 37599 2496 37611 2499
rect 38838 2496 38844 2508
rect 37599 2468 38844 2496
rect 37599 2465 37611 2468
rect 37553 2459 37611 2465
rect 38838 2456 38844 2468
rect 38896 2456 38902 2508
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2774 2428 2780 2440
rect 2280 2400 2780 2428
rect 2280 2388 2286 2400
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5040 2400 6377 2428
rect 5040 2388 5046 2400
rect 6365 2397 6377 2400
rect 6411 2428 6423 2431
rect 6454 2428 6460 2440
rect 6411 2400 6460 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 6886 2400 7757 2428
rect 1394 2320 1400 2372
rect 1452 2360 1458 2372
rect 1762 2360 1768 2372
rect 1452 2332 1768 2360
rect 1452 2320 1458 2332
rect 1762 2320 1768 2332
rect 1820 2320 1826 2372
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3016 2332 3893 2360
rect 3016 2320 3022 2332
rect 3881 2329 3893 2332
rect 3927 2360 3939 2363
rect 3970 2360 3976 2372
rect 3927 2332 3976 2360
rect 3927 2329 3939 2332
rect 3881 2323 3939 2329
rect 3970 2320 3976 2332
rect 4028 2320 4034 2372
rect 6086 2320 6092 2372
rect 6144 2360 6150 2372
rect 6886 2360 6914 2400
rect 7745 2397 7757 2400
rect 7791 2428 7803 2431
rect 8110 2428 8116 2440
rect 7791 2400 8116 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8846 2388 8852 2440
rect 8904 2428 8910 2440
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 8904 2400 9505 2428
rect 8904 2388 8910 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10594 2428 10600 2440
rect 10284 2400 10600 2428
rect 10284 2388 10290 2400
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 14056 2400 14105 2428
rect 14056 2388 14062 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15712 2400 15761 2428
rect 15712 2388 15718 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 15749 2391 15807 2397
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 17310 2388 17316 2440
rect 17368 2428 17374 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17368 2400 17509 2428
rect 17368 2388 17374 2400
rect 17497 2397 17509 2400
rect 17543 2428 17555 2431
rect 17586 2428 17592 2440
rect 17543 2400 17592 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 19886 2428 19892 2440
rect 19847 2400 19892 2428
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 20349 2431 20407 2437
rect 20349 2428 20361 2431
rect 20312 2400 20361 2428
rect 20312 2388 20318 2400
rect 20349 2397 20361 2400
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 23661 2431 23719 2437
rect 23661 2397 23673 2431
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 6144 2332 6914 2360
rect 7929 2363 7987 2369
rect 6144 2320 6150 2332
rect 7929 2329 7941 2363
rect 7975 2360 7987 2363
rect 10962 2360 10968 2372
rect 7975 2332 10968 2360
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 14182 2360 14188 2372
rect 11900 2332 14188 2360
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 11900 2292 11928 2332
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 18138 2320 18144 2372
rect 18196 2360 18202 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 18196 2332 18337 2360
rect 18196 2320 18202 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 18325 2323 18383 2329
rect 18414 2320 18420 2372
rect 18472 2360 18478 2372
rect 19150 2360 19156 2372
rect 18472 2332 19156 2360
rect 18472 2320 18478 2332
rect 19150 2320 19156 2332
rect 19208 2360 19214 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19208 2332 19717 2360
rect 19208 2320 19214 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 23676 2360 23704 2391
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 24394 2428 24400 2440
rect 23992 2400 24400 2428
rect 23992 2388 23998 2400
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 26329 2431 26387 2437
rect 24719 2400 26234 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 24762 2360 24768 2372
rect 21315 2332 24768 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 12066 2292 12072 2304
rect 8812 2264 11928 2292
rect 12027 2264 12072 2292
rect 8812 2252 8818 2264
rect 12066 2252 12072 2264
rect 12124 2252 12130 2304
rect 14274 2292 14280 2304
rect 14235 2264 14280 2292
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 23842 2292 23848 2304
rect 23803 2264 23848 2292
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 26206 2292 26234 2400
rect 26329 2397 26341 2431
rect 26375 2428 26387 2431
rect 26694 2428 26700 2440
rect 26375 2400 26700 2428
rect 26375 2397 26387 2400
rect 26329 2391 26387 2397
rect 26694 2388 26700 2400
rect 26752 2388 26758 2440
rect 27154 2388 27160 2440
rect 27212 2428 27218 2440
rect 28258 2428 28264 2440
rect 27212 2400 28264 2428
rect 27212 2388 27218 2400
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 28994 2428 29000 2440
rect 28955 2400 29000 2428
rect 28994 2388 29000 2400
rect 29052 2388 29058 2440
rect 29086 2388 29092 2440
rect 29144 2428 29150 2440
rect 30098 2428 30104 2440
rect 29144 2400 30104 2428
rect 29144 2388 29150 2400
rect 30098 2388 30104 2400
rect 30156 2428 30162 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 30156 2400 31217 2428
rect 30156 2388 30162 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 32214 2428 32220 2440
rect 32175 2400 32220 2428
rect 31205 2391 31263 2397
rect 32214 2388 32220 2400
rect 32272 2388 32278 2440
rect 33686 2388 33692 2440
rect 33744 2428 33750 2440
rect 34057 2431 34115 2437
rect 34057 2428 34069 2431
rect 33744 2400 34069 2428
rect 33744 2388 33750 2400
rect 34057 2397 34069 2400
rect 34103 2397 34115 2431
rect 34057 2391 34115 2397
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34664 2400 34713 2428
rect 34664 2388 34670 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 36170 2428 36176 2440
rect 36131 2400 36176 2428
rect 34701 2391 34759 2397
rect 36170 2388 36176 2400
rect 36228 2388 36234 2440
rect 37292 2428 37320 2456
rect 37918 2428 37924 2440
rect 37292 2400 37924 2428
rect 37918 2388 37924 2400
rect 37976 2388 37982 2440
rect 26418 2320 26424 2372
rect 26476 2360 26482 2372
rect 27338 2360 27344 2372
rect 26476 2332 27344 2360
rect 26476 2320 26482 2332
rect 27338 2320 27344 2332
rect 27396 2360 27402 2372
rect 27525 2363 27583 2369
rect 27525 2360 27537 2363
rect 27396 2332 27537 2360
rect 27396 2320 27402 2332
rect 27525 2329 27537 2332
rect 27571 2329 27583 2363
rect 28074 2360 28080 2372
rect 27525 2323 27583 2329
rect 27632 2332 28080 2360
rect 27632 2292 27660 2332
rect 28074 2320 28080 2332
rect 28132 2320 28138 2372
rect 28166 2292 28172 2304
rect 26206 2264 27660 2292
rect 28127 2264 28172 2292
rect 28166 2252 28172 2264
rect 28224 2252 28230 2304
rect 31110 2292 31116 2304
rect 31071 2264 31116 2292
rect 31110 2252 31116 2264
rect 31168 2252 31174 2304
rect 33962 2292 33968 2304
rect 33923 2264 33968 2292
rect 33962 2252 33968 2264
rect 34020 2252 34026 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 16114 2048 16120 2100
rect 16172 2088 16178 2100
rect 36170 2088 36176 2100
rect 16172 2060 36176 2088
rect 16172 2048 16178 2060
rect 36170 2048 36176 2060
rect 36228 2048 36234 2100
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 31110 2020 31116 2032
rect 9824 1992 31116 2020
rect 9824 1980 9830 1992
rect 31110 1980 31116 1992
rect 31168 1980 31174 2032
rect 4890 1912 4896 1964
rect 4948 1952 4954 1964
rect 27522 1952 27528 1964
rect 4948 1924 27528 1952
rect 4948 1912 4954 1924
rect 27522 1912 27528 1924
rect 27580 1912 27586 1964
rect 2866 1844 2872 1896
rect 2924 1884 2930 1896
rect 12526 1884 12532 1896
rect 2924 1856 12532 1884
rect 2924 1844 2930 1856
rect 12526 1844 12532 1856
rect 12584 1844 12590 1896
rect 18874 1844 18880 1896
rect 18932 1884 18938 1896
rect 28166 1884 28172 1896
rect 18932 1856 28172 1884
rect 18932 1844 18938 1856
rect 28166 1844 28172 1856
rect 28224 1844 28230 1896
rect 14458 1776 14464 1828
rect 14516 1816 14522 1828
rect 33962 1816 33968 1828
rect 14516 1788 33968 1816
rect 14516 1776 14522 1788
rect 33962 1776 33968 1788
rect 34020 1776 34026 1828
rect 12066 1708 12072 1760
rect 12124 1748 12130 1760
rect 23014 1748 23020 1760
rect 12124 1720 23020 1748
rect 12124 1708 12130 1720
rect 23014 1708 23020 1720
rect 23072 1708 23078 1760
<< via1 >>
rect 2228 37816 2280 37868
rect 23664 37816 23716 37868
rect 7288 37748 7340 37800
rect 26700 37748 26752 37800
rect 12256 37680 12308 37732
rect 31484 37680 31536 37732
rect 13176 37612 13228 37664
rect 31576 37612 31628 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2228 37408 2280 37460
rect 4896 37408 4948 37460
rect 7288 37408 7340 37460
rect 12256 37451 12308 37460
rect 12256 37417 12265 37451
rect 12265 37417 12299 37451
rect 12299 37417 12308 37451
rect 12256 37408 12308 37417
rect 29092 37408 29144 37460
rect 13176 37383 13228 37392
rect 13176 37349 13185 37383
rect 13185 37349 13219 37383
rect 13219 37349 13228 37383
rect 13176 37340 13228 37349
rect 3700 37272 3752 37324
rect 5264 37272 5316 37324
rect 1124 37204 1176 37256
rect 1952 37204 2004 37256
rect 2136 37204 2188 37256
rect 2596 37204 2648 37256
rect 4160 37204 4212 37256
rect 5080 37247 5132 37256
rect 5080 37213 5089 37247
rect 5089 37213 5123 37247
rect 5123 37213 5132 37247
rect 5080 37204 5132 37213
rect 5724 37204 5776 37256
rect 6368 37204 6420 37256
rect 7472 37204 7524 37256
rect 8484 37204 8536 37256
rect 9404 37247 9456 37256
rect 9404 37213 9413 37247
rect 9413 37213 9447 37247
rect 9447 37213 9456 37247
rect 9404 37204 9456 37213
rect 10140 37204 10192 37256
rect 10600 37204 10652 37256
rect 12164 37204 12216 37256
rect 13820 37204 13872 37256
rect 35992 37340 36044 37392
rect 15844 37272 15896 37324
rect 17408 37272 17460 37324
rect 21916 37272 21968 37324
rect 14832 37204 14884 37256
rect 15108 37204 15160 37256
rect 15936 37204 15988 37256
rect 17500 37204 17552 37256
rect 17960 37204 18012 37256
rect 19064 37204 19116 37256
rect 20076 37204 20128 37256
rect 20904 37247 20956 37256
rect 20904 37213 20913 37247
rect 20913 37213 20947 37247
rect 20947 37213 20956 37247
rect 20904 37204 20956 37213
rect 21088 37204 21140 37256
rect 30656 37315 30708 37324
rect 30656 37281 30665 37315
rect 30665 37281 30699 37315
rect 30699 37281 30708 37315
rect 30656 37272 30708 37281
rect 32496 37315 32548 37324
rect 32496 37281 32505 37315
rect 32505 37281 32539 37315
rect 32539 37281 32548 37315
rect 32496 37272 32548 37281
rect 3240 37136 3292 37188
rect 4068 37136 4120 37188
rect 11612 37136 11664 37188
rect 13176 37136 13228 37188
rect 18052 37136 18104 37188
rect 3056 37068 3108 37120
rect 7840 37111 7892 37120
rect 7840 37077 7849 37111
rect 7849 37077 7883 37111
rect 7883 37077 7892 37111
rect 7840 37068 7892 37077
rect 10416 37111 10468 37120
rect 10416 37077 10425 37111
rect 10425 37077 10459 37111
rect 10459 37077 10468 37111
rect 10416 37068 10468 37077
rect 14004 37068 14056 37120
rect 19432 37111 19484 37120
rect 19432 37077 19441 37111
rect 19441 37077 19475 37111
rect 19475 37077 19484 37111
rect 19432 37068 19484 37077
rect 20352 37111 20404 37120
rect 20352 37077 20361 37111
rect 20361 37077 20395 37111
rect 20395 37077 20404 37111
rect 20352 37068 20404 37077
rect 20444 37068 20496 37120
rect 22192 37136 22244 37188
rect 24308 37204 24360 37256
rect 25320 37204 25372 37256
rect 25504 37204 25556 37256
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 24124 37136 24176 37188
rect 26608 37136 26660 37188
rect 28540 37204 28592 37256
rect 28816 37247 28868 37256
rect 28816 37213 28825 37247
rect 28825 37213 28859 37247
rect 28859 37213 28868 37247
rect 28816 37204 28868 37213
rect 29552 37247 29604 37256
rect 29552 37213 29561 37247
rect 29561 37213 29595 37247
rect 29595 37213 29604 37247
rect 29552 37204 29604 37213
rect 30564 37204 30616 37256
rect 31208 37204 31260 37256
rect 31760 37204 31812 37256
rect 32772 37204 32824 37256
rect 33508 37247 33560 37256
rect 33508 37213 33517 37247
rect 33517 37213 33551 37247
rect 33551 37213 33560 37247
rect 33508 37204 33560 37213
rect 33784 37204 33836 37256
rect 35440 37204 35492 37256
rect 35716 37247 35768 37256
rect 35716 37213 35725 37247
rect 35725 37213 35759 37247
rect 35759 37213 35768 37247
rect 35716 37204 35768 37213
rect 35900 37204 35952 37256
rect 37280 37247 37332 37256
rect 37280 37213 37289 37247
rect 37289 37213 37323 37247
rect 37323 37213 37332 37247
rect 37280 37204 37332 37213
rect 28448 37136 28500 37188
rect 23296 37068 23348 37120
rect 24584 37111 24636 37120
rect 24584 37077 24593 37111
rect 24593 37077 24627 37111
rect 24627 37077 24636 37111
rect 24584 37068 24636 37077
rect 25596 37111 25648 37120
rect 25596 37077 25605 37111
rect 25605 37077 25639 37111
rect 25639 37077 25648 37111
rect 25596 37068 25648 37077
rect 25688 37068 25740 37120
rect 26792 37068 26844 37120
rect 27804 37068 27856 37120
rect 28724 37111 28776 37120
rect 28724 37077 28733 37111
rect 28733 37077 28767 37111
rect 28767 37077 28776 37111
rect 28724 37068 28776 37077
rect 29736 37111 29788 37120
rect 29736 37077 29745 37111
rect 29745 37077 29779 37111
rect 29779 37077 29788 37111
rect 29736 37068 29788 37077
rect 29828 37068 29880 37120
rect 31208 37068 31260 37120
rect 34336 37136 34388 37188
rect 34796 37111 34848 37120
rect 34796 37077 34805 37111
rect 34805 37077 34839 37111
rect 34839 37077 34848 37111
rect 34796 37068 34848 37077
rect 35532 37111 35584 37120
rect 35532 37077 35541 37111
rect 35541 37077 35575 37111
rect 35575 37077 35584 37111
rect 35532 37068 35584 37077
rect 36268 37111 36320 37120
rect 36268 37077 36277 37111
rect 36277 37077 36311 37111
rect 36311 37077 36320 37111
rect 36268 37068 36320 37077
rect 38384 37136 38436 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2504 36864 2556 36916
rect 3608 36864 3660 36916
rect 4620 36864 4672 36916
rect 4988 36864 5040 36916
rect 5816 36864 5868 36916
rect 7748 36864 7800 36916
rect 8852 36864 8904 36916
rect 10968 36864 11020 36916
rect 11980 36864 12032 36916
rect 13084 36864 13136 36916
rect 14096 36864 14148 36916
rect 15200 36864 15252 36916
rect 17224 36864 17276 36916
rect 18328 36864 18380 36916
rect 19340 36864 19392 36916
rect 19984 36864 20036 36916
rect 20812 36864 20864 36916
rect 21456 36864 21508 36916
rect 22560 36864 22612 36916
rect 23572 36864 23624 36916
rect 24860 36864 24912 36916
rect 25044 36864 25096 36916
rect 27068 36864 27120 36916
rect 28172 36864 28224 36916
rect 29184 36864 29236 36916
rect 29920 36864 29972 36916
rect 30932 36864 30984 36916
rect 32036 36864 32088 36916
rect 33140 36864 33192 36916
rect 34152 36864 34204 36916
rect 35348 36864 35400 36916
rect 36360 36864 36412 36916
rect 112 36796 164 36848
rect 1584 36796 1636 36848
rect 3056 36796 3108 36848
rect 7472 36796 7524 36848
rect 12716 36796 12768 36848
rect 13176 36796 13228 36848
rect 16948 36796 17000 36848
rect 2964 36728 3016 36780
rect 4620 36728 4672 36780
rect 5356 36728 5408 36780
rect 5540 36728 5592 36780
rect 5632 36728 5684 36780
rect 6184 36728 6236 36780
rect 7104 36771 7156 36780
rect 7104 36737 7113 36771
rect 7113 36737 7147 36771
rect 7147 36737 7156 36771
rect 7104 36728 7156 36737
rect 7932 36728 7984 36780
rect 8576 36771 8628 36780
rect 8576 36737 8585 36771
rect 8585 36737 8619 36771
rect 8619 36737 8628 36771
rect 8576 36728 8628 36737
rect 9680 36728 9732 36780
rect 10692 36771 10744 36780
rect 10692 36737 10701 36771
rect 10701 36737 10735 36771
rect 10735 36737 10744 36771
rect 10692 36728 10744 36737
rect 12532 36728 12584 36780
rect 14280 36771 14332 36780
rect 9404 36660 9456 36712
rect 14280 36737 14289 36771
rect 14289 36737 14323 36771
rect 14323 36737 14332 36771
rect 14280 36728 14332 36737
rect 15936 36771 15988 36780
rect 15936 36737 15945 36771
rect 15945 36737 15979 36771
rect 15979 36737 15988 36771
rect 15936 36728 15988 36737
rect 14832 36660 14884 36712
rect 14924 36660 14976 36712
rect 18788 36771 18840 36780
rect 2044 36635 2096 36644
rect 2044 36601 2053 36635
rect 2053 36601 2087 36635
rect 2087 36601 2096 36635
rect 2044 36592 2096 36601
rect 6644 36635 6696 36644
rect 6644 36601 6653 36635
rect 6653 36601 6687 36635
rect 6687 36601 6696 36635
rect 6644 36592 6696 36601
rect 6920 36592 6972 36644
rect 13268 36592 13320 36644
rect 17316 36635 17368 36644
rect 17316 36601 17325 36635
rect 17325 36601 17359 36635
rect 17359 36601 17368 36635
rect 17316 36592 17368 36601
rect 18788 36737 18797 36771
rect 18797 36737 18831 36771
rect 18831 36737 18840 36771
rect 18788 36728 18840 36737
rect 20260 36728 20312 36780
rect 20536 36728 20588 36780
rect 20996 36728 21048 36780
rect 22560 36771 22612 36780
rect 22560 36737 22569 36771
rect 22569 36737 22603 36771
rect 22603 36737 22612 36771
rect 22560 36728 22612 36737
rect 23204 36728 23256 36780
rect 23480 36728 23532 36780
rect 24124 36796 24176 36848
rect 31116 36796 31168 36848
rect 34888 36796 34940 36848
rect 35716 36796 35768 36848
rect 38016 36796 38068 36848
rect 21088 36660 21140 36712
rect 21180 36660 21232 36712
rect 25412 36728 25464 36780
rect 26424 36771 26476 36780
rect 26424 36737 26433 36771
rect 26433 36737 26467 36771
rect 26467 36737 26476 36771
rect 26424 36728 26476 36737
rect 26884 36728 26936 36780
rect 27252 36728 27304 36780
rect 28632 36728 28684 36780
rect 29276 36771 29328 36780
rect 29276 36737 29285 36771
rect 29285 36737 29319 36771
rect 29319 36737 29328 36771
rect 29276 36728 29328 36737
rect 30012 36771 30064 36780
rect 30012 36737 30021 36771
rect 30021 36737 30055 36771
rect 30055 36737 30064 36771
rect 30012 36728 30064 36737
rect 31024 36771 31076 36780
rect 31024 36737 31033 36771
rect 31033 36737 31067 36771
rect 31067 36737 31076 36771
rect 31024 36728 31076 36737
rect 31944 36728 31996 36780
rect 33140 36771 33192 36780
rect 33140 36737 33149 36771
rect 33149 36737 33183 36771
rect 33183 36737 33192 36771
rect 33140 36728 33192 36737
rect 34244 36771 34296 36780
rect 34244 36737 34253 36771
rect 34253 36737 34287 36771
rect 34287 36737 34296 36771
rect 34244 36728 34296 36737
rect 34520 36728 34572 36780
rect 36268 36728 36320 36780
rect 24860 36660 24912 36712
rect 37556 36660 37608 36712
rect 18604 36592 18656 36644
rect 1492 36524 1544 36576
rect 6368 36524 6420 36576
rect 6736 36524 6788 36576
rect 23388 36567 23440 36576
rect 23388 36533 23397 36567
rect 23397 36533 23431 36567
rect 23431 36533 23440 36567
rect 23388 36524 23440 36533
rect 23664 36592 23716 36644
rect 24676 36524 24728 36576
rect 26332 36592 26384 36644
rect 38200 36592 38252 36644
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 388 36320 440 36372
rect 1860 36320 1912 36372
rect 2872 36320 2924 36372
rect 3884 36320 3936 36372
rect 5356 36363 5408 36372
rect 5356 36329 5365 36363
rect 5365 36329 5399 36363
rect 5399 36329 5408 36363
rect 5356 36320 5408 36329
rect 6000 36320 6052 36372
rect 7196 36320 7248 36372
rect 7932 36363 7984 36372
rect 7932 36329 7941 36363
rect 7941 36329 7975 36363
rect 7975 36329 7984 36363
rect 7932 36320 7984 36329
rect 8300 36320 8352 36372
rect 9864 36320 9916 36372
rect 10232 36320 10284 36372
rect 11336 36320 11388 36372
rect 12440 36320 12492 36372
rect 13452 36320 13504 36372
rect 14464 36320 14516 36372
rect 16212 36320 16264 36372
rect 16580 36320 16632 36372
rect 17592 36320 17644 36372
rect 18696 36320 18748 36372
rect 20536 36320 20588 36372
rect 20996 36320 21048 36372
rect 21824 36320 21876 36372
rect 14924 36252 14976 36304
rect 15108 36252 15160 36304
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 3240 36159 3292 36168
rect 3240 36125 3249 36159
rect 3249 36125 3283 36159
rect 3283 36125 3292 36159
rect 3240 36116 3292 36125
rect 4712 36116 4764 36168
rect 3148 36048 3200 36100
rect 7012 36116 7064 36168
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 8024 36116 8076 36168
rect 9220 36159 9272 36168
rect 9220 36125 9229 36159
rect 9229 36125 9263 36159
rect 9263 36125 9272 36159
rect 9220 36116 9272 36125
rect 10232 36159 10284 36168
rect 10232 36125 10241 36159
rect 10241 36125 10275 36159
rect 10275 36125 10284 36159
rect 10232 36116 10284 36125
rect 11704 36159 11756 36168
rect 6460 36048 6512 36100
rect 11704 36125 11713 36159
rect 11713 36125 11747 36159
rect 11747 36125 11756 36159
rect 11704 36116 11756 36125
rect 12900 36184 12952 36236
rect 23664 36295 23716 36304
rect 23664 36261 23673 36295
rect 23673 36261 23707 36295
rect 23707 36261 23716 36295
rect 23664 36252 23716 36261
rect 23940 36320 23992 36372
rect 25320 36363 25372 36372
rect 25320 36329 25329 36363
rect 25329 36329 25363 36363
rect 25363 36329 25372 36363
rect 25320 36320 25372 36329
rect 26332 36320 26384 36372
rect 26608 36363 26660 36372
rect 26608 36329 26617 36363
rect 26617 36329 26651 36363
rect 26651 36329 26660 36363
rect 26608 36320 26660 36329
rect 27252 36363 27304 36372
rect 27252 36329 27261 36363
rect 27261 36329 27295 36363
rect 27295 36329 27304 36363
rect 27252 36320 27304 36329
rect 28632 36363 28684 36372
rect 28632 36329 28641 36363
rect 28641 36329 28675 36363
rect 28675 36329 28684 36363
rect 28632 36320 28684 36329
rect 28816 36320 28868 36372
rect 31300 36320 31352 36372
rect 34428 36320 34480 36372
rect 35440 36363 35492 36372
rect 35440 36329 35449 36363
rect 35449 36329 35483 36363
rect 35483 36329 35492 36363
rect 35440 36320 35492 36329
rect 26424 36252 26476 36304
rect 29276 36252 29328 36304
rect 29368 36252 29420 36304
rect 28448 36184 28500 36236
rect 13452 36116 13504 36168
rect 13912 36116 13964 36168
rect 14188 36116 14240 36168
rect 16488 36116 16540 36168
rect 17132 36116 17184 36168
rect 18052 36116 18104 36168
rect 12072 36048 12124 36100
rect 20168 36116 20220 36168
rect 20720 36116 20772 36168
rect 22008 36116 22060 36168
rect 24860 36116 24912 36168
rect 26516 36116 26568 36168
rect 27068 36159 27120 36168
rect 27068 36125 27077 36159
rect 27077 36125 27111 36159
rect 27111 36125 27120 36159
rect 27068 36116 27120 36125
rect 27988 36159 28040 36168
rect 27988 36125 27997 36159
rect 27997 36125 28031 36159
rect 28031 36125 28040 36159
rect 27988 36116 28040 36125
rect 20444 36048 20496 36100
rect 23296 36091 23348 36100
rect 23296 36057 23305 36091
rect 23305 36057 23339 36091
rect 23339 36057 23348 36091
rect 23296 36048 23348 36057
rect 24952 36048 25004 36100
rect 31116 36184 31168 36236
rect 37556 36227 37608 36236
rect 37556 36193 37565 36227
rect 37565 36193 37599 36227
rect 37599 36193 37608 36227
rect 37556 36184 37608 36193
rect 28816 36159 28868 36168
rect 28816 36125 28825 36159
rect 28825 36125 28859 36159
rect 28859 36125 28868 36159
rect 28816 36116 28868 36125
rect 30196 36159 30248 36168
rect 30196 36125 30205 36159
rect 30205 36125 30239 36159
rect 30239 36125 30248 36159
rect 30196 36116 30248 36125
rect 31668 36159 31720 36168
rect 31668 36125 31677 36159
rect 31677 36125 31711 36159
rect 31711 36125 31720 36159
rect 31668 36116 31720 36125
rect 34704 36159 34756 36168
rect 34704 36125 34713 36159
rect 34713 36125 34747 36159
rect 34747 36125 34756 36159
rect 34704 36116 34756 36125
rect 30472 36048 30524 36100
rect 30932 36048 30984 36100
rect 33232 36048 33284 36100
rect 33968 36048 34020 36100
rect 38568 36116 38620 36168
rect 38844 36048 38896 36100
rect 22836 36023 22888 36032
rect 22836 35989 22845 36023
rect 22845 35989 22879 36023
rect 22879 35989 22888 36023
rect 22836 35980 22888 35989
rect 23664 35980 23716 36032
rect 26332 35980 26384 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 756 35776 808 35828
rect 3148 35776 3200 35828
rect 4068 35776 4120 35828
rect 5080 35819 5132 35828
rect 5080 35785 5089 35819
rect 5089 35785 5123 35819
rect 5123 35785 5132 35819
rect 5080 35776 5132 35785
rect 7104 35776 7156 35828
rect 8576 35819 8628 35828
rect 8576 35785 8585 35819
rect 8585 35785 8619 35819
rect 8619 35785 8628 35819
rect 8576 35776 8628 35785
rect 9312 35776 9364 35828
rect 10692 35776 10744 35828
rect 11704 35776 11756 35828
rect 14280 35776 14332 35828
rect 14832 35819 14884 35828
rect 14832 35785 14841 35819
rect 14841 35785 14875 35819
rect 14875 35785 14884 35819
rect 14832 35776 14884 35785
rect 15476 35776 15528 35828
rect 15936 35776 15988 35828
rect 20904 35776 20956 35828
rect 22192 35776 22244 35828
rect 22928 35776 22980 35828
rect 23480 35776 23532 35828
rect 24308 35819 24360 35828
rect 24308 35785 24317 35819
rect 24317 35785 24351 35819
rect 24351 35785 24360 35819
rect 24308 35776 24360 35785
rect 26976 35776 27028 35828
rect 28908 35776 28960 35828
rect 29736 35776 29788 35828
rect 30288 35776 30340 35828
rect 31208 35819 31260 35828
rect 31208 35785 31217 35819
rect 31217 35785 31251 35819
rect 31251 35785 31260 35819
rect 31208 35776 31260 35785
rect 33416 35776 33468 35828
rect 35624 35776 35676 35828
rect 37280 35819 37332 35828
rect 37280 35785 37289 35819
rect 37289 35785 37323 35819
rect 37323 35785 37332 35819
rect 37280 35776 37332 35785
rect 3516 35683 3568 35692
rect 3516 35649 3525 35683
rect 3525 35649 3559 35683
rect 3559 35649 3568 35683
rect 3516 35640 3568 35649
rect 5172 35572 5224 35624
rect 5724 35479 5776 35488
rect 5724 35445 5733 35479
rect 5733 35445 5767 35479
rect 5767 35445 5776 35479
rect 5724 35436 5776 35445
rect 9036 35640 9088 35692
rect 10968 35683 11020 35692
rect 10968 35649 10977 35683
rect 10977 35649 11011 35683
rect 11011 35649 11020 35683
rect 10968 35640 11020 35649
rect 11428 35640 11480 35692
rect 11244 35572 11296 35624
rect 22560 35708 22612 35760
rect 27436 35708 27488 35760
rect 14464 35640 14516 35692
rect 14924 35640 14976 35692
rect 16120 35640 16172 35692
rect 16764 35640 16816 35692
rect 17868 35640 17920 35692
rect 23020 35683 23072 35692
rect 16580 35572 16632 35624
rect 23020 35649 23029 35683
rect 23029 35649 23063 35683
rect 23063 35649 23072 35683
rect 23020 35640 23072 35649
rect 26332 35640 26384 35692
rect 27528 35683 27580 35692
rect 27528 35649 27537 35683
rect 27537 35649 27571 35683
rect 27571 35649 27580 35683
rect 27528 35640 27580 35649
rect 30564 35708 30616 35760
rect 31300 35640 31352 35692
rect 32956 35640 33008 35692
rect 33692 35640 33744 35692
rect 33876 35640 33928 35692
rect 35348 35640 35400 35692
rect 35624 35683 35676 35692
rect 35624 35649 35633 35683
rect 35633 35649 35667 35683
rect 35667 35649 35676 35683
rect 35624 35640 35676 35649
rect 36360 35640 36412 35692
rect 37924 35640 37976 35692
rect 39028 35640 39080 35692
rect 13360 35504 13412 35556
rect 16488 35504 16540 35556
rect 29552 35504 29604 35556
rect 32404 35504 32456 35556
rect 36544 35504 36596 35556
rect 37372 35504 37424 35556
rect 37832 35547 37884 35556
rect 37832 35513 37841 35547
rect 37841 35513 37875 35547
rect 37875 35513 37884 35547
rect 37832 35504 37884 35513
rect 7748 35436 7800 35488
rect 8116 35479 8168 35488
rect 8116 35445 8125 35479
rect 8125 35445 8159 35479
rect 8159 35445 8168 35479
rect 8116 35436 8168 35445
rect 13452 35479 13504 35488
rect 13452 35445 13461 35479
rect 13461 35445 13495 35479
rect 13495 35445 13504 35479
rect 13452 35436 13504 35445
rect 17868 35436 17920 35488
rect 20168 35479 20220 35488
rect 20168 35445 20177 35479
rect 20177 35445 20211 35479
rect 20211 35445 20220 35479
rect 20168 35436 20220 35445
rect 20720 35479 20772 35488
rect 20720 35445 20729 35479
rect 20729 35445 20763 35479
rect 20763 35445 20772 35479
rect 20720 35436 20772 35445
rect 22008 35479 22060 35488
rect 22008 35445 22017 35479
rect 22017 35445 22051 35479
rect 22051 35445 22060 35479
rect 22008 35436 22060 35445
rect 24860 35479 24912 35488
rect 24860 35445 24869 35479
rect 24869 35445 24903 35479
rect 24903 35445 24912 35479
rect 24860 35436 24912 35445
rect 25412 35479 25464 35488
rect 25412 35445 25421 35479
rect 25421 35445 25455 35479
rect 25455 35445 25464 35479
rect 25412 35436 25464 35445
rect 26976 35479 27028 35488
rect 26976 35445 26985 35479
rect 26985 35445 27019 35479
rect 27019 35445 27028 35479
rect 26976 35436 27028 35445
rect 28172 35479 28224 35488
rect 28172 35445 28181 35479
rect 28181 35445 28215 35479
rect 28215 35445 28224 35479
rect 28172 35436 28224 35445
rect 29460 35436 29512 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1584 35275 1636 35284
rect 1584 35241 1593 35275
rect 1593 35241 1627 35275
rect 1627 35241 1636 35275
rect 1584 35232 1636 35241
rect 1952 35232 2004 35284
rect 6184 35275 6236 35284
rect 6184 35241 6193 35275
rect 6193 35241 6227 35275
rect 6227 35241 6236 35275
rect 6184 35232 6236 35241
rect 6736 35275 6788 35284
rect 6736 35241 6745 35275
rect 6745 35241 6779 35275
rect 6779 35241 6788 35275
rect 6736 35232 6788 35241
rect 7472 35232 7524 35284
rect 9588 35232 9640 35284
rect 10140 35232 10192 35284
rect 10232 35232 10284 35284
rect 12164 35275 12216 35284
rect 12164 35241 12173 35275
rect 12173 35241 12207 35275
rect 12207 35241 12216 35275
rect 12164 35232 12216 35241
rect 12716 35275 12768 35284
rect 12716 35241 12725 35275
rect 12725 35241 12759 35275
rect 12759 35241 12768 35275
rect 12716 35232 12768 35241
rect 17500 35275 17552 35284
rect 17500 35241 17509 35275
rect 17509 35241 17543 35275
rect 17543 35241 17552 35275
rect 17500 35232 17552 35241
rect 17960 35232 18012 35284
rect 18604 35275 18656 35284
rect 18604 35241 18613 35275
rect 18613 35241 18647 35275
rect 18647 35241 18656 35275
rect 18604 35232 18656 35241
rect 19064 35232 19116 35284
rect 20076 35275 20128 35284
rect 20076 35241 20085 35275
rect 20085 35241 20119 35275
rect 20119 35241 20128 35275
rect 20076 35232 20128 35241
rect 28816 35232 28868 35284
rect 33508 35275 33560 35284
rect 33508 35241 33517 35275
rect 33517 35241 33551 35275
rect 33551 35241 33560 35275
rect 33508 35232 33560 35241
rect 35808 35232 35860 35284
rect 38292 35232 38344 35284
rect 1676 35164 1728 35216
rect 17224 35164 17276 35216
rect 18788 35164 18840 35216
rect 20536 35207 20588 35216
rect 20536 35173 20545 35207
rect 20545 35173 20579 35207
rect 20579 35173 20588 35207
rect 20536 35164 20588 35173
rect 28172 35164 28224 35216
rect 28908 35164 28960 35216
rect 34520 35164 34572 35216
rect 12532 35096 12584 35148
rect 18420 35096 18472 35148
rect 18604 35096 18656 35148
rect 29460 35096 29512 35148
rect 10784 35028 10836 35080
rect 15108 35071 15160 35080
rect 15108 35037 15117 35071
rect 15117 35037 15151 35071
rect 15151 35037 15160 35071
rect 15108 35028 15160 35037
rect 15752 35071 15804 35080
rect 15752 35037 15761 35071
rect 15761 35037 15795 35071
rect 15795 35037 15804 35071
rect 15752 35028 15804 35037
rect 17224 35028 17276 35080
rect 21180 35028 21232 35080
rect 28448 35028 28500 35080
rect 30564 35028 30616 35080
rect 31668 35028 31720 35080
rect 10968 34960 11020 35012
rect 13176 34960 13228 35012
rect 3884 34935 3936 34944
rect 3884 34901 3893 34935
rect 3893 34901 3927 34935
rect 3927 34901 3936 34935
rect 3884 34892 3936 34901
rect 4712 34892 4764 34944
rect 4804 34892 4856 34944
rect 5540 34935 5592 34944
rect 5540 34901 5549 34935
rect 5549 34901 5583 34935
rect 5583 34901 5592 34935
rect 5540 34892 5592 34901
rect 7104 34892 7156 34944
rect 9036 34935 9088 34944
rect 9036 34901 9045 34935
rect 9045 34901 9079 34935
rect 9079 34901 9088 34935
rect 9036 34892 9088 34901
rect 11428 34892 11480 34944
rect 14464 34935 14516 34944
rect 14464 34901 14473 34935
rect 14473 34901 14507 34935
rect 14507 34901 14516 34935
rect 14464 34892 14516 34901
rect 25504 34960 25556 35012
rect 26240 34960 26292 35012
rect 33140 34960 33192 35012
rect 16764 34892 16816 34944
rect 21088 34935 21140 34944
rect 21088 34901 21097 34935
rect 21097 34901 21131 34935
rect 21131 34901 21140 34935
rect 21088 34892 21140 34901
rect 22468 34892 22520 34944
rect 23020 34892 23072 34944
rect 26424 34935 26476 34944
rect 26424 34901 26433 34935
rect 26433 34901 26467 34935
rect 26467 34901 26476 34935
rect 26424 34892 26476 34901
rect 29000 34935 29052 34944
rect 29000 34901 29009 34935
rect 29009 34901 29043 34935
rect 29043 34901 29052 34935
rect 29000 34892 29052 34901
rect 30380 34892 30432 34944
rect 31024 34892 31076 34944
rect 31944 34935 31996 34944
rect 31944 34901 31953 34935
rect 31953 34901 31987 34935
rect 31987 34901 31996 34935
rect 31944 34892 31996 34901
rect 32956 34935 33008 34944
rect 32956 34901 32965 34935
rect 32965 34901 32999 34935
rect 32999 34901 33008 34935
rect 32956 34892 33008 34901
rect 33600 34892 33652 34944
rect 34244 34892 34296 34944
rect 35900 35028 35952 35080
rect 37280 35028 37332 35080
rect 38752 35028 38804 35080
rect 36452 34960 36504 35012
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2596 34731 2648 34740
rect 2596 34697 2605 34731
rect 2605 34697 2639 34731
rect 2639 34697 2648 34731
rect 2596 34688 2648 34697
rect 12072 34731 12124 34740
rect 12072 34697 12081 34731
rect 12081 34697 12115 34731
rect 12115 34697 12124 34731
rect 12072 34688 12124 34697
rect 12900 34731 12952 34740
rect 12900 34697 12909 34731
rect 12909 34697 12943 34731
rect 12943 34697 12952 34731
rect 12900 34688 12952 34697
rect 13544 34688 13596 34740
rect 15108 34688 15160 34740
rect 16948 34731 17000 34740
rect 16948 34697 16957 34731
rect 16957 34697 16991 34731
rect 16991 34697 17000 34731
rect 16948 34688 17000 34697
rect 2780 34552 2832 34604
rect 3240 34552 3292 34604
rect 9496 34620 9548 34672
rect 27528 34688 27580 34740
rect 36636 34688 36688 34740
rect 5264 34552 5316 34604
rect 9220 34595 9272 34604
rect 9220 34561 9229 34595
rect 9229 34561 9263 34595
rect 9263 34561 9272 34595
rect 13912 34595 13964 34604
rect 9220 34552 9272 34561
rect 13912 34561 13921 34595
rect 13921 34561 13955 34595
rect 13955 34561 13964 34595
rect 13912 34552 13964 34561
rect 14188 34552 14240 34604
rect 14924 34552 14976 34604
rect 18328 34595 18380 34604
rect 18328 34561 18362 34595
rect 18362 34561 18380 34595
rect 18328 34552 18380 34561
rect 2872 34484 2924 34536
rect 9680 34484 9732 34536
rect 9864 34484 9916 34536
rect 10784 34527 10836 34536
rect 10784 34493 10793 34527
rect 10793 34493 10827 34527
rect 10827 34493 10836 34527
rect 10784 34484 10836 34493
rect 11244 34484 11296 34536
rect 13728 34484 13780 34536
rect 20260 34484 20312 34536
rect 20444 34527 20496 34536
rect 20444 34493 20453 34527
rect 20453 34493 20487 34527
rect 20487 34493 20496 34527
rect 20444 34484 20496 34493
rect 27988 34620 28040 34672
rect 37280 34688 37332 34740
rect 38016 34688 38068 34740
rect 37188 34620 37240 34672
rect 39764 34620 39816 34672
rect 23296 34552 23348 34604
rect 26240 34552 26292 34604
rect 27528 34552 27580 34604
rect 37556 34552 37608 34604
rect 24952 34484 25004 34536
rect 32864 34484 32916 34536
rect 33048 34484 33100 34536
rect 33692 34527 33744 34536
rect 33692 34493 33701 34527
rect 33701 34493 33735 34527
rect 33735 34493 33744 34527
rect 33692 34484 33744 34493
rect 34428 34484 34480 34536
rect 36268 34484 36320 34536
rect 37096 34484 37148 34536
rect 24032 34459 24084 34468
rect 5816 34391 5868 34400
rect 5816 34357 5825 34391
rect 5825 34357 5859 34391
rect 5859 34357 5868 34391
rect 5816 34348 5868 34357
rect 19432 34391 19484 34400
rect 19432 34357 19441 34391
rect 19441 34357 19475 34391
rect 19475 34357 19484 34391
rect 19432 34348 19484 34357
rect 19984 34348 20036 34400
rect 24032 34425 24041 34459
rect 24041 34425 24075 34459
rect 24075 34425 24084 34459
rect 24032 34416 24084 34425
rect 39396 34484 39448 34536
rect 35808 34348 35860 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 18052 34187 18104 34196
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 31300 34187 31352 34196
rect 31300 34153 31309 34187
rect 31309 34153 31343 34187
rect 31343 34153 31352 34187
rect 31300 34144 31352 34153
rect 33140 34144 33192 34196
rect 37188 34187 37240 34196
rect 37188 34153 37197 34187
rect 37197 34153 37231 34187
rect 37231 34153 37240 34187
rect 37188 34144 37240 34153
rect 37648 34144 37700 34196
rect 31484 34076 31536 34128
rect 31668 34076 31720 34128
rect 35900 34119 35952 34128
rect 35900 34085 35909 34119
rect 35909 34085 35943 34119
rect 35943 34085 35952 34119
rect 35900 34076 35952 34085
rect 28724 34008 28776 34060
rect 35624 34008 35676 34060
rect 9496 33940 9548 33992
rect 31484 33983 31536 33992
rect 10140 33872 10192 33924
rect 11060 33804 11112 33856
rect 31484 33949 31493 33983
rect 31493 33949 31527 33983
rect 31527 33949 31536 33983
rect 31484 33940 31536 33949
rect 33508 33940 33560 33992
rect 34704 33983 34756 33992
rect 34704 33949 34713 33983
rect 34713 33949 34747 33983
rect 34747 33949 34756 33983
rect 34704 33940 34756 33949
rect 35716 33940 35768 33992
rect 36636 33940 36688 33992
rect 38016 33940 38068 33992
rect 20536 33872 20588 33924
rect 38476 33872 38528 33924
rect 13728 33804 13780 33856
rect 16120 33804 16172 33856
rect 17132 33847 17184 33856
rect 17132 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17184 33847
rect 17132 33804 17184 33813
rect 21272 33804 21324 33856
rect 24032 33804 24084 33856
rect 33876 33847 33928 33856
rect 33876 33813 33885 33847
rect 33885 33813 33919 33847
rect 33919 33813 33928 33847
rect 33876 33804 33928 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 5264 33643 5316 33652
rect 5264 33609 5273 33643
rect 5273 33609 5307 33643
rect 5307 33609 5316 33643
rect 5264 33600 5316 33609
rect 10140 33643 10192 33652
rect 10140 33609 10149 33643
rect 10149 33609 10183 33643
rect 10183 33609 10192 33643
rect 10140 33600 10192 33609
rect 11060 33600 11112 33652
rect 11704 33600 11756 33652
rect 18328 33600 18380 33652
rect 30012 33600 30064 33652
rect 35716 33600 35768 33652
rect 37924 33600 37976 33652
rect 38660 33600 38712 33652
rect 6920 33464 6972 33516
rect 5816 33396 5868 33448
rect 6368 33396 6420 33448
rect 11060 33464 11112 33516
rect 18604 33507 18656 33516
rect 10508 33439 10560 33448
rect 10508 33405 10517 33439
rect 10517 33405 10551 33439
rect 10551 33405 10560 33439
rect 10508 33396 10560 33405
rect 18604 33473 18613 33507
rect 18613 33473 18647 33507
rect 18647 33473 18656 33507
rect 18604 33464 18656 33473
rect 27528 33507 27580 33516
rect 27528 33473 27537 33507
rect 27537 33473 27571 33507
rect 27571 33473 27580 33507
rect 27528 33464 27580 33473
rect 29184 33507 29236 33516
rect 29184 33473 29193 33507
rect 29193 33473 29227 33507
rect 29227 33473 29236 33507
rect 29184 33464 29236 33473
rect 19432 33396 19484 33448
rect 27804 33439 27856 33448
rect 27804 33405 27813 33439
rect 27813 33405 27847 33439
rect 27847 33405 27856 33439
rect 27804 33396 27856 33405
rect 38752 33396 38804 33448
rect 19524 33328 19576 33380
rect 4896 33260 4948 33312
rect 8024 33260 8076 33312
rect 10508 33260 10560 33312
rect 19248 33260 19300 33312
rect 27896 33260 27948 33312
rect 35348 33260 35400 33312
rect 36360 33260 36412 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 18604 33056 18656 33108
rect 28448 33031 28500 33040
rect 28448 32997 28457 33031
rect 28457 32997 28491 33031
rect 28491 32997 28500 33031
rect 28448 32988 28500 32997
rect 36268 32920 36320 32972
rect 37096 32920 37148 32972
rect 19248 32895 19300 32904
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 19524 32895 19576 32904
rect 19524 32861 19533 32895
rect 19533 32861 19567 32895
rect 19567 32861 19576 32895
rect 19524 32852 19576 32861
rect 20536 32852 20588 32904
rect 27804 32852 27856 32904
rect 32772 32852 32824 32904
rect 38108 32895 38160 32904
rect 38108 32861 38117 32895
rect 38117 32861 38151 32895
rect 38151 32861 38160 32895
rect 38108 32852 38160 32861
rect 9036 32716 9088 32768
rect 18880 32716 18932 32768
rect 19432 32716 19484 32768
rect 36544 32716 36596 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 9772 32512 9824 32564
rect 23112 32512 23164 32564
rect 26332 32512 26384 32564
rect 31484 32512 31536 32564
rect 10416 32444 10468 32496
rect 27804 32444 27856 32496
rect 38108 32487 38160 32496
rect 38108 32453 38117 32487
rect 38117 32453 38151 32487
rect 38151 32453 38160 32487
rect 38108 32444 38160 32453
rect 8024 32376 8076 32428
rect 13728 32376 13780 32428
rect 14372 32419 14424 32428
rect 14372 32385 14406 32419
rect 14406 32385 14424 32419
rect 14372 32376 14424 32385
rect 25320 32376 25372 32428
rect 26240 32376 26292 32428
rect 6920 32283 6972 32292
rect 6920 32249 6929 32283
rect 6929 32249 6963 32283
rect 6963 32249 6972 32283
rect 6920 32240 6972 32249
rect 7472 32215 7524 32224
rect 7472 32181 7481 32215
rect 7481 32181 7515 32215
rect 7515 32181 7524 32215
rect 7472 32172 7524 32181
rect 14832 32172 14884 32224
rect 25320 32215 25372 32224
rect 25320 32181 25329 32215
rect 25329 32181 25363 32215
rect 25363 32181 25372 32215
rect 25320 32172 25372 32181
rect 26332 32172 26384 32224
rect 35348 32376 35400 32428
rect 32772 32351 32824 32360
rect 32772 32317 32781 32351
rect 32781 32317 32815 32351
rect 32815 32317 32824 32351
rect 32772 32308 32824 32317
rect 38016 32172 38068 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 18512 31968 18564 32020
rect 26332 31968 26384 32020
rect 26516 32011 26568 32020
rect 26516 31977 26525 32011
rect 26525 31977 26559 32011
rect 26559 31977 26568 32011
rect 26516 31968 26568 31977
rect 29184 31968 29236 32020
rect 30104 31968 30156 32020
rect 32864 31968 32916 32020
rect 27528 31900 27580 31952
rect 21456 31832 21508 31884
rect 13268 31764 13320 31816
rect 13636 31764 13688 31816
rect 15108 31696 15160 31748
rect 26240 31764 26292 31816
rect 27528 31764 27580 31816
rect 28448 31764 28500 31816
rect 36176 31628 36228 31680
rect 36452 31628 36504 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 35348 31424 35400 31476
rect 36176 31356 36228 31408
rect 33048 31288 33100 31340
rect 35900 31288 35952 31340
rect 36452 31331 36504 31340
rect 36452 31297 36470 31331
rect 36470 31297 36504 31331
rect 36452 31288 36504 31297
rect 38108 31331 38160 31340
rect 38108 31297 38117 31331
rect 38117 31297 38151 31331
rect 38151 31297 38160 31331
rect 38108 31288 38160 31297
rect 17316 31084 17368 31136
rect 22652 31084 22704 31136
rect 33416 31084 33468 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 27068 30923 27120 30932
rect 27068 30889 27077 30923
rect 27077 30889 27111 30923
rect 27111 30889 27120 30923
rect 27068 30880 27120 30889
rect 33048 30923 33100 30932
rect 33048 30889 33057 30923
rect 33057 30889 33091 30923
rect 33091 30889 33100 30923
rect 33048 30880 33100 30889
rect 35900 30880 35952 30932
rect 32864 30855 32916 30864
rect 32864 30821 32873 30855
rect 32873 30821 32907 30855
rect 32907 30821 32916 30855
rect 32864 30812 32916 30821
rect 27528 30744 27580 30796
rect 2688 30608 2740 30660
rect 4896 30676 4948 30728
rect 3148 30540 3200 30592
rect 4068 30540 4120 30592
rect 4896 30583 4948 30592
rect 4896 30549 4905 30583
rect 4905 30549 4939 30583
rect 4939 30549 4948 30583
rect 4896 30540 4948 30549
rect 18788 30608 18840 30660
rect 7472 30540 7524 30592
rect 22284 30583 22336 30592
rect 22284 30549 22293 30583
rect 22293 30549 22327 30583
rect 22327 30549 22336 30583
rect 22284 30540 22336 30549
rect 22744 30608 22796 30660
rect 27160 30608 27212 30660
rect 32588 30651 32640 30660
rect 32588 30617 32597 30651
rect 32597 30617 32631 30651
rect 32631 30617 32640 30651
rect 32588 30608 32640 30617
rect 37924 30540 37976 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4988 30379 5040 30388
rect 4988 30345 4997 30379
rect 4997 30345 5031 30379
rect 5031 30345 5040 30379
rect 4988 30336 5040 30345
rect 3148 30268 3200 30320
rect 1584 30200 1636 30252
rect 4896 30200 4948 30252
rect 5632 30268 5684 30320
rect 6368 30311 6420 30320
rect 6368 30277 6377 30311
rect 6377 30277 6411 30311
rect 6411 30277 6420 30311
rect 6368 30268 6420 30277
rect 11888 30336 11940 30388
rect 22744 30379 22796 30388
rect 8024 30311 8076 30320
rect 8024 30277 8033 30311
rect 8033 30277 8067 30311
rect 8067 30277 8076 30311
rect 8024 30268 8076 30277
rect 11612 30268 11664 30320
rect 12992 30311 13044 30320
rect 4068 30175 4120 30184
rect 4068 30141 4077 30175
rect 4077 30141 4111 30175
rect 4111 30141 4120 30175
rect 4068 30132 4120 30141
rect 6184 30064 6236 30116
rect 3976 30039 4028 30048
rect 3976 30005 3985 30039
rect 3985 30005 4019 30039
rect 4019 30005 4028 30039
rect 3976 29996 4028 30005
rect 4620 29996 4672 30048
rect 11336 30200 11388 30252
rect 12992 30277 13001 30311
rect 13001 30277 13035 30311
rect 13035 30277 13044 30311
rect 12992 30268 13044 30277
rect 14372 30311 14424 30320
rect 14372 30277 14381 30311
rect 14381 30277 14415 30311
rect 14415 30277 14424 30311
rect 14372 30268 14424 30277
rect 11796 30200 11848 30252
rect 15936 30268 15988 30320
rect 11612 30064 11664 30116
rect 11704 30039 11756 30048
rect 11704 30005 11713 30039
rect 11713 30005 11747 30039
rect 11747 30005 11756 30039
rect 11704 29996 11756 30005
rect 11888 30039 11940 30048
rect 11888 30005 11897 30039
rect 11897 30005 11931 30039
rect 11931 30005 11940 30039
rect 14832 30175 14884 30184
rect 14832 30141 14841 30175
rect 14841 30141 14875 30175
rect 14875 30141 14884 30175
rect 14832 30132 14884 30141
rect 11888 29996 11940 30005
rect 15936 29996 15988 30048
rect 19248 30268 19300 30320
rect 18696 30200 18748 30252
rect 19432 30268 19484 30320
rect 22744 30345 22753 30379
rect 22753 30345 22787 30379
rect 22787 30345 22796 30379
rect 22744 30336 22796 30345
rect 24952 30268 25004 30320
rect 26976 30268 27028 30320
rect 32588 30336 32640 30388
rect 32404 30268 32456 30320
rect 32956 30268 33008 30320
rect 33324 30268 33376 30320
rect 22928 30200 22980 30252
rect 32220 30243 32272 30252
rect 32220 30209 32229 30243
rect 32229 30209 32263 30243
rect 32263 30209 32272 30243
rect 32220 30200 32272 30209
rect 33416 30200 33468 30252
rect 19432 30132 19484 30184
rect 22284 30175 22336 30184
rect 22284 30141 22293 30175
rect 22293 30141 22327 30175
rect 22327 30141 22336 30175
rect 22284 30132 22336 30141
rect 32128 30175 32180 30184
rect 32128 30141 32137 30175
rect 32137 30141 32171 30175
rect 32171 30141 32180 30175
rect 32128 30132 32180 30141
rect 18328 30064 18380 30116
rect 30288 30064 30340 30116
rect 16212 29996 16264 30048
rect 18420 29996 18472 30048
rect 19432 29996 19484 30048
rect 22284 29996 22336 30048
rect 30748 29996 30800 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 6920 29792 6972 29844
rect 7472 29792 7524 29844
rect 16212 29792 16264 29844
rect 32864 29792 32916 29844
rect 37924 29835 37976 29844
rect 37924 29801 37933 29835
rect 37933 29801 37967 29835
rect 37967 29801 37976 29835
rect 37924 29792 37976 29801
rect 11520 29724 11572 29776
rect 32312 29724 32364 29776
rect 33876 29724 33928 29776
rect 8024 29588 8076 29640
rect 11796 29656 11848 29708
rect 15292 29656 15344 29708
rect 25596 29656 25648 29708
rect 11704 29588 11756 29640
rect 22284 29588 22336 29640
rect 32128 29656 32180 29708
rect 32220 29631 32272 29640
rect 32220 29597 32229 29631
rect 32229 29597 32263 29631
rect 32263 29597 32272 29631
rect 32220 29588 32272 29597
rect 8668 29520 8720 29572
rect 9588 29520 9640 29572
rect 10140 29520 10192 29572
rect 11336 29563 11388 29572
rect 11336 29529 11345 29563
rect 11345 29529 11379 29563
rect 11379 29529 11388 29563
rect 11336 29520 11388 29529
rect 11612 29520 11664 29572
rect 25228 29563 25280 29572
rect 25228 29529 25237 29563
rect 25237 29529 25271 29563
rect 25271 29529 25280 29563
rect 25228 29520 25280 29529
rect 31392 29520 31444 29572
rect 32404 29631 32456 29640
rect 32404 29597 32413 29631
rect 32413 29597 32447 29631
rect 32447 29597 32456 29631
rect 32404 29588 32456 29597
rect 32588 29588 32640 29640
rect 38108 29631 38160 29640
rect 38108 29597 38117 29631
rect 38117 29597 38151 29631
rect 38151 29597 38160 29631
rect 38108 29588 38160 29597
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9588 29248 9640 29300
rect 22928 29291 22980 29300
rect 22928 29257 22937 29291
rect 22937 29257 22971 29291
rect 22971 29257 22980 29291
rect 22928 29248 22980 29257
rect 11520 29155 11572 29164
rect 11520 29121 11529 29155
rect 11529 29121 11563 29155
rect 11563 29121 11572 29155
rect 11520 29112 11572 29121
rect 11888 29112 11940 29164
rect 16212 29112 16264 29164
rect 25228 29112 25280 29164
rect 30288 29112 30340 29164
rect 8668 29087 8720 29096
rect 8668 29053 8677 29087
rect 8677 29053 8711 29087
rect 8711 29053 8720 29087
rect 8668 29044 8720 29053
rect 13084 29044 13136 29096
rect 11336 28976 11388 29028
rect 31392 28976 31444 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6184 28747 6236 28756
rect 6184 28713 6193 28747
rect 6193 28713 6227 28747
rect 6227 28713 6236 28747
rect 6184 28704 6236 28713
rect 6920 28747 6972 28756
rect 6920 28713 6929 28747
rect 6929 28713 6963 28747
rect 6963 28713 6972 28747
rect 6920 28704 6972 28713
rect 18328 28679 18380 28688
rect 18328 28645 18337 28679
rect 18337 28645 18371 28679
rect 18371 28645 18380 28679
rect 18328 28636 18380 28645
rect 15384 28568 15436 28620
rect 29000 28568 29052 28620
rect 6184 28500 6236 28552
rect 6736 28543 6788 28552
rect 6736 28509 6745 28543
rect 6745 28509 6779 28543
rect 6779 28509 6788 28543
rect 6736 28500 6788 28509
rect 9864 28500 9916 28552
rect 18420 28543 18472 28552
rect 18420 28509 18429 28543
rect 18429 28509 18463 28543
rect 18463 28509 18472 28543
rect 18420 28500 18472 28509
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 25780 28432 25832 28484
rect 29000 28432 29052 28484
rect 30840 28475 30892 28484
rect 30840 28441 30849 28475
rect 30849 28441 30883 28475
rect 30883 28441 30892 28475
rect 30840 28432 30892 28441
rect 35900 28432 35952 28484
rect 18420 28407 18472 28416
rect 17592 28364 17644 28373
rect 18420 28373 18429 28407
rect 18429 28373 18463 28407
rect 18463 28373 18472 28407
rect 18420 28364 18472 28373
rect 26424 28364 26476 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 30840 28160 30892 28212
rect 31392 28092 31444 28144
rect 25228 28024 25280 28076
rect 26148 28067 26200 28076
rect 26148 28033 26157 28067
rect 26157 28033 26191 28067
rect 26191 28033 26200 28067
rect 26148 28024 26200 28033
rect 26240 28067 26292 28076
rect 26240 28033 26249 28067
rect 26249 28033 26283 28067
rect 26283 28033 26292 28067
rect 26424 28067 26476 28076
rect 26240 28024 26292 28033
rect 26424 28033 26433 28067
rect 26433 28033 26467 28067
rect 26467 28033 26476 28067
rect 26424 28024 26476 28033
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 27436 28067 27488 28076
rect 27436 28033 27470 28067
rect 27470 28033 27488 28067
rect 27436 28024 27488 28033
rect 31760 28024 31812 28076
rect 32588 28024 32640 28076
rect 38108 28067 38160 28076
rect 38108 28033 38117 28067
rect 38117 28033 38151 28067
rect 38151 28033 38160 28067
rect 38108 28024 38160 28033
rect 30288 27888 30340 27940
rect 27068 27820 27120 27872
rect 32404 27863 32456 27872
rect 32404 27829 32413 27863
rect 32413 27829 32447 27863
rect 32447 27829 32456 27863
rect 32404 27820 32456 27829
rect 36084 27820 36136 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 27436 27616 27488 27668
rect 3976 27548 4028 27600
rect 4528 27455 4580 27464
rect 4528 27421 4537 27455
rect 4537 27421 4571 27455
rect 4571 27421 4580 27455
rect 4528 27412 4580 27421
rect 6920 27548 6972 27600
rect 10784 27548 10836 27600
rect 13544 27548 13596 27600
rect 18696 27591 18748 27600
rect 18696 27557 18705 27591
rect 18705 27557 18739 27591
rect 18739 27557 18748 27591
rect 18696 27548 18748 27557
rect 26148 27548 26200 27600
rect 37556 27591 37608 27600
rect 37556 27557 37565 27591
rect 37565 27557 37599 27591
rect 37599 27557 37608 27591
rect 37556 27548 37608 27557
rect 31760 27523 31812 27532
rect 31760 27489 31769 27523
rect 31769 27489 31803 27523
rect 31803 27489 31812 27523
rect 31760 27480 31812 27489
rect 5632 27344 5684 27396
rect 5356 27319 5408 27328
rect 5356 27285 5365 27319
rect 5365 27285 5399 27319
rect 5399 27285 5408 27319
rect 5356 27276 5408 27285
rect 8116 27276 8168 27328
rect 14372 27276 14424 27328
rect 15476 27276 15528 27328
rect 18420 27412 18472 27464
rect 26240 27412 26292 27464
rect 27068 27412 27120 27464
rect 30840 27412 30892 27464
rect 32404 27455 32456 27464
rect 31392 27344 31444 27396
rect 30840 27319 30892 27328
rect 30840 27285 30849 27319
rect 30849 27285 30883 27319
rect 30883 27285 30892 27319
rect 30840 27276 30892 27285
rect 32404 27421 32413 27455
rect 32413 27421 32447 27455
rect 32447 27421 32456 27455
rect 32404 27412 32456 27421
rect 35900 27480 35952 27532
rect 35440 27344 35492 27396
rect 32588 27276 32640 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 19340 27072 19392 27124
rect 14372 27004 14424 27056
rect 26240 27004 26292 27056
rect 15844 26936 15896 26988
rect 16856 26936 16908 26988
rect 19984 26936 20036 26988
rect 32588 27072 32640 27124
rect 3884 26868 3936 26920
rect 24676 26868 24728 26920
rect 13084 26732 13136 26784
rect 17224 26800 17276 26852
rect 17592 26800 17644 26852
rect 15844 26775 15896 26784
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 15844 26732 15896 26741
rect 35440 26979 35492 26988
rect 35440 26945 35458 26979
rect 35458 26945 35492 26979
rect 35440 26936 35492 26945
rect 35900 26936 35952 26988
rect 37188 26732 37240 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 15844 26528 15896 26580
rect 30840 26528 30892 26580
rect 5632 26460 5684 26512
rect 5356 26392 5408 26444
rect 4620 26324 4672 26376
rect 3792 26231 3844 26240
rect 3792 26197 3801 26231
rect 3801 26197 3835 26231
rect 3835 26197 3844 26231
rect 3792 26188 3844 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4620 25984 4672 26036
rect 26424 25984 26476 26036
rect 30840 26027 30892 26036
rect 30840 25993 30849 26027
rect 30849 25993 30883 26027
rect 30883 25993 30892 26027
rect 30840 25984 30892 25993
rect 2688 25916 2740 25968
rect 6920 25916 6972 25968
rect 8668 25916 8720 25968
rect 17040 25916 17092 25968
rect 21456 25916 21508 25968
rect 3792 25848 3844 25900
rect 27160 25916 27212 25968
rect 22100 25891 22152 25900
rect 22100 25857 22134 25891
rect 22134 25857 22152 25891
rect 30748 25959 30800 25968
rect 30748 25925 30757 25959
rect 30757 25925 30791 25959
rect 30791 25925 30800 25959
rect 30748 25916 30800 25925
rect 22100 25848 22152 25857
rect 8668 25712 8720 25764
rect 15476 25712 15528 25764
rect 38108 25755 38160 25764
rect 14372 25644 14424 25696
rect 38108 25721 38117 25755
rect 38117 25721 38151 25755
rect 38151 25721 38160 25755
rect 38108 25712 38160 25721
rect 23112 25644 23164 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 6736 25440 6788 25492
rect 13084 25483 13136 25492
rect 13084 25449 13093 25483
rect 13093 25449 13127 25483
rect 13127 25449 13136 25483
rect 13084 25440 13136 25449
rect 22100 25440 22152 25492
rect 6920 25347 6972 25356
rect 6920 25313 6929 25347
rect 6929 25313 6963 25347
rect 6963 25313 6972 25347
rect 6920 25304 6972 25313
rect 20536 25372 20588 25424
rect 22836 25372 22888 25424
rect 7932 25168 7984 25220
rect 14372 25304 14424 25356
rect 15476 25347 15528 25356
rect 15476 25313 15485 25347
rect 15485 25313 15519 25347
rect 15519 25313 15528 25347
rect 15476 25304 15528 25313
rect 11612 25236 11664 25288
rect 23112 25279 23164 25288
rect 11520 25168 11572 25220
rect 12992 25168 13044 25220
rect 23112 25245 23121 25279
rect 23121 25245 23155 25279
rect 23155 25245 23164 25279
rect 23112 25236 23164 25245
rect 30932 25440 30984 25492
rect 31392 25304 31444 25356
rect 23388 25236 23440 25288
rect 36084 25236 36136 25288
rect 22836 25168 22888 25220
rect 25688 25168 25740 25220
rect 26424 25168 26476 25220
rect 29000 25211 29052 25220
rect 9680 25143 9732 25152
rect 9680 25109 9689 25143
rect 9689 25109 9723 25143
rect 9723 25109 9732 25143
rect 9680 25100 9732 25109
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 22192 25100 22244 25152
rect 28172 25143 28224 25152
rect 28172 25109 28181 25143
rect 28181 25109 28215 25143
rect 28215 25109 28224 25143
rect 29000 25177 29009 25211
rect 29009 25177 29043 25211
rect 29043 25177 29052 25211
rect 29000 25168 29052 25177
rect 28172 25100 28224 25109
rect 31300 25100 31352 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7932 24939 7984 24948
rect 7932 24905 7941 24939
rect 7941 24905 7975 24939
rect 7975 24905 7984 24939
rect 7932 24896 7984 24905
rect 12992 24939 13044 24948
rect 12992 24905 13001 24939
rect 13001 24905 13035 24939
rect 13035 24905 13044 24939
rect 12992 24896 13044 24905
rect 9680 24828 9732 24880
rect 12624 24871 12676 24880
rect 12624 24837 12633 24871
rect 12633 24837 12667 24871
rect 12667 24837 12676 24871
rect 12624 24828 12676 24837
rect 10140 24803 10192 24812
rect 10140 24769 10149 24803
rect 10149 24769 10183 24803
rect 10183 24769 10192 24803
rect 10140 24760 10192 24769
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 11612 24760 11664 24812
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 12440 24692 12492 24744
rect 13084 24760 13136 24812
rect 14096 24760 14148 24812
rect 20904 24556 20956 24608
rect 28172 24556 28224 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 12440 24352 12492 24404
rect 20904 24395 20956 24404
rect 20904 24361 20913 24395
rect 20913 24361 20947 24395
rect 20947 24361 20956 24395
rect 20904 24352 20956 24361
rect 25688 24395 25740 24404
rect 25688 24361 25697 24395
rect 25697 24361 25731 24395
rect 25731 24361 25740 24395
rect 25688 24352 25740 24361
rect 14096 24216 14148 24268
rect 11612 24148 11664 24200
rect 18880 24148 18932 24200
rect 19432 24080 19484 24132
rect 23388 24148 23440 24200
rect 26240 24284 26292 24336
rect 29920 24123 29972 24132
rect 12532 24012 12584 24064
rect 25136 24055 25188 24064
rect 25136 24021 25145 24055
rect 25145 24021 25179 24055
rect 25179 24021 25188 24055
rect 25136 24012 25188 24021
rect 29920 24089 29929 24123
rect 29929 24089 29963 24123
rect 29963 24089 29972 24123
rect 29920 24080 29972 24089
rect 31392 24148 31444 24200
rect 30840 24080 30892 24132
rect 33784 24080 33836 24132
rect 38016 24123 38068 24132
rect 38016 24089 38025 24123
rect 38025 24089 38059 24123
rect 38059 24089 38068 24123
rect 38016 24080 38068 24089
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 37740 23851 37792 23860
rect 37740 23817 37749 23851
rect 37749 23817 37783 23851
rect 37783 23817 37792 23851
rect 37740 23808 37792 23817
rect 13544 23740 13596 23792
rect 31392 23783 31444 23792
rect 31392 23749 31401 23783
rect 31401 23749 31435 23783
rect 31435 23749 31444 23783
rect 31392 23740 31444 23749
rect 17592 23715 17644 23724
rect 17592 23681 17626 23715
rect 17626 23681 17644 23715
rect 17592 23672 17644 23681
rect 31852 23672 31904 23724
rect 37556 23672 37608 23724
rect 15936 23468 15988 23520
rect 36636 23604 36688 23656
rect 20996 23536 21048 23588
rect 38844 23536 38896 23588
rect 19432 23511 19484 23520
rect 19432 23477 19441 23511
rect 19441 23477 19475 23511
rect 19475 23477 19484 23511
rect 19432 23468 19484 23477
rect 29920 23468 29972 23520
rect 31852 23468 31904 23520
rect 33968 23468 34020 23520
rect 34520 23468 34572 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 17224 23307 17276 23316
rect 17224 23273 17233 23307
rect 17233 23273 17267 23307
rect 17267 23273 17276 23307
rect 17224 23264 17276 23273
rect 17592 23264 17644 23316
rect 17776 23171 17828 23180
rect 17776 23137 17785 23171
rect 17785 23137 17819 23171
rect 17819 23137 17828 23171
rect 17776 23128 17828 23137
rect 17960 23103 18012 23112
rect 17960 23069 17969 23103
rect 17969 23069 18003 23103
rect 18003 23069 18012 23103
rect 17960 23060 18012 23069
rect 31392 23128 31444 23180
rect 21180 23060 21232 23112
rect 28264 23060 28316 23112
rect 33784 23060 33836 23112
rect 37556 23060 37608 23112
rect 20996 23035 21048 23044
rect 20996 23001 21005 23035
rect 21005 23001 21039 23035
rect 21039 23001 21048 23035
rect 20996 22992 21048 23001
rect 26056 23035 26108 23044
rect 26056 23001 26090 23035
rect 26090 23001 26108 23035
rect 26056 22992 26108 23001
rect 22192 22924 22244 22976
rect 27252 22924 27304 22976
rect 37648 22924 37700 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 10232 22720 10284 22772
rect 20352 22720 20404 22772
rect 26056 22720 26108 22772
rect 33232 22763 33284 22772
rect 33232 22729 33241 22763
rect 33241 22729 33275 22763
rect 33275 22729 33284 22763
rect 33232 22720 33284 22729
rect 37096 22720 37148 22772
rect 38476 22720 38528 22772
rect 20996 22652 21048 22704
rect 22744 22652 22796 22704
rect 25136 22584 25188 22636
rect 32956 22584 33008 22636
rect 22192 22516 22244 22568
rect 27252 22516 27304 22568
rect 33784 22559 33836 22568
rect 33784 22525 33793 22559
rect 33793 22525 33827 22559
rect 33827 22525 33836 22559
rect 33784 22516 33836 22525
rect 35900 22652 35952 22704
rect 36636 22652 36688 22704
rect 37648 22584 37700 22636
rect 20996 22380 21048 22432
rect 26424 22380 26476 22432
rect 32956 22380 33008 22432
rect 36084 22423 36136 22432
rect 36084 22389 36093 22423
rect 36093 22389 36127 22423
rect 36127 22389 36136 22423
rect 36084 22380 36136 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 17960 22040 18012 22092
rect 21180 22083 21232 22092
rect 21180 22049 21189 22083
rect 21189 22049 21223 22083
rect 21223 22049 21232 22083
rect 21180 22040 21232 22049
rect 23388 22040 23440 22092
rect 31392 22108 31444 22160
rect 20996 22015 21048 22024
rect 6368 21904 6420 21956
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 20996 21972 21048 21981
rect 38108 22015 38160 22024
rect 38108 21981 38117 22015
rect 38117 21981 38151 22015
rect 38151 21981 38160 22015
rect 38108 21972 38160 21981
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 29552 21836 29604 21888
rect 37096 21904 37148 21956
rect 30472 21836 30524 21888
rect 37740 21836 37792 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3516 21632 3568 21684
rect 3056 21496 3108 21548
rect 3424 21335 3476 21344
rect 3424 21301 3433 21335
rect 3433 21301 3467 21335
rect 3467 21301 3476 21335
rect 3424 21292 3476 21301
rect 13176 21632 13228 21684
rect 32220 21632 32272 21684
rect 11428 21564 11480 21616
rect 31024 21564 31076 21616
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 23756 21496 23808 21548
rect 7840 21428 7892 21480
rect 27988 21428 28040 21480
rect 25872 21360 25924 21412
rect 6552 21292 6604 21344
rect 9956 21292 10008 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6368 21131 6420 21140
rect 6368 21097 6377 21131
rect 6377 21097 6411 21131
rect 6411 21097 6420 21131
rect 6368 21088 6420 21097
rect 26608 21088 26660 21140
rect 35532 21088 35584 21140
rect 5632 20952 5684 21004
rect 6552 20995 6604 21004
rect 6552 20961 6561 20995
rect 6561 20961 6595 20995
rect 6595 20961 6604 20995
rect 6552 20952 6604 20961
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 36084 20952 36136 21004
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 9956 20748 10008 20800
rect 37096 20884 37148 20936
rect 11060 20816 11112 20868
rect 13084 20748 13136 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 7012 20544 7064 20596
rect 11060 20544 11112 20596
rect 37740 20544 37792 20596
rect 3424 20476 3476 20528
rect 28264 20519 28316 20528
rect 28264 20485 28273 20519
rect 28273 20485 28307 20519
rect 28307 20485 28316 20519
rect 28264 20476 28316 20485
rect 29000 20476 29052 20528
rect 6000 20340 6052 20392
rect 6828 20272 6880 20324
rect 7288 20408 7340 20460
rect 15200 20451 15252 20460
rect 7380 20340 7432 20392
rect 12256 20340 12308 20392
rect 8208 20272 8260 20324
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15844 20408 15896 20460
rect 38108 20451 38160 20460
rect 38108 20417 38117 20451
rect 38117 20417 38151 20451
rect 38151 20417 38160 20451
rect 38108 20408 38160 20417
rect 25044 20272 25096 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6736 20000 6788 20052
rect 6920 20000 6972 20052
rect 4620 19932 4672 19984
rect 17960 20000 18012 20052
rect 23756 20000 23808 20052
rect 13084 19975 13136 19984
rect 13084 19941 13093 19975
rect 13093 19941 13127 19975
rect 13127 19941 13136 19975
rect 13084 19932 13136 19941
rect 9956 19864 10008 19916
rect 3424 19796 3476 19848
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 7380 19796 7432 19848
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 12532 19796 12584 19848
rect 17776 19864 17828 19916
rect 23296 19932 23348 19984
rect 27252 19975 27304 19984
rect 15936 19839 15988 19848
rect 9956 19771 10008 19780
rect 9956 19737 9965 19771
rect 9965 19737 9999 19771
rect 9999 19737 10008 19771
rect 9956 19728 10008 19737
rect 12624 19728 12676 19780
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 19984 19864 20036 19916
rect 25044 19864 25096 19916
rect 26056 19864 26108 19916
rect 27252 19941 27261 19975
rect 27261 19941 27295 19975
rect 27295 19941 27304 19975
rect 27252 19932 27304 19941
rect 23112 19796 23164 19848
rect 30196 19864 30248 19916
rect 27252 19796 27304 19848
rect 27344 19728 27396 19780
rect 33232 19796 33284 19848
rect 8208 19660 8260 19712
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 15476 19703 15528 19712
rect 15476 19669 15485 19703
rect 15485 19669 15519 19703
rect 15519 19669 15528 19703
rect 15476 19660 15528 19669
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 26976 19703 27028 19712
rect 26976 19669 26985 19703
rect 26985 19669 27019 19703
rect 27019 19669 27028 19703
rect 30932 19703 30984 19712
rect 26976 19660 27028 19669
rect 30932 19669 30941 19703
rect 30941 19669 30975 19703
rect 30975 19669 30984 19703
rect 30932 19660 30984 19669
rect 34336 19660 34388 19712
rect 35900 19660 35952 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 12256 19499 12308 19508
rect 12256 19465 12265 19499
rect 12265 19465 12299 19499
rect 12299 19465 12308 19499
rect 12256 19456 12308 19465
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 26148 19456 26200 19508
rect 26976 19456 27028 19508
rect 30196 19499 30248 19508
rect 30196 19465 30205 19499
rect 30205 19465 30239 19499
rect 30239 19465 30248 19499
rect 30196 19456 30248 19465
rect 33232 19456 33284 19508
rect 34336 19499 34388 19508
rect 34336 19465 34345 19499
rect 34345 19465 34379 19499
rect 34379 19465 34388 19499
rect 34336 19456 34388 19465
rect 35900 19456 35952 19508
rect 12532 19388 12584 19440
rect 19892 19431 19944 19440
rect 19892 19397 19901 19431
rect 19901 19397 19935 19431
rect 19935 19397 19944 19431
rect 19892 19388 19944 19397
rect 13084 19320 13136 19372
rect 17776 19320 17828 19372
rect 19800 19363 19852 19372
rect 19800 19329 19809 19363
rect 19809 19329 19843 19363
rect 19843 19329 19852 19363
rect 19800 19320 19852 19329
rect 20996 19320 21048 19372
rect 23756 19388 23808 19440
rect 23112 19320 23164 19372
rect 27252 19388 27304 19440
rect 27344 19431 27396 19440
rect 27344 19397 27353 19431
rect 27353 19397 27387 19431
rect 27387 19397 27396 19431
rect 27344 19388 27396 19397
rect 12624 19295 12676 19304
rect 12624 19261 12633 19295
rect 12633 19261 12667 19295
rect 12667 19261 12676 19295
rect 12624 19252 12676 19261
rect 28264 19252 28316 19304
rect 30932 19320 30984 19372
rect 34704 19388 34756 19440
rect 33232 19320 33284 19372
rect 34796 19320 34848 19372
rect 38844 19320 38896 19372
rect 38568 19252 38620 19304
rect 12808 19184 12860 19236
rect 20168 19227 20220 19236
rect 20168 19193 20177 19227
rect 20177 19193 20211 19227
rect 20211 19193 20220 19227
rect 20168 19184 20220 19193
rect 23204 19184 23256 19236
rect 26148 19184 26200 19236
rect 20260 19116 20312 19168
rect 25688 19116 25740 19168
rect 26240 19116 26292 19168
rect 26516 19116 26568 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19892 18912 19944 18964
rect 23112 18955 23164 18964
rect 23112 18921 23121 18955
rect 23121 18921 23155 18955
rect 23155 18921 23164 18955
rect 23112 18912 23164 18921
rect 34704 18955 34756 18964
rect 34704 18921 34713 18955
rect 34713 18921 34747 18955
rect 34747 18921 34756 18955
rect 34704 18912 34756 18921
rect 5172 18844 5224 18896
rect 24216 18844 24268 18896
rect 26424 18844 26476 18896
rect 5724 18708 5776 18760
rect 18052 18640 18104 18692
rect 18880 18640 18932 18692
rect 19800 18683 19852 18692
rect 3148 18572 3200 18624
rect 19432 18572 19484 18624
rect 19800 18649 19827 18683
rect 19827 18649 19852 18683
rect 19800 18640 19852 18649
rect 19984 18683 20036 18692
rect 19984 18649 19993 18683
rect 19993 18649 20027 18683
rect 20027 18649 20036 18683
rect 19984 18640 20036 18649
rect 22376 18708 22428 18760
rect 23204 18776 23256 18828
rect 26056 18776 26108 18828
rect 23296 18751 23348 18760
rect 23296 18717 23305 18751
rect 23305 18717 23339 18751
rect 23339 18717 23348 18751
rect 23296 18708 23348 18717
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 25596 18640 25648 18692
rect 25688 18640 25740 18692
rect 37372 18844 37424 18896
rect 38108 18751 38160 18760
rect 38108 18717 38117 18751
rect 38117 18717 38151 18751
rect 38151 18717 38160 18751
rect 38108 18708 38160 18717
rect 23480 18615 23532 18624
rect 23480 18581 23489 18615
rect 23489 18581 23523 18615
rect 23523 18581 23532 18615
rect 23480 18572 23532 18581
rect 26240 18615 26292 18624
rect 26240 18581 26249 18615
rect 26249 18581 26283 18615
rect 26283 18581 26292 18615
rect 37924 18615 37976 18624
rect 26240 18572 26292 18581
rect 37924 18581 37933 18615
rect 37933 18581 37967 18615
rect 37967 18581 37976 18615
rect 37924 18572 37976 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3056 18368 3108 18420
rect 17960 18368 18012 18420
rect 21088 18368 21140 18420
rect 37280 18368 37332 18420
rect 3240 18232 3292 18284
rect 17684 18275 17736 18284
rect 17684 18241 17693 18275
rect 17693 18241 17727 18275
rect 17727 18241 17736 18275
rect 17684 18232 17736 18241
rect 18052 18232 18104 18284
rect 4620 18164 4672 18216
rect 3976 18028 4028 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3240 17867 3292 17876
rect 3240 17833 3249 17867
rect 3249 17833 3283 17867
rect 3283 17833 3292 17867
rect 3240 17824 3292 17833
rect 7380 17824 7432 17876
rect 3792 17527 3844 17536
rect 3792 17493 3801 17527
rect 3801 17493 3835 17527
rect 3835 17493 3844 17527
rect 3792 17484 3844 17493
rect 4620 17688 4672 17740
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 7380 17620 7432 17672
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 8484 17620 8536 17672
rect 15200 17824 15252 17876
rect 22376 17867 22428 17876
rect 22376 17833 22385 17867
rect 22385 17833 22419 17867
rect 22419 17833 22428 17867
rect 22376 17824 22428 17833
rect 21548 17756 21600 17808
rect 34612 17824 34664 17876
rect 23480 17663 23532 17672
rect 23480 17629 23498 17663
rect 23498 17629 23532 17663
rect 23480 17620 23532 17629
rect 38108 17663 38160 17672
rect 12900 17552 12952 17604
rect 23388 17552 23440 17604
rect 4896 17484 4948 17536
rect 12440 17484 12492 17536
rect 38108 17629 38117 17663
rect 38117 17629 38151 17663
rect 38151 17629 38160 17663
rect 38108 17620 38160 17629
rect 28264 17484 28316 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8484 17323 8536 17332
rect 8484 17289 8493 17323
rect 8493 17289 8527 17323
rect 8527 17289 8536 17323
rect 8484 17280 8536 17289
rect 7380 17144 7432 17196
rect 12716 17280 12768 17332
rect 13360 17280 13412 17332
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 17684 17212 17736 17264
rect 20444 17280 20496 17332
rect 32128 17212 32180 17264
rect 12440 17144 12492 17153
rect 12808 17144 12860 17196
rect 17776 17144 17828 17196
rect 20536 17144 20588 17196
rect 34244 17212 34296 17264
rect 33692 17144 33744 17196
rect 7012 17076 7064 17128
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 12532 17076 12584 17128
rect 34152 17119 34204 17128
rect 34152 17085 34161 17119
rect 34161 17085 34195 17119
rect 34195 17085 34204 17119
rect 34152 17076 34204 17085
rect 37556 17008 37608 17060
rect 7288 16940 7340 16992
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4620 16736 4672 16788
rect 7748 16736 7800 16788
rect 12808 16736 12860 16788
rect 17776 16600 17828 16652
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 12532 16575 12584 16584
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 12532 16532 12584 16541
rect 14464 16532 14516 16584
rect 15200 16532 15252 16584
rect 17684 16575 17736 16584
rect 31944 16600 31996 16652
rect 17684 16541 17699 16575
rect 17699 16541 17733 16575
rect 17733 16541 17736 16575
rect 17684 16532 17736 16541
rect 31392 16575 31444 16584
rect 31392 16541 31401 16575
rect 31401 16541 31435 16575
rect 31435 16541 31444 16575
rect 31392 16532 31444 16541
rect 7196 16507 7248 16516
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 14740 16464 14792 16516
rect 18788 16464 18840 16516
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 8208 16396 8260 16448
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 17776 16439 17828 16448
rect 17776 16405 17785 16439
rect 17785 16405 17819 16439
rect 17819 16405 17828 16439
rect 17776 16396 17828 16405
rect 37464 16439 37516 16448
rect 37464 16405 37473 16439
rect 37473 16405 37507 16439
rect 37507 16405 37516 16439
rect 37464 16396 37516 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 30380 16192 30432 16244
rect 30564 16192 30616 16244
rect 34152 16192 34204 16244
rect 38016 16192 38068 16244
rect 4896 16124 4948 16176
rect 25504 16124 25556 16176
rect 37464 16124 37516 16176
rect 38752 16124 38804 16176
rect 6828 16056 6880 16108
rect 17776 16056 17828 16108
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 20168 16056 20220 16108
rect 29000 16056 29052 16108
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 3976 15852 4028 15904
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 27252 15852 27304 15904
rect 35348 15988 35400 16040
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3792 15648 3844 15700
rect 12532 15648 12584 15700
rect 20168 15648 20220 15700
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4160 15444 4212 15496
rect 15476 15512 15528 15564
rect 28264 15648 28316 15700
rect 31392 15648 31444 15700
rect 27344 15580 27396 15632
rect 32588 15648 32640 15700
rect 34796 15691 34848 15700
rect 34796 15657 34805 15691
rect 34805 15657 34839 15691
rect 34839 15657 34848 15691
rect 34796 15648 34848 15657
rect 35348 15648 35400 15700
rect 29184 15512 29236 15564
rect 18512 15444 18564 15496
rect 20352 15444 20404 15496
rect 34796 15444 34848 15496
rect 37188 15487 37240 15496
rect 37188 15453 37197 15487
rect 37197 15453 37231 15487
rect 37231 15453 37240 15487
rect 37188 15444 37240 15453
rect 38016 15487 38068 15496
rect 38016 15453 38025 15487
rect 38025 15453 38059 15487
rect 38059 15453 38068 15487
rect 38016 15444 38068 15453
rect 12072 15376 12124 15428
rect 26240 15376 26292 15428
rect 36636 15376 36688 15428
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 31484 15351 31536 15360
rect 31484 15317 31493 15351
rect 31493 15317 31527 15351
rect 31527 15317 31536 15351
rect 31484 15308 31536 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 7564 15104 7616 15156
rect 10600 15104 10652 15156
rect 11520 15104 11572 15156
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 22928 15104 22980 15156
rect 29000 15104 29052 15156
rect 30564 15104 30616 15156
rect 36544 15104 36596 15156
rect 37372 15104 37424 15156
rect 38016 15147 38068 15156
rect 38016 15113 38025 15147
rect 38025 15113 38059 15147
rect 38059 15113 38068 15147
rect 38016 15104 38068 15113
rect 22008 15036 22060 15088
rect 29184 15079 29236 15088
rect 29184 15045 29193 15079
rect 29193 15045 29227 15079
rect 29227 15045 29236 15079
rect 29184 15036 29236 15045
rect 4068 14968 4120 15020
rect 7196 14968 7248 15020
rect 17684 14968 17736 15020
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 24492 14968 24544 15020
rect 38476 14968 38528 15020
rect 7748 14900 7800 14952
rect 11612 14900 11664 14952
rect 24400 14900 24452 14952
rect 17960 14832 18012 14884
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 23756 14807 23808 14816
rect 23756 14773 23765 14807
rect 23765 14773 23799 14807
rect 23799 14773 23808 14807
rect 23756 14764 23808 14773
rect 23940 14764 23992 14816
rect 29460 14875 29512 14884
rect 29460 14841 29469 14875
rect 29469 14841 29503 14875
rect 29503 14841 29512 14875
rect 29460 14832 29512 14841
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 13636 14560 13688 14612
rect 14924 14560 14976 14612
rect 19340 14560 19392 14612
rect 23940 14560 23992 14612
rect 24400 14603 24452 14612
rect 24400 14569 24409 14603
rect 24409 14569 24443 14603
rect 24443 14569 24452 14603
rect 24400 14560 24452 14569
rect 29460 14560 29512 14612
rect 10784 14492 10836 14544
rect 6828 14424 6880 14476
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 20812 14424 20864 14476
rect 22928 14424 22980 14476
rect 22744 14356 22796 14408
rect 23756 14492 23808 14544
rect 24860 14492 24912 14544
rect 37280 14399 37332 14408
rect 37280 14365 37289 14399
rect 37289 14365 37323 14399
rect 37323 14365 37332 14399
rect 37280 14356 37332 14365
rect 37556 14399 37608 14408
rect 37556 14365 37565 14399
rect 37565 14365 37599 14399
rect 37599 14365 37608 14399
rect 37556 14356 37608 14365
rect 14648 14288 14700 14340
rect 16212 14288 16264 14340
rect 25320 14288 25372 14340
rect 7196 14220 7248 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 15568 14016 15620 14068
rect 6920 13948 6972 14000
rect 9956 13948 10008 14000
rect 14188 13991 14240 14000
rect 14188 13957 14197 13991
rect 14197 13957 14231 13991
rect 14231 13957 14240 13991
rect 14188 13948 14240 13957
rect 16120 13948 16172 14000
rect 3792 13880 3844 13932
rect 14464 13880 14516 13932
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 24400 13948 24452 14000
rect 25412 13948 25464 14000
rect 23664 13880 23716 13932
rect 25320 13880 25372 13932
rect 11796 13812 11848 13864
rect 13452 13812 13504 13864
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 17868 13812 17920 13864
rect 18512 13812 18564 13864
rect 37280 14016 37332 14068
rect 37740 14016 37792 14068
rect 26332 13948 26384 14000
rect 31484 13991 31536 14000
rect 31484 13957 31493 13991
rect 31493 13957 31527 13991
rect 31527 13957 31536 13991
rect 31484 13948 31536 13957
rect 38660 13948 38712 14000
rect 37740 13923 37792 13932
rect 37740 13889 37749 13923
rect 37749 13889 37783 13923
rect 37783 13889 37792 13923
rect 37740 13880 37792 13889
rect 13636 13744 13688 13796
rect 14096 13676 14148 13728
rect 15752 13676 15804 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 22560 13472 22612 13524
rect 23664 13472 23716 13524
rect 23756 13336 23808 13388
rect 37556 13268 37608 13320
rect 24124 13200 24176 13252
rect 37740 13200 37792 13252
rect 13084 13132 13136 13184
rect 14648 13132 14700 13184
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7748 12928 7800 12980
rect 13912 12860 13964 12912
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7196 12835 7248 12844
rect 7196 12801 7230 12835
rect 7230 12801 7248 12835
rect 7196 12792 7248 12801
rect 12164 12792 12216 12844
rect 10692 12724 10744 12776
rect 22284 12928 22336 12980
rect 25780 12971 25832 12980
rect 25780 12937 25789 12971
rect 25789 12937 25823 12971
rect 25823 12937 25832 12971
rect 25780 12928 25832 12937
rect 17868 12860 17920 12912
rect 28908 12792 28960 12844
rect 32404 12767 32456 12776
rect 32404 12733 32413 12767
rect 32413 12733 32447 12767
rect 32447 12733 32456 12767
rect 32404 12724 32456 12733
rect 33784 12724 33836 12776
rect 19800 12631 19852 12640
rect 19800 12597 19809 12631
rect 19809 12597 19843 12631
rect 19843 12597 19852 12631
rect 19800 12588 19852 12597
rect 23756 12631 23808 12640
rect 23756 12597 23765 12631
rect 23765 12597 23799 12631
rect 23799 12597 23808 12631
rect 23756 12588 23808 12597
rect 33876 12588 33928 12640
rect 38108 12631 38160 12640
rect 38108 12597 38117 12631
rect 38117 12597 38151 12631
rect 38151 12597 38160 12631
rect 38108 12588 38160 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10232 12427 10284 12436
rect 10232 12393 10241 12427
rect 10241 12393 10275 12427
rect 10275 12393 10284 12427
rect 10232 12384 10284 12393
rect 20720 12384 20772 12436
rect 31024 12384 31076 12436
rect 4712 12316 4764 12368
rect 21824 12316 21876 12368
rect 10232 12180 10284 12232
rect 4620 12112 4672 12164
rect 10324 12112 10376 12164
rect 19432 12155 19484 12164
rect 19432 12121 19441 12155
rect 19441 12121 19475 12155
rect 19475 12121 19484 12155
rect 19432 12112 19484 12121
rect 19800 12112 19852 12164
rect 11336 12044 11388 12096
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 23756 12112 23808 12164
rect 27988 12087 28040 12096
rect 27988 12053 27997 12087
rect 27997 12053 28031 12087
rect 28031 12053 28040 12087
rect 27988 12044 28040 12053
rect 28356 12044 28408 12096
rect 31116 12112 31168 12164
rect 37924 12044 37976 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2780 11840 2832 11892
rect 12440 11840 12492 11892
rect 16580 11840 16632 11892
rect 20076 11840 20128 11892
rect 28908 11840 28960 11892
rect 31116 11883 31168 11892
rect 31116 11849 31125 11883
rect 31125 11849 31159 11883
rect 31159 11849 31168 11883
rect 31116 11840 31168 11849
rect 4804 11772 4856 11824
rect 19432 11772 19484 11824
rect 22468 11815 22520 11824
rect 22468 11781 22477 11815
rect 22477 11781 22511 11815
rect 22511 11781 22520 11815
rect 22468 11772 22520 11781
rect 27988 11772 28040 11824
rect 32404 11772 32456 11824
rect 2412 11704 2464 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 20444 11704 20496 11756
rect 22008 11704 22060 11756
rect 11980 11636 12032 11688
rect 10876 11568 10928 11620
rect 12532 11543 12584 11552
rect 12532 11509 12541 11543
rect 12541 11509 12575 11543
rect 12575 11509 12584 11543
rect 12532 11500 12584 11509
rect 15016 11568 15068 11620
rect 24584 11636 24636 11688
rect 26792 11568 26844 11620
rect 28356 11611 28408 11620
rect 28356 11577 28365 11611
rect 28365 11577 28399 11611
rect 28399 11577 28408 11611
rect 28356 11568 28408 11577
rect 31208 11611 31260 11620
rect 31208 11577 31217 11611
rect 31217 11577 31251 11611
rect 31251 11577 31260 11611
rect 31208 11568 31260 11577
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 28540 11543 28592 11552
rect 28540 11509 28549 11543
rect 28549 11509 28583 11543
rect 28583 11509 28592 11543
rect 28540 11500 28592 11509
rect 32036 11500 32088 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 13728 11296 13780 11348
rect 19432 11296 19484 11348
rect 26792 11296 26844 11348
rect 37924 11339 37976 11348
rect 37924 11305 37933 11339
rect 37933 11305 37967 11339
rect 37967 11305 37976 11339
rect 37924 11296 37976 11305
rect 8760 11228 8812 11280
rect 15016 11228 15068 11280
rect 27804 11228 27856 11280
rect 33600 11228 33652 11280
rect 27988 11203 28040 11212
rect 27988 11169 27997 11203
rect 27997 11169 28031 11203
rect 28031 11169 28040 11203
rect 27988 11160 28040 11169
rect 28448 11203 28500 11212
rect 28448 11169 28457 11203
rect 28457 11169 28491 11203
rect 28491 11169 28500 11203
rect 28448 11160 28500 11169
rect 2044 11092 2096 11144
rect 11152 11092 11204 11144
rect 11980 11092 12032 11144
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 10416 11024 10468 11076
rect 13544 11024 13596 11076
rect 20996 11024 21048 11076
rect 22008 11024 22060 11076
rect 26884 11024 26936 11076
rect 35348 11024 35400 11076
rect 37280 11024 37332 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 27804 10795 27856 10804
rect 27804 10761 27813 10795
rect 27813 10761 27847 10795
rect 27847 10761 27856 10795
rect 27804 10752 27856 10761
rect 35992 10795 36044 10804
rect 35992 10761 36001 10795
rect 36001 10761 36035 10795
rect 36035 10761 36044 10795
rect 35992 10752 36044 10761
rect 37372 10752 37424 10804
rect 5540 10684 5592 10736
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 12532 10616 12584 10668
rect 37280 10659 37332 10668
rect 37280 10625 37289 10659
rect 37289 10625 37323 10659
rect 37323 10625 37332 10659
rect 37280 10616 37332 10625
rect 12992 10412 13044 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 36728 10455 36780 10464
rect 36728 10421 36737 10455
rect 36737 10421 36771 10455
rect 36771 10421 36780 10455
rect 36728 10412 36780 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 7104 10140 7156 10192
rect 15292 10208 15344 10260
rect 17776 10208 17828 10260
rect 17408 10140 17460 10192
rect 27160 10004 27212 10056
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 6000 9979 6052 9988
rect 2780 9936 2832 9945
rect 6000 9945 6009 9979
rect 6009 9945 6043 9979
rect 6043 9945 6052 9979
rect 6000 9936 6052 9945
rect 14280 9936 14332 9988
rect 17040 9936 17092 9988
rect 17500 9936 17552 9988
rect 37004 9936 37056 9988
rect 13820 9868 13872 9920
rect 17132 9911 17184 9920
rect 17132 9877 17141 9911
rect 17141 9877 17175 9911
rect 17175 9877 17184 9911
rect 17132 9868 17184 9877
rect 30748 9868 30800 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 17132 9664 17184 9716
rect 33048 9664 33100 9716
rect 9772 9639 9824 9648
rect 9772 9605 9781 9639
rect 9781 9605 9815 9639
rect 9815 9605 9824 9639
rect 9772 9596 9824 9605
rect 14096 9639 14148 9648
rect 14096 9605 14105 9639
rect 14105 9605 14139 9639
rect 14139 9605 14148 9639
rect 14096 9596 14148 9605
rect 14280 9639 14332 9648
rect 14280 9605 14289 9639
rect 14289 9605 14323 9639
rect 14323 9605 14332 9639
rect 14280 9596 14332 9605
rect 17408 9596 17460 9648
rect 24216 9596 24268 9648
rect 28448 9596 28500 9648
rect 13820 9528 13872 9580
rect 14372 9528 14424 9580
rect 7288 9392 7340 9444
rect 25136 9528 25188 9580
rect 28540 9528 28592 9580
rect 37740 9571 37792 9580
rect 37740 9537 37749 9571
rect 37749 9537 37783 9571
rect 37783 9537 37792 9571
rect 37740 9528 37792 9537
rect 13728 9324 13780 9376
rect 27988 9460 28040 9512
rect 31024 9392 31076 9444
rect 24860 9324 24912 9376
rect 31944 9324 31996 9376
rect 37464 9324 37516 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3700 9120 3752 9172
rect 5356 9120 5408 9172
rect 26148 9120 26200 9172
rect 34520 9120 34572 9172
rect 9772 9052 9824 9104
rect 10600 9052 10652 9104
rect 21548 9095 21600 9104
rect 21548 9061 21557 9095
rect 21557 9061 21591 9095
rect 21591 9061 21600 9095
rect 21548 9052 21600 9061
rect 2872 8848 2924 8900
rect 5172 8848 5224 8900
rect 9128 8848 9180 8900
rect 9588 8848 9640 8900
rect 10416 8916 10468 8968
rect 25044 8984 25096 9036
rect 25596 9027 25648 9036
rect 25596 8993 25605 9027
rect 25605 8993 25639 9027
rect 25639 8993 25648 9027
rect 25596 8984 25648 8993
rect 24032 8916 24084 8968
rect 20628 8891 20680 8900
rect 20628 8857 20637 8891
rect 20637 8857 20671 8891
rect 20671 8857 20680 8891
rect 20628 8848 20680 8857
rect 24860 8848 24912 8900
rect 33048 8916 33100 8968
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 9772 8780 9824 8832
rect 20168 8780 20220 8832
rect 24676 8823 24728 8832
rect 24676 8789 24685 8823
rect 24685 8789 24719 8823
rect 24719 8789 24728 8823
rect 24676 8780 24728 8789
rect 26976 8848 27028 8900
rect 34796 8848 34848 8900
rect 35808 8848 35860 8900
rect 27436 8780 27488 8832
rect 36452 8780 36504 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2780 8576 2832 8628
rect 2964 8508 3016 8560
rect 6460 8508 6512 8560
rect 7288 8551 7340 8560
rect 7288 8517 7297 8551
rect 7297 8517 7331 8551
rect 7331 8517 7340 8551
rect 7288 8508 7340 8517
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 5172 8440 5224 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 2964 8372 3016 8424
rect 10968 8372 11020 8424
rect 12256 8372 12308 8424
rect 12900 8508 12952 8560
rect 20168 8440 20220 8492
rect 18788 8372 18840 8424
rect 20352 8372 20404 8424
rect 17500 8304 17552 8356
rect 19340 8304 19392 8356
rect 20260 8304 20312 8356
rect 20628 8440 20680 8492
rect 23572 8576 23624 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 38292 8576 38344 8628
rect 26884 8508 26936 8560
rect 32128 8508 32180 8560
rect 33324 8508 33376 8560
rect 26700 8440 26752 8492
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 24860 8372 24912 8424
rect 32128 8372 32180 8424
rect 35808 8508 35860 8560
rect 33600 8483 33652 8492
rect 33600 8449 33609 8483
rect 33609 8449 33643 8483
rect 33643 8449 33652 8483
rect 33600 8440 33652 8449
rect 37924 8372 37976 8424
rect 20720 8304 20772 8356
rect 23572 8304 23624 8356
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 37464 8347 37516 8356
rect 37464 8313 37473 8347
rect 37473 8313 37507 8347
rect 37507 8313 37516 8347
rect 37464 8304 37516 8313
rect 11520 8236 11572 8288
rect 23940 8279 23992 8288
rect 23940 8245 23949 8279
rect 23949 8245 23983 8279
rect 23983 8245 23992 8279
rect 23940 8236 23992 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 30104 8075 30156 8084
rect 30104 8041 30113 8075
rect 30113 8041 30147 8075
rect 30147 8041 30156 8075
rect 30104 8032 30156 8041
rect 36176 8032 36228 8084
rect 11796 8007 11848 8016
rect 11796 7973 11805 8007
rect 11805 7973 11839 8007
rect 11839 7973 11848 8007
rect 11796 7964 11848 7973
rect 32220 7896 32272 7948
rect 9864 7828 9916 7880
rect 10968 7828 11020 7880
rect 23940 7828 23992 7880
rect 32404 7871 32456 7880
rect 32404 7837 32413 7871
rect 32413 7837 32447 7871
rect 32447 7837 32456 7871
rect 32404 7828 32456 7837
rect 35716 7828 35768 7880
rect 38108 7871 38160 7880
rect 38108 7837 38117 7871
rect 38117 7837 38151 7871
rect 38151 7837 38160 7871
rect 38108 7828 38160 7837
rect 11428 7803 11480 7812
rect 11428 7769 11437 7803
rect 11437 7769 11471 7803
rect 11471 7769 11480 7803
rect 11428 7760 11480 7769
rect 23204 7760 23256 7812
rect 29000 7760 29052 7812
rect 30012 7803 30064 7812
rect 30012 7769 30021 7803
rect 30021 7769 30055 7803
rect 30055 7769 30064 7803
rect 30012 7760 30064 7769
rect 32128 7760 32180 7812
rect 3056 7692 3108 7744
rect 15016 7692 15068 7744
rect 20628 7692 20680 7744
rect 25964 7692 26016 7744
rect 28356 7692 28408 7744
rect 35532 7735 35584 7744
rect 35532 7701 35541 7735
rect 35541 7701 35575 7735
rect 35575 7701 35584 7735
rect 35532 7692 35584 7701
rect 36544 7735 36596 7744
rect 36544 7701 36553 7735
rect 36553 7701 36587 7735
rect 36587 7701 36596 7735
rect 36544 7692 36596 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 7656 7488 7708 7540
rect 18420 7488 18472 7540
rect 26148 7488 26200 7540
rect 28632 7531 28684 7540
rect 28632 7497 28641 7531
rect 28641 7497 28675 7531
rect 28675 7497 28684 7531
rect 28632 7488 28684 7497
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 6644 7216 6696 7268
rect 12624 7148 12676 7200
rect 14188 7284 14240 7336
rect 16120 7352 16172 7404
rect 26148 7352 26200 7404
rect 20168 7284 20220 7336
rect 26240 7284 26292 7336
rect 38292 7420 38344 7472
rect 37188 7352 37240 7404
rect 29368 7284 29420 7336
rect 36176 7284 36228 7336
rect 14004 7216 14056 7268
rect 14832 7216 14884 7268
rect 19340 7216 19392 7268
rect 20536 7216 20588 7268
rect 21088 7216 21140 7268
rect 26792 7216 26844 7268
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 27804 7148 27856 7200
rect 29000 7216 29052 7268
rect 34336 7148 34388 7200
rect 34612 7191 34664 7200
rect 34612 7157 34621 7191
rect 34621 7157 34655 7191
rect 34655 7157 34664 7191
rect 34612 7148 34664 7157
rect 35900 7148 35952 7200
rect 38108 7148 38160 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 14832 6987 14884 6996
rect 14832 6953 14841 6987
rect 14841 6953 14875 6987
rect 14875 6953 14884 6987
rect 14832 6944 14884 6953
rect 16120 6944 16172 6996
rect 26792 6944 26844 6996
rect 6644 6808 6696 6860
rect 16028 6851 16080 6860
rect 16028 6817 16037 6851
rect 16037 6817 16071 6851
rect 16071 6817 16080 6851
rect 18420 6876 18472 6928
rect 33784 6944 33836 6996
rect 16028 6808 16080 6817
rect 20812 6740 20864 6792
rect 21088 6740 21140 6792
rect 24952 6808 25004 6860
rect 30012 6808 30064 6860
rect 31576 6808 31628 6860
rect 32128 6851 32180 6860
rect 32128 6817 32137 6851
rect 32137 6817 32171 6851
rect 32171 6817 32180 6851
rect 32128 6808 32180 6817
rect 36728 6808 36780 6860
rect 27620 6783 27672 6792
rect 27620 6749 27629 6783
rect 27629 6749 27663 6783
rect 27663 6749 27672 6783
rect 27620 6740 27672 6749
rect 16488 6672 16540 6724
rect 19984 6715 20036 6724
rect 5356 6604 5408 6656
rect 19432 6604 19484 6656
rect 19984 6681 19993 6715
rect 19993 6681 20027 6715
rect 20027 6681 20036 6715
rect 19984 6672 20036 6681
rect 20168 6715 20220 6724
rect 20168 6681 20177 6715
rect 20177 6681 20211 6715
rect 20211 6681 20220 6715
rect 20168 6672 20220 6681
rect 24860 6715 24912 6724
rect 24860 6681 24869 6715
rect 24869 6681 24903 6715
rect 24903 6681 24912 6715
rect 24860 6672 24912 6681
rect 35440 6740 35492 6792
rect 37372 6740 37424 6792
rect 38476 6740 38528 6792
rect 28172 6604 28224 6656
rect 30012 6604 30064 6656
rect 30564 6647 30616 6656
rect 30564 6613 30573 6647
rect 30573 6613 30607 6647
rect 30607 6613 30616 6647
rect 30564 6604 30616 6613
rect 32220 6604 32272 6656
rect 32588 6647 32640 6656
rect 32588 6613 32597 6647
rect 32597 6613 32631 6647
rect 32631 6613 32640 6647
rect 32588 6604 32640 6613
rect 33324 6604 33376 6656
rect 33968 6604 34020 6656
rect 34520 6604 34572 6656
rect 35808 6604 35860 6656
rect 38476 6604 38528 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 25688 6400 25740 6452
rect 37740 6400 37792 6452
rect 2964 6196 3016 6248
rect 5264 6332 5316 6384
rect 15568 6375 15620 6384
rect 15568 6341 15577 6375
rect 15577 6341 15611 6375
rect 15611 6341 15620 6375
rect 15568 6332 15620 6341
rect 16764 6332 16816 6384
rect 15844 6264 15896 6316
rect 16488 6264 16540 6316
rect 15016 6196 15068 6248
rect 1584 6060 1636 6112
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 15016 6103 15068 6112
rect 15016 6069 15025 6103
rect 15025 6069 15059 6103
rect 15059 6069 15068 6103
rect 15016 6060 15068 6069
rect 19340 6332 19392 6384
rect 27620 6332 27672 6384
rect 35532 6332 35584 6384
rect 37832 6375 37884 6384
rect 35624 6264 35676 6316
rect 36176 6264 36228 6316
rect 36728 6264 36780 6316
rect 19156 6196 19208 6248
rect 29828 6196 29880 6248
rect 37832 6341 37841 6375
rect 37841 6341 37875 6375
rect 37875 6341 37884 6375
rect 37832 6332 37884 6341
rect 37372 6264 37424 6316
rect 39580 6264 39632 6316
rect 39856 6196 39908 6248
rect 27252 6128 27304 6180
rect 30104 6128 30156 6180
rect 37280 6128 37332 6180
rect 18696 6060 18748 6112
rect 29644 6103 29696 6112
rect 29644 6069 29653 6103
rect 29653 6069 29687 6103
rect 29687 6069 29696 6103
rect 29644 6060 29696 6069
rect 30472 6103 30524 6112
rect 30472 6069 30481 6103
rect 30481 6069 30515 6103
rect 30515 6069 30524 6103
rect 30472 6060 30524 6069
rect 30932 6103 30984 6112
rect 30932 6069 30941 6103
rect 30941 6069 30975 6103
rect 30975 6069 30984 6103
rect 30932 6060 30984 6069
rect 31392 6060 31444 6112
rect 32864 6103 32916 6112
rect 32864 6069 32873 6103
rect 32873 6069 32907 6103
rect 32907 6069 32916 6103
rect 32864 6060 32916 6069
rect 33508 6060 33560 6112
rect 34060 6060 34112 6112
rect 35992 6060 36044 6112
rect 37740 6103 37792 6112
rect 37740 6069 37749 6103
rect 37749 6069 37783 6103
rect 37783 6069 37792 6103
rect 37740 6060 37792 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4620 5856 4672 5908
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 18696 5856 18748 5908
rect 25044 5856 25096 5908
rect 25412 5856 25464 5908
rect 26516 5856 26568 5908
rect 26700 5856 26752 5908
rect 29828 5856 29880 5908
rect 30656 5899 30708 5908
rect 30656 5865 30665 5899
rect 30665 5865 30699 5899
rect 30699 5865 30708 5899
rect 30656 5856 30708 5865
rect 31668 5856 31720 5908
rect 32680 5856 32732 5908
rect 33784 5856 33836 5908
rect 34796 5856 34848 5908
rect 36084 5856 36136 5908
rect 35532 5788 35584 5840
rect 39304 5788 39356 5840
rect 10968 5720 11020 5772
rect 14280 5720 14332 5772
rect 24768 5720 24820 5772
rect 37740 5720 37792 5772
rect 18880 5652 18932 5704
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 30656 5652 30708 5704
rect 1768 5584 1820 5636
rect 2964 5584 3016 5636
rect 7012 5584 7064 5636
rect 1400 5559 1452 5568
rect 1400 5525 1409 5559
rect 1409 5525 1443 5559
rect 1443 5525 1452 5559
rect 1400 5516 1452 5525
rect 1676 5516 1728 5568
rect 3700 5516 3752 5568
rect 4068 5516 4120 5568
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 24860 5584 24912 5636
rect 34060 5652 34112 5704
rect 35440 5695 35492 5704
rect 35440 5661 35449 5695
rect 35449 5661 35483 5695
rect 35483 5661 35492 5695
rect 35440 5652 35492 5661
rect 36636 5695 36688 5704
rect 36636 5661 36645 5695
rect 36645 5661 36679 5695
rect 36679 5661 36688 5695
rect 36636 5652 36688 5661
rect 37096 5695 37148 5704
rect 37096 5661 37105 5695
rect 37105 5661 37139 5695
rect 37139 5661 37148 5695
rect 37096 5652 37148 5661
rect 35808 5584 35860 5636
rect 38016 5627 38068 5636
rect 38016 5593 38025 5627
rect 38025 5593 38059 5627
rect 38059 5593 38068 5627
rect 38016 5584 38068 5593
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 15660 5559 15712 5568
rect 15660 5525 15669 5559
rect 15669 5525 15703 5559
rect 15703 5525 15712 5559
rect 15660 5516 15712 5525
rect 20076 5516 20128 5568
rect 20904 5516 20956 5568
rect 22192 5516 22244 5568
rect 24584 5559 24636 5568
rect 24584 5525 24593 5559
rect 24593 5525 24627 5559
rect 24627 5525 24636 5559
rect 24584 5516 24636 5525
rect 26792 5516 26844 5568
rect 29736 5516 29788 5568
rect 30656 5516 30708 5568
rect 30932 5516 30984 5568
rect 31116 5516 31168 5568
rect 31852 5516 31904 5568
rect 33232 5516 33284 5568
rect 36084 5516 36136 5568
rect 37556 5516 37608 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 26056 5312 26108 5364
rect 26608 5312 26660 5364
rect 29276 5355 29328 5364
rect 29276 5321 29285 5355
rect 29285 5321 29319 5355
rect 29319 5321 29328 5355
rect 29276 5312 29328 5321
rect 30932 5312 30984 5364
rect 32036 5312 32088 5364
rect 32404 5312 32456 5364
rect 33600 5312 33652 5364
rect 34428 5312 34480 5364
rect 37832 5312 37884 5364
rect 21640 5244 21692 5296
rect 26884 5244 26936 5296
rect 27436 5244 27488 5296
rect 31484 5244 31536 5296
rect 32772 5244 32824 5296
rect 35440 5287 35492 5296
rect 35440 5253 35449 5287
rect 35449 5253 35483 5287
rect 35483 5253 35492 5287
rect 35440 5244 35492 5253
rect 29276 5176 29328 5228
rect 31668 5176 31720 5228
rect 31852 5176 31904 5228
rect 32864 5176 32916 5228
rect 33968 5176 34020 5228
rect 36452 5219 36504 5228
rect 8300 5108 8352 5160
rect 22284 5108 22336 5160
rect 30380 5108 30432 5160
rect 36452 5185 36461 5219
rect 36461 5185 36495 5219
rect 36495 5185 36504 5219
rect 36452 5176 36504 5185
rect 38108 5219 38160 5228
rect 38108 5185 38117 5219
rect 38117 5185 38151 5219
rect 38151 5185 38160 5219
rect 38108 5176 38160 5185
rect 4712 5040 4764 5092
rect 6092 5040 6144 5092
rect 23388 5040 23440 5092
rect 24860 5040 24912 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 2780 4972 2832 5024
rect 3240 4972 3292 5024
rect 3792 5015 3844 5024
rect 3792 4981 3801 5015
rect 3801 4981 3835 5015
rect 3835 4981 3844 5015
rect 3792 4972 3844 4981
rect 4620 4972 4672 5024
rect 5632 4972 5684 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 7748 4972 7800 5024
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 9220 4972 9272 5024
rect 9680 4972 9732 5024
rect 10600 4972 10652 5024
rect 11520 4972 11572 5024
rect 11888 4972 11940 5024
rect 12532 4972 12584 5024
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 14832 5015 14884 5024
rect 14832 4981 14841 5015
rect 14841 4981 14875 5015
rect 14875 4981 14884 5015
rect 14832 4972 14884 4981
rect 15752 5015 15804 5024
rect 15752 4981 15761 5015
rect 15761 4981 15795 5015
rect 15795 4981 15804 5015
rect 15752 4972 15804 4981
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 18972 5015 19024 5024
rect 18972 4981 18981 5015
rect 18981 4981 19015 5015
rect 19015 4981 19024 5015
rect 18972 4972 19024 4981
rect 19340 4972 19392 5024
rect 20444 5015 20496 5024
rect 20444 4981 20453 5015
rect 20453 4981 20487 5015
rect 20487 4981 20496 5015
rect 20444 4972 20496 4981
rect 21180 4972 21232 5024
rect 21456 4972 21508 5024
rect 22468 5015 22520 5024
rect 22468 4981 22477 5015
rect 22477 4981 22511 5015
rect 22511 4981 22520 5015
rect 22468 4972 22520 4981
rect 22652 4972 22704 5024
rect 23756 5015 23808 5024
rect 23756 4981 23765 5015
rect 23765 4981 23799 5015
rect 23799 4981 23808 5015
rect 23756 4972 23808 4981
rect 24400 4972 24452 5024
rect 25044 5015 25096 5024
rect 25044 4981 25053 5015
rect 25053 4981 25087 5015
rect 25087 4981 25096 5015
rect 25044 4972 25096 4981
rect 26608 4972 26660 5024
rect 27528 5015 27580 5024
rect 27528 4981 27537 5015
rect 27537 4981 27571 5015
rect 27571 4981 27580 5015
rect 27528 4972 27580 4981
rect 27988 5015 28040 5024
rect 27988 4981 27997 5015
rect 27997 4981 28031 5015
rect 28031 4981 28040 5015
rect 27988 4972 28040 4981
rect 28724 5015 28776 5024
rect 28724 4981 28733 5015
rect 28733 4981 28767 5015
rect 28767 4981 28776 5015
rect 28724 4972 28776 4981
rect 28816 4972 28868 5024
rect 33508 5040 33560 5092
rect 33784 5040 33836 5092
rect 31944 4972 31996 5024
rect 36820 4972 36872 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 5264 4768 5316 4820
rect 6092 4811 6144 4820
rect 6092 4777 6101 4811
rect 6101 4777 6135 4811
rect 6135 4777 6144 4811
rect 6092 4768 6144 4777
rect 8300 4811 8352 4820
rect 8300 4777 8309 4811
rect 8309 4777 8343 4811
rect 8343 4777 8352 4811
rect 8300 4768 8352 4777
rect 12716 4768 12768 4820
rect 2872 4700 2924 4752
rect 3884 4743 3936 4752
rect 3884 4709 3893 4743
rect 3893 4709 3927 4743
rect 3927 4709 3936 4743
rect 3884 4700 3936 4709
rect 8852 4700 8904 4752
rect 20996 4768 21048 4820
rect 25136 4811 25188 4820
rect 25136 4777 25145 4811
rect 25145 4777 25179 4811
rect 25179 4777 25188 4811
rect 25136 4768 25188 4777
rect 27436 4811 27488 4820
rect 1584 4564 1636 4616
rect 1768 4564 1820 4616
rect 2504 4564 2556 4616
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 8300 4632 8352 4684
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 6920 4564 6972 4616
rect 9128 4564 9180 4616
rect 11060 4564 11112 4616
rect 13084 4632 13136 4684
rect 3976 4428 4028 4480
rect 7656 4496 7708 4548
rect 7748 4496 7800 4548
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 8392 4428 8444 4480
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 12808 4564 12860 4616
rect 13360 4564 13412 4616
rect 13452 4564 13504 4616
rect 14096 4564 14148 4616
rect 26240 4700 26292 4752
rect 22744 4632 22796 4684
rect 25872 4632 25924 4684
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 21456 4564 21508 4616
rect 22192 4607 22244 4616
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 25044 4564 25096 4616
rect 27436 4777 27445 4811
rect 27445 4777 27479 4811
rect 27479 4777 27488 4811
rect 27436 4768 27488 4777
rect 31208 4768 31260 4820
rect 32312 4811 32364 4820
rect 32312 4777 32321 4811
rect 32321 4777 32355 4811
rect 32355 4777 32364 4811
rect 32312 4768 32364 4777
rect 33416 4811 33468 4820
rect 33416 4777 33425 4811
rect 33425 4777 33459 4811
rect 33459 4777 33468 4811
rect 33416 4768 33468 4777
rect 33508 4768 33560 4820
rect 35992 4700 36044 4752
rect 37004 4700 37056 4752
rect 26884 4632 26936 4684
rect 26700 4607 26752 4616
rect 26700 4573 26709 4607
rect 26709 4573 26743 4607
rect 26743 4573 26752 4607
rect 26700 4564 26752 4573
rect 28632 4564 28684 4616
rect 31024 4607 31076 4616
rect 11244 4428 11296 4480
rect 13360 4428 13412 4480
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 15476 4428 15528 4480
rect 16212 4428 16264 4480
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 17592 4471 17644 4480
rect 17592 4437 17601 4471
rect 17601 4437 17635 4471
rect 17635 4437 17644 4471
rect 17592 4428 17644 4437
rect 18052 4428 18104 4480
rect 20168 4428 20220 4480
rect 20536 4428 20588 4480
rect 21548 4428 21600 4480
rect 27344 4496 27396 4548
rect 31024 4573 31033 4607
rect 31033 4573 31067 4607
rect 31067 4573 31076 4607
rect 31024 4564 31076 4573
rect 31116 4564 31168 4616
rect 33692 4564 33744 4616
rect 36084 4607 36136 4616
rect 36084 4573 36093 4607
rect 36093 4573 36127 4607
rect 36127 4573 36136 4607
rect 36084 4564 36136 4573
rect 37188 4564 37240 4616
rect 30564 4496 30616 4548
rect 31576 4496 31628 4548
rect 35164 4539 35216 4548
rect 35164 4505 35173 4539
rect 35173 4505 35207 4539
rect 35207 4505 35216 4539
rect 35164 4496 35216 4505
rect 37372 4539 37424 4548
rect 37372 4505 37381 4539
rect 37381 4505 37415 4539
rect 37415 4505 37424 4539
rect 37372 4496 37424 4505
rect 37924 4496 37976 4548
rect 22376 4471 22428 4480
rect 22376 4437 22385 4471
rect 22385 4437 22419 4471
rect 22419 4437 22428 4471
rect 22376 4428 22428 4437
rect 23020 4428 23072 4480
rect 23848 4471 23900 4480
rect 23848 4437 23857 4471
rect 23857 4437 23891 4471
rect 23891 4437 23900 4471
rect 23848 4428 23900 4437
rect 24676 4471 24728 4480
rect 24676 4437 24685 4471
rect 24685 4437 24719 4471
rect 24719 4437 24728 4471
rect 24676 4428 24728 4437
rect 28264 4428 28316 4480
rect 29276 4428 29328 4480
rect 30380 4428 30432 4480
rect 31484 4428 31536 4480
rect 33784 4428 33836 4480
rect 34152 4471 34204 4480
rect 34152 4437 34161 4471
rect 34161 4437 34195 4471
rect 34195 4437 34204 4471
rect 34152 4428 34204 4437
rect 35992 4428 36044 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3884 4224 3936 4276
rect 5540 4224 5592 4276
rect 7288 4224 7340 4276
rect 20536 4267 20588 4276
rect 20536 4233 20545 4267
rect 20545 4233 20579 4267
rect 20579 4233 20588 4267
rect 20536 4224 20588 4233
rect 21640 4224 21692 4276
rect 22284 4224 22336 4276
rect 24676 4224 24728 4276
rect 29000 4224 29052 4276
rect 32404 4224 32456 4276
rect 4804 4156 4856 4208
rect 572 4088 624 4140
rect 1952 4088 2004 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3148 4088 3200 4140
rect 4068 4088 4120 4140
rect 296 4020 348 4072
rect 1584 4020 1636 4072
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 4988 4088 5040 4140
rect 5448 4088 5500 4140
rect 7196 4156 7248 4208
rect 7656 4156 7708 4208
rect 5724 4088 5776 4140
rect 6368 4088 6420 4140
rect 8576 4088 8628 4140
rect 9036 4088 9088 4140
rect 11888 4131 11940 4140
rect 4804 4020 4856 4072
rect 2412 3995 2464 4004
rect 2412 3961 2421 3995
rect 2421 3961 2455 3995
rect 2455 3961 2464 3995
rect 2412 3952 2464 3961
rect 3608 3952 3660 4004
rect 5080 3995 5132 4004
rect 2872 3884 2924 3936
rect 5080 3961 5089 3995
rect 5089 3961 5123 3995
rect 5123 3961 5132 3995
rect 5080 3952 5132 3961
rect 5172 3952 5224 4004
rect 5448 3952 5500 4004
rect 8392 4020 8444 4072
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 9864 4020 9916 4072
rect 7564 3952 7616 4004
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 11980 4088 12032 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 16120 4088 16172 4140
rect 19800 4156 19852 4208
rect 19156 4088 19208 4140
rect 19340 4131 19392 4140
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 31116 4156 31168 4208
rect 15568 4020 15620 4072
rect 17040 4020 17092 4072
rect 12992 3952 13044 4004
rect 14096 3952 14148 4004
rect 17776 4020 17828 4072
rect 19064 4063 19116 4072
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 17316 3952 17368 4004
rect 21732 4088 21784 4140
rect 22192 4088 22244 4140
rect 23204 4131 23256 4140
rect 19800 4020 19852 4072
rect 7012 3884 7064 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 10784 3884 10836 3936
rect 11428 3884 11480 3936
rect 12164 3884 12216 3936
rect 13728 3884 13780 3936
rect 14740 3884 14792 3936
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17040 3884 17092 3936
rect 18144 3884 18196 3936
rect 20352 4020 20404 4072
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 24768 4088 24820 4140
rect 25596 4020 25648 4072
rect 20628 3952 20680 4004
rect 22928 3952 22980 4004
rect 26056 3995 26108 4004
rect 20536 3884 20588 3936
rect 22008 3884 22060 3936
rect 22836 3884 22888 3936
rect 23664 3884 23716 3936
rect 24676 3884 24728 3936
rect 25320 3884 25372 3936
rect 26056 3961 26065 3995
rect 26065 3961 26099 3995
rect 26099 3961 26108 3995
rect 26056 3952 26108 3961
rect 25688 3884 25740 3936
rect 27528 4088 27580 4140
rect 28172 4088 28224 4140
rect 28816 4088 28868 4140
rect 30288 4131 30340 4140
rect 28080 4020 28132 4072
rect 29276 4020 29328 4072
rect 30288 4097 30297 4131
rect 30297 4097 30331 4131
rect 30331 4097 30340 4131
rect 30288 4088 30340 4097
rect 30564 4088 30616 4140
rect 30748 4088 30800 4140
rect 32220 4156 32272 4208
rect 32772 4156 32824 4208
rect 36268 4156 36320 4208
rect 32128 4131 32180 4140
rect 32128 4097 32137 4131
rect 32137 4097 32171 4131
rect 32171 4097 32180 4131
rect 32128 4088 32180 4097
rect 32312 4088 32364 4140
rect 34152 4088 34204 4140
rect 35532 4088 35584 4140
rect 34428 4020 34480 4072
rect 38384 4088 38436 4140
rect 26700 3952 26752 4004
rect 28172 3952 28224 4004
rect 28356 3952 28408 4004
rect 29184 3952 29236 4004
rect 29552 3952 29604 4004
rect 32220 3952 32272 4004
rect 32404 3952 32456 4004
rect 34336 3952 34388 4004
rect 35624 3952 35676 4004
rect 37096 3952 37148 4004
rect 37372 3952 37424 4004
rect 38200 3952 38252 4004
rect 26976 3927 27028 3936
rect 26976 3893 26985 3927
rect 26985 3893 27019 3927
rect 27019 3893 27028 3927
rect 26976 3884 27028 3893
rect 28540 3884 28592 3936
rect 29000 3884 29052 3936
rect 29828 3884 29880 3936
rect 31852 3884 31904 3936
rect 33784 3884 33836 3936
rect 34244 3884 34296 3936
rect 35348 3884 35400 3936
rect 36728 3884 36780 3936
rect 39028 3884 39080 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4896 3680 4948 3732
rect 2228 3544 2280 3596
rect 1676 3476 1728 3528
rect 3240 3519 3292 3528
rect 848 3408 900 3460
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 3700 3476 3752 3528
rect 4160 3476 4212 3528
rect 4988 3476 5040 3528
rect 5448 3544 5500 3596
rect 6000 3680 6052 3732
rect 11612 3680 11664 3732
rect 12072 3680 12124 3732
rect 14464 3680 14516 3732
rect 17132 3680 17184 3732
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 19800 3680 19852 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 7932 3612 7984 3664
rect 20352 3612 20404 3664
rect 22560 3655 22612 3664
rect 22560 3621 22569 3655
rect 22569 3621 22603 3655
rect 22603 3621 22612 3655
rect 22560 3612 22612 3621
rect 24492 3612 24544 3664
rect 6552 3544 6604 3596
rect 1952 3408 2004 3460
rect 2964 3340 3016 3392
rect 4436 3340 4488 3392
rect 4896 3340 4948 3392
rect 5264 3340 5316 3392
rect 5724 3476 5776 3528
rect 7472 3476 7524 3528
rect 8484 3476 8536 3528
rect 9404 3544 9456 3596
rect 10876 3476 10928 3528
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 6276 3408 6328 3460
rect 6736 3408 6788 3460
rect 7012 3340 7064 3392
rect 7932 3340 7984 3392
rect 11152 3408 11204 3460
rect 12716 3587 12768 3596
rect 12716 3553 12725 3587
rect 12725 3553 12759 3587
rect 12759 3553 12768 3587
rect 12716 3544 12768 3553
rect 14188 3544 14240 3596
rect 15844 3587 15896 3596
rect 13084 3476 13136 3528
rect 14096 3476 14148 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14924 3476 14976 3528
rect 14556 3451 14608 3460
rect 14556 3417 14565 3451
rect 14565 3417 14599 3451
rect 14599 3417 14608 3451
rect 14556 3408 14608 3417
rect 9312 3340 9364 3392
rect 13636 3340 13688 3392
rect 14096 3340 14148 3392
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 16488 3544 16540 3596
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 17776 3544 17828 3596
rect 22284 3544 22336 3596
rect 23020 3544 23072 3596
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 17684 3408 17736 3460
rect 18512 3476 18564 3528
rect 18972 3476 19024 3528
rect 19248 3476 19300 3528
rect 20444 3476 20496 3528
rect 20628 3476 20680 3528
rect 21180 3519 21232 3528
rect 21180 3485 21189 3519
rect 21189 3485 21223 3519
rect 21223 3485 21232 3519
rect 21180 3476 21232 3485
rect 21548 3476 21600 3528
rect 22376 3476 22428 3528
rect 23756 3476 23808 3528
rect 24216 3476 24268 3528
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 17868 3340 17920 3392
rect 20720 3340 20772 3392
rect 24860 3340 24912 3392
rect 25872 3680 25924 3732
rect 27528 3680 27580 3732
rect 29552 3680 29604 3732
rect 31300 3680 31352 3732
rect 28816 3612 28868 3664
rect 29184 3612 29236 3664
rect 30196 3612 30248 3664
rect 32220 3680 32272 3732
rect 34244 3680 34296 3732
rect 25596 3544 25648 3596
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 26792 3476 26844 3528
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 28632 3519 28684 3528
rect 28632 3485 28641 3519
rect 28641 3485 28675 3519
rect 28675 3485 28684 3519
rect 28632 3476 28684 3485
rect 25320 3408 25372 3460
rect 28356 3408 28408 3460
rect 29276 3408 29328 3460
rect 29552 3544 29604 3596
rect 29828 3544 29880 3596
rect 30012 3587 30064 3596
rect 30012 3553 30021 3587
rect 30021 3553 30055 3587
rect 30055 3553 30064 3587
rect 30012 3544 30064 3553
rect 29460 3476 29512 3528
rect 31944 3544 31996 3596
rect 30932 3476 30984 3528
rect 37648 3544 37700 3596
rect 31392 3451 31444 3460
rect 26148 3340 26200 3392
rect 26884 3340 26936 3392
rect 27712 3340 27764 3392
rect 28448 3340 28500 3392
rect 30564 3340 30616 3392
rect 30748 3340 30800 3392
rect 31392 3417 31401 3451
rect 31401 3417 31435 3451
rect 31435 3417 31444 3451
rect 31392 3408 31444 3417
rect 33876 3519 33928 3528
rect 33876 3485 33885 3519
rect 33885 3485 33919 3519
rect 33919 3485 33928 3519
rect 33876 3476 33928 3485
rect 34520 3476 34572 3528
rect 34796 3476 34848 3528
rect 36544 3476 36596 3528
rect 38200 3476 38252 3528
rect 33048 3408 33100 3460
rect 38384 3408 38436 3460
rect 31024 3340 31076 3392
rect 32680 3340 32732 3392
rect 34336 3340 34388 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3516 3136 3568 3188
rect 5724 3136 5776 3188
rect 9312 3136 9364 3188
rect 9588 3179 9640 3188
rect 9588 3145 9597 3179
rect 9597 3145 9631 3179
rect 9631 3145 9640 3179
rect 9588 3136 9640 3145
rect 10508 3136 10560 3188
rect 13544 3136 13596 3188
rect 14372 3136 14424 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 16856 3179 16908 3188
rect 3332 3068 3384 3120
rect 3792 3068 3844 3120
rect 4712 3111 4764 3120
rect 4712 3077 4721 3111
rect 4721 3077 4755 3111
rect 4755 3077 4764 3111
rect 4712 3068 4764 3077
rect 5540 3068 5592 3120
rect 6644 3068 6696 3120
rect 7932 3068 7984 3120
rect 1124 3000 1176 3052
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 2872 2975 2924 2984
rect 112 2796 164 2848
rect 1400 2796 1452 2848
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 3884 3000 3936 3052
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 8024 3000 8076 3052
rect 4896 2932 4948 2984
rect 14096 3068 14148 3120
rect 14280 3068 14332 3120
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 18604 3179 18656 3188
rect 18604 3145 18613 3179
rect 18613 3145 18647 3179
rect 18647 3145 18656 3179
rect 18604 3136 18656 3145
rect 19984 3136 20036 3188
rect 20536 3136 20588 3188
rect 16396 3068 16448 3120
rect 17408 3068 17460 3120
rect 17960 3111 18012 3120
rect 17960 3077 17969 3111
rect 17969 3077 18003 3111
rect 18003 3077 18012 3111
rect 17960 3068 18012 3077
rect 18972 3068 19024 3120
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 9680 3000 9732 3052
rect 9956 3000 10008 3052
rect 10140 3000 10192 3052
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 11336 3000 11388 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 12624 3000 12676 3052
rect 14372 3043 14424 3052
rect 8852 2932 8904 2984
rect 9128 2932 9180 2984
rect 5448 2796 5500 2848
rect 7012 2796 7064 2848
rect 9588 2864 9640 2916
rect 12440 2932 12492 2984
rect 13360 2932 13412 2984
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14648 3000 14700 3052
rect 15016 3000 15068 3052
rect 10784 2864 10836 2916
rect 11336 2864 11388 2916
rect 13268 2864 13320 2916
rect 15752 3000 15804 3052
rect 15936 2932 15988 2984
rect 17224 3000 17276 3052
rect 17684 3000 17736 3052
rect 18052 3000 18104 3052
rect 18328 3000 18380 3052
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 20168 3068 20220 3120
rect 19984 3000 20036 3052
rect 20444 3000 20496 3052
rect 22928 3068 22980 3120
rect 23112 3068 23164 3120
rect 23848 3068 23900 3120
rect 24124 3068 24176 3120
rect 24584 3068 24636 3120
rect 25504 3068 25556 3120
rect 27436 3068 27488 3120
rect 27988 3068 28040 3120
rect 28356 3111 28408 3120
rect 28356 3077 28365 3111
rect 28365 3077 28399 3111
rect 28399 3077 28408 3111
rect 28356 3068 28408 3077
rect 28816 3068 28868 3120
rect 29736 3111 29788 3120
rect 29736 3077 29745 3111
rect 29745 3077 29779 3111
rect 29779 3077 29788 3111
rect 29736 3068 29788 3077
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22652 3043 22704 3052
rect 22100 3000 22152 3009
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 23388 3000 23440 3052
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 25964 3000 26016 3052
rect 28080 3000 28132 3052
rect 28724 3000 28776 3052
rect 29368 3000 29420 3052
rect 30472 3000 30524 3052
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 16764 2932 16816 2984
rect 34428 3068 34480 3120
rect 35440 3068 35492 3120
rect 35716 3111 35768 3120
rect 35716 3077 35725 3111
rect 35725 3077 35759 3111
rect 35759 3077 35768 3111
rect 35716 3068 35768 3077
rect 32404 3000 32456 3052
rect 32588 3000 32640 3052
rect 32956 3000 33008 3052
rect 33784 3043 33836 3052
rect 33784 3009 33793 3043
rect 33793 3009 33827 3043
rect 33827 3009 33836 3043
rect 33784 3000 33836 3009
rect 33324 2932 33376 2984
rect 35532 3000 35584 3052
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 37464 3000 37516 3052
rect 38752 2932 38804 2984
rect 16304 2864 16356 2916
rect 20720 2864 20772 2916
rect 24492 2864 24544 2916
rect 8944 2796 8996 2848
rect 12532 2796 12584 2848
rect 13084 2796 13136 2848
rect 13360 2796 13412 2848
rect 13636 2796 13688 2848
rect 18696 2796 18748 2848
rect 20352 2796 20404 2848
rect 21180 2796 21232 2848
rect 25320 2864 25372 2916
rect 27528 2907 27580 2916
rect 27528 2873 27537 2907
rect 27537 2873 27571 2907
rect 27571 2873 27580 2907
rect 27528 2864 27580 2873
rect 27896 2864 27948 2916
rect 33600 2864 33652 2916
rect 35716 2864 35768 2916
rect 36360 2864 36412 2916
rect 25688 2796 25740 2848
rect 33508 2796 33560 2848
rect 35624 2839 35676 2848
rect 35624 2805 35633 2839
rect 35633 2805 35667 2839
rect 35667 2805 35676 2839
rect 35624 2796 35676 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 9864 2592 9916 2644
rect 10692 2635 10744 2644
rect 10692 2601 10701 2635
rect 10701 2601 10735 2635
rect 10735 2601 10744 2635
rect 10692 2592 10744 2601
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 15108 2635 15160 2644
rect 15108 2601 15117 2635
rect 15117 2601 15151 2635
rect 15151 2601 15160 2635
rect 15108 2592 15160 2601
rect 16948 2592 17000 2644
rect 17500 2592 17552 2644
rect 8760 2524 8812 2576
rect 9128 2524 9180 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 3056 2456 3108 2508
rect 4436 2456 4488 2508
rect 4620 2456 4672 2508
rect 9036 2456 9088 2508
rect 9220 2499 9272 2508
rect 9220 2465 9229 2499
rect 9229 2465 9263 2499
rect 9263 2465 9272 2499
rect 9220 2456 9272 2465
rect 9680 2524 9732 2576
rect 21272 2592 21324 2644
rect 22100 2592 22152 2644
rect 34704 2592 34756 2644
rect 18788 2524 18840 2576
rect 19432 2524 19484 2576
rect 27252 2524 27304 2576
rect 22284 2456 22336 2508
rect 22468 2456 22520 2508
rect 36452 2524 36504 2576
rect 29644 2456 29696 2508
rect 29920 2456 29972 2508
rect 31760 2456 31812 2508
rect 35900 2499 35952 2508
rect 35900 2465 35909 2499
rect 35909 2465 35943 2499
rect 35943 2465 35952 2499
rect 35900 2456 35952 2465
rect 36544 2456 36596 2508
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 38844 2456 38896 2508
rect 2228 2388 2280 2440
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 4988 2388 5040 2440
rect 6460 2388 6512 2440
rect 1400 2320 1452 2372
rect 1768 2320 1820 2372
rect 2964 2320 3016 2372
rect 3976 2320 4028 2372
rect 6092 2320 6144 2372
rect 8116 2388 8168 2440
rect 8852 2388 8904 2440
rect 10232 2388 10284 2440
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 14004 2388 14056 2440
rect 14832 2388 14884 2440
rect 15660 2388 15712 2440
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17316 2388 17368 2440
rect 17592 2388 17644 2440
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 20260 2388 20312 2440
rect 10968 2320 11020 2372
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 8760 2252 8812 2304
rect 14188 2320 14240 2372
rect 18144 2320 18196 2372
rect 18420 2320 18472 2372
rect 19156 2320 19208 2372
rect 23940 2388 23992 2440
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 24768 2320 24820 2372
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 23848 2295 23900 2304
rect 23848 2261 23857 2295
rect 23857 2261 23891 2295
rect 23891 2261 23900 2295
rect 23848 2252 23900 2261
rect 26700 2388 26752 2440
rect 27160 2388 27212 2440
rect 28264 2431 28316 2440
rect 28264 2397 28273 2431
rect 28273 2397 28307 2431
rect 28307 2397 28316 2431
rect 28264 2388 28316 2397
rect 29000 2431 29052 2440
rect 29000 2397 29009 2431
rect 29009 2397 29043 2431
rect 29043 2397 29052 2431
rect 29000 2388 29052 2397
rect 29092 2388 29144 2440
rect 30104 2388 30156 2440
rect 32220 2431 32272 2440
rect 32220 2397 32229 2431
rect 32229 2397 32263 2431
rect 32263 2397 32272 2431
rect 32220 2388 32272 2397
rect 33692 2388 33744 2440
rect 34612 2388 34664 2440
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 37924 2388 37976 2440
rect 26424 2320 26476 2372
rect 27344 2320 27396 2372
rect 28080 2320 28132 2372
rect 28172 2295 28224 2304
rect 28172 2261 28181 2295
rect 28181 2261 28215 2295
rect 28215 2261 28224 2295
rect 28172 2252 28224 2261
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 33968 2295 34020 2304
rect 33968 2261 33977 2295
rect 33977 2261 34011 2295
rect 34011 2261 34020 2295
rect 33968 2252 34020 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 16120 2048 16172 2100
rect 36176 2048 36228 2100
rect 9772 1980 9824 2032
rect 31116 1980 31168 2032
rect 4896 1912 4948 1964
rect 27528 1912 27580 1964
rect 2872 1844 2924 1896
rect 12532 1844 12584 1896
rect 18880 1844 18932 1896
rect 28172 1844 28224 1896
rect 14464 1776 14516 1828
rect 33968 1776 34020 1828
rect 12072 1708 12124 1760
rect 23020 1708 23072 1760
<< metal2 >>
rect 110 39200 166 40000
rect 386 39200 442 40000
rect 754 39200 810 40000
rect 1122 39200 1178 40000
rect 1490 39200 1546 40000
rect 1858 39200 1914 40000
rect 2134 39200 2190 40000
rect 2502 39200 2558 40000
rect 2870 39200 2926 40000
rect 3238 39200 3294 40000
rect 3606 39200 3662 40000
rect 3882 39200 3938 40000
rect 4250 39200 4306 40000
rect 4618 39200 4674 40000
rect 4986 39200 5042 40000
rect 5354 39200 5410 40000
rect 5722 39200 5778 40000
rect 5998 39200 6054 40000
rect 6366 39200 6422 40000
rect 6734 39200 6790 40000
rect 7102 39200 7158 40000
rect 7470 39200 7526 40000
rect 7746 39200 7802 40000
rect 8114 39200 8170 40000
rect 8482 39200 8538 40000
rect 8850 39200 8906 40000
rect 9218 39200 9274 40000
rect 9586 39200 9642 40000
rect 9862 39200 9918 40000
rect 10230 39200 10286 40000
rect 10598 39200 10654 40000
rect 10966 39200 11022 40000
rect 11334 39200 11390 40000
rect 11610 39200 11666 40000
rect 11978 39200 12034 40000
rect 12346 39200 12402 40000
rect 12714 39200 12770 40000
rect 13082 39200 13138 40000
rect 13450 39200 13506 40000
rect 13726 39200 13782 40000
rect 14094 39200 14150 40000
rect 14462 39200 14518 40000
rect 14830 39200 14886 40000
rect 15198 39200 15254 40000
rect 15474 39200 15530 40000
rect 15842 39200 15898 40000
rect 16210 39200 16266 40000
rect 16578 39200 16634 40000
rect 16946 39200 17002 40000
rect 17222 39200 17278 40000
rect 17590 39200 17646 40000
rect 17958 39200 18014 40000
rect 18326 39200 18382 40000
rect 18694 39200 18750 40000
rect 19062 39200 19118 40000
rect 19338 39200 19394 40000
rect 19706 39200 19762 40000
rect 19812 39222 20024 39250
rect 124 36854 152 39200
rect 112 36848 164 36854
rect 112 36790 164 36796
rect 400 36378 428 39200
rect 388 36372 440 36378
rect 388 36314 440 36320
rect 768 35834 796 39200
rect 1136 37262 1164 39200
rect 1124 37256 1176 37262
rect 1124 37198 1176 37204
rect 1504 36582 1532 39200
rect 1584 36848 1636 36854
rect 1584 36790 1636 36796
rect 1492 36576 1544 36582
rect 1492 36518 1544 36524
rect 756 35828 808 35834
rect 756 35770 808 35776
rect 1596 35290 1624 36790
rect 1872 36378 1900 39200
rect 2148 37262 2176 39200
rect 2228 37868 2280 37874
rect 2228 37810 2280 37816
rect 2240 37466 2268 37810
rect 2228 37460 2280 37466
rect 2228 37402 2280 37408
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 2136 37256 2188 37262
rect 2136 37198 2188 37204
rect 1860 36372 1912 36378
rect 1860 36314 1912 36320
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1584 35284 1636 35290
rect 1584 35226 1636 35232
rect 1688 35222 1716 36110
rect 1964 35290 1992 37198
rect 2516 36922 2544 39200
rect 2596 37256 2648 37262
rect 2596 37198 2648 37204
rect 2504 36916 2556 36922
rect 2504 36858 2556 36864
rect 2044 36644 2096 36650
rect 2044 36586 2096 36592
rect 1952 35284 2004 35290
rect 1952 35226 2004 35232
rect 1676 35216 1728 35222
rect 1676 35158 1728 35164
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 30025 1624 30194
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1596 29850 1624 29951
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 2056 11354 2084 36586
rect 2608 34746 2636 37198
rect 2884 36378 2912 39200
rect 3252 37194 3280 39200
rect 3240 37188 3292 37194
rect 3240 37130 3292 37136
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 3068 36854 3096 37062
rect 3620 36922 3648 39200
rect 3700 37324 3752 37330
rect 3700 37266 3752 37272
rect 3608 36916 3660 36922
rect 3608 36858 3660 36864
rect 3056 36848 3108 36854
rect 3056 36790 3108 36796
rect 2964 36780 3016 36786
rect 2964 36722 3016 36728
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 2976 35894 3004 36722
rect 3240 36168 3292 36174
rect 3240 36110 3292 36116
rect 3148 36100 3200 36106
rect 3148 36042 3200 36048
rect 2884 35866 3004 35894
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 2780 34604 2832 34610
rect 2780 34546 2832 34552
rect 2688 30660 2740 30666
rect 2688 30602 2740 30608
rect 2700 25974 2728 30602
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 2792 11898 2820 34546
rect 2884 34542 2912 35866
rect 3160 35834 3188 36042
rect 3148 35828 3200 35834
rect 3148 35770 3200 35776
rect 3252 34610 3280 36110
rect 3516 35692 3568 35698
rect 3516 35634 3568 35640
rect 3240 34604 3292 34610
rect 3240 34546 3292 34552
rect 2872 34536 2924 34542
rect 2872 34478 2924 34484
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2056 11150 2084 11290
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 296 4072 348 4078
rect 296 4014 348 4020
rect 112 2848 164 2854
rect 112 2790 164 2796
rect 124 800 152 2790
rect 308 800 336 4014
rect 584 800 612 4082
rect 848 3460 900 3466
rect 848 3402 900 3408
rect 860 800 888 3402
rect 1412 3058 1440 5510
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1124 3052 1176 3058
rect 1124 2994 1176 3000
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1136 800 1164 2994
rect 1400 2848 1452 2854
rect 1504 2836 1532 4966
rect 1596 4622 1624 6054
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 4078 1624 4558
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1688 3534 1716 5510
rect 1780 4622 1808 5578
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1452 2808 1532 2836
rect 1400 2790 1452 2796
rect 1412 2514 1440 2790
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1412 800 1440 2314
rect 1688 800 1716 3470
rect 1780 2378 1808 4558
rect 1964 4146 1992 4966
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2240 3602 2268 4422
rect 2424 4010 2452 11698
rect 2884 10266 2912 34478
rect 3148 30592 3200 30598
rect 3148 30534 3200 30540
rect 3160 30326 3188 30534
rect 3148 30320 3200 30326
rect 3148 30262 3200 30268
rect 3528 21690 3556 35634
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 18426 3096 21490
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3436 20534 3464 21286
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3436 19854 3464 20470
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3160 10033 3188 18566
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3252 17882 3280 18226
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3146 10024 3202 10033
rect 2780 9988 2832 9994
rect 3146 9959 3202 9968
rect 2780 9930 2832 9936
rect 2792 8634 2820 9930
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2884 8498 2912 8842
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8566 3004 8774
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 7562 3004 8366
rect 3068 7750 3096 8434
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 2976 7534 3096 7562
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 4622 2544 6054
rect 2976 5642 3004 6190
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 1964 800 1992 3402
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 2516 800 2544 4558
rect 2792 2446 2820 4966
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2884 4146 2912 4694
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2976 4026 3004 5578
rect 3068 4078 3096 7534
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2884 3998 3004 4026
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2884 3942 2912 3998
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 2990 2912 3878
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3194 3004 3334
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 3068 2514 3096 4014
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 2780 2440 2832 2446
rect 3160 2394 3188 4082
rect 3252 3534 3280 4966
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3528 3194 3556 11698
rect 3712 9178 3740 37266
rect 3896 36378 3924 39200
rect 4264 37754 4292 39200
rect 4080 37726 4292 37754
rect 4080 37448 4108 37726
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4080 37420 4200 37448
rect 4172 37262 4200 37420
rect 4160 37256 4212 37262
rect 4160 37198 4212 37204
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 3884 36372 3936 36378
rect 3884 36314 3936 36320
rect 4080 35834 4108 37130
rect 4632 36922 4660 39200
rect 4896 37460 4948 37466
rect 4896 37402 4948 37408
rect 4620 36916 4672 36922
rect 4620 36858 4672 36864
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4068 35828 4120 35834
rect 4068 35770 4120 35776
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 3884 34944 3936 34950
rect 4632 34932 4660 36722
rect 4712 36168 4764 36174
rect 4712 36110 4764 36116
rect 4724 35894 4752 36110
rect 4724 35866 4844 35894
rect 4816 34950 4844 35866
rect 4908 35714 4936 37402
rect 5000 36922 5028 39200
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 4988 36916 5040 36922
rect 4988 36858 5040 36864
rect 5092 35834 5120 37198
rect 5276 35894 5304 37266
rect 5368 36938 5396 39200
rect 5736 37346 5764 39200
rect 5736 37318 5856 37346
rect 5724 37256 5776 37262
rect 5724 37198 5776 37204
rect 5368 36910 5672 36938
rect 5644 36786 5672 36910
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 5540 36780 5592 36786
rect 5540 36722 5592 36728
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 5368 36378 5396 36722
rect 5356 36372 5408 36378
rect 5356 36314 5408 36320
rect 5276 35866 5488 35894
rect 5080 35828 5132 35834
rect 5080 35770 5132 35776
rect 4908 35686 5396 35714
rect 5172 35624 5224 35630
rect 5172 35566 5224 35572
rect 4712 34944 4764 34950
rect 4632 34904 4712 34932
rect 3884 34886 3936 34892
rect 4712 34886 4764 34892
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 3896 26926 3924 34886
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 4080 30190 4108 30534
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 3976 30048 4028 30054
rect 3976 29990 4028 29996
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 3988 27606 4016 29990
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 3976 27600 4028 27606
rect 4632 27554 4660 29990
rect 3976 27542 4028 27548
rect 4540 27526 4660 27554
rect 4540 27470 4568 27526
rect 4528 27464 4580 27470
rect 4528 27406 4580 27412
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4632 26382 4660 27526
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3804 25906 3832 26182
rect 4632 26042 4660 26318
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4632 18222 4660 19926
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3988 17678 4016 18022
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4632 17746 4660 18158
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3804 15706 3832 17478
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4632 16794 4660 17682
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3988 15502 4016 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 3976 15496 4028 15502
rect 4160 15496 4212 15502
rect 3976 15438 4028 15444
rect 4080 15444 4160 15450
rect 4080 15438 4212 15444
rect 4080 15422 4200 15438
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 13938 3832 15302
rect 4080 15026 4108 15422
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14074 4108 14962
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4724 12374 4752 34886
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4632 5914 4660 12106
rect 4816 11830 4844 34886
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4908 30734 4936 33254
rect 4896 30728 4948 30734
rect 4948 30676 5028 30682
rect 4896 30670 5028 30676
rect 4908 30654 5028 30670
rect 4896 30592 4948 30598
rect 4896 30534 4948 30540
rect 4908 30258 4936 30534
rect 5000 30394 5028 30654
rect 4988 30388 5040 30394
rect 4988 30330 5040 30336
rect 4896 30252 4948 30258
rect 4896 30194 4948 30200
rect 5184 18902 5212 35566
rect 5264 34604 5316 34610
rect 5264 34546 5316 34552
rect 5276 33658 5304 34546
rect 5264 33652 5316 33658
rect 5264 33594 5316 33600
rect 5368 33538 5396 35686
rect 5276 33510 5396 33538
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 16182 4936 17478
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 2780 2382 2832 2388
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 3068 2366 3188 2394
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 1902 2912 2246
rect 2872 1896 2924 1902
rect 2872 1838 2924 1844
rect 2976 1714 3004 2314
rect 2792 1686 3004 1714
rect 2792 800 2820 1686
rect 3068 800 3096 2366
rect 3344 800 3372 3062
rect 3620 800 3648 3946
rect 3712 3534 3740 5510
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3804 3126 3832 4966
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3896 4282 3924 4694
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3896 800 3924 2994
rect 3988 2378 4016 4422
rect 4080 4146 4108 5510
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4434 3496 4490 3505
rect 4172 2836 4200 3470
rect 4434 3431 4490 3440
rect 4448 3398 4476 3431
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4080 2808 4200 2836
rect 4080 2530 4108 2808
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4080 2502 4200 2530
rect 4632 2514 4660 4966
rect 4724 3126 4752 5034
rect 4816 4214 4844 6054
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4816 2774 4844 4014
rect 4908 3738 4936 10610
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8498 5212 8842
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5000 3534 5028 4082
rect 5078 4040 5134 4049
rect 5184 4010 5212 8434
rect 5276 6390 5304 33510
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5368 26450 5396 27270
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5460 22094 5488 35866
rect 5552 34950 5580 36722
rect 5736 35494 5764 37198
rect 5828 36922 5856 37318
rect 5816 36916 5868 36922
rect 5816 36858 5868 36864
rect 6012 36378 6040 39200
rect 6380 37262 6408 39200
rect 6368 37256 6420 37262
rect 6368 37198 6420 37204
rect 6184 36780 6236 36786
rect 6184 36722 6236 36728
rect 6000 36372 6052 36378
rect 6000 36314 6052 36320
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5540 34944 5592 34950
rect 5540 34886 5592 34892
rect 5368 22066 5488 22094
rect 5368 9178 5396 22066
rect 5552 10742 5580 34886
rect 5632 30320 5684 30326
rect 5632 30262 5684 30268
rect 5644 27402 5672 30262
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 5644 26518 5672 27338
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 5644 21010 5672 26454
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5736 18766 5764 35430
rect 6196 35290 6224 36722
rect 6380 36582 6408 37198
rect 6748 36666 6776 39200
rect 7116 37210 7144 39200
rect 7288 37800 7340 37806
rect 7288 37742 7340 37748
rect 7300 37466 7328 37742
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7484 37262 7512 39200
rect 7472 37256 7524 37262
rect 7116 37182 7236 37210
rect 7472 37198 7524 37204
rect 7104 36780 7156 36786
rect 7104 36722 7156 36728
rect 6748 36650 6960 36666
rect 6644 36644 6696 36650
rect 6748 36644 6972 36650
rect 6748 36638 6920 36644
rect 6644 36586 6696 36592
rect 6920 36586 6972 36592
rect 6368 36576 6420 36582
rect 6368 36518 6420 36524
rect 6460 36100 6512 36106
rect 6460 36042 6512 36048
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 5816 34400 5868 34406
rect 5816 34342 5868 34348
rect 5828 33454 5856 34342
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 6368 33448 6420 33454
rect 6368 33390 6420 33396
rect 6380 30326 6408 33390
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 6184 30116 6236 30122
rect 6184 30058 6236 30064
rect 6196 28762 6224 30058
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6196 28558 6224 28698
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6012 20398 6040 21830
rect 6380 21146 6408 21898
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5078 3975 5080 3984
rect 5132 3975 5134 3984
rect 5172 4004 5224 4010
rect 5080 3946 5132 3952
rect 5172 3946 5224 3952
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5276 3398 5304 4762
rect 5368 4622 5396 6598
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 4908 2990 4936 3334
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4724 2746 4844 2774
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 4172 800 4200 2502
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4448 800 4476 2450
rect 4724 800 4752 2746
rect 4908 1970 4936 2926
rect 5368 2774 5396 4558
rect 5460 4146 5488 6054
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3602 5488 3946
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 2854 5488 3538
rect 5552 3369 5580 4218
rect 5538 3360 5594 3369
rect 5538 3295 5594 3304
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5276 2746 5396 2774
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 5000 800 5028 2382
rect 5276 800 5304 2746
rect 5552 800 5580 3062
rect 5644 3058 5672 4966
rect 5736 4146 5764 5510
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 6012 3738 6040 9930
rect 6472 8566 6500 36042
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21350 6592 21830
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6564 20602 6592 20946
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4826 6132 5034
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6380 4146 6408 5510
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 6274 3496 6330 3505
rect 5736 3194 5764 3470
rect 6274 3431 6276 3440
rect 6328 3431 6330 3440
rect 6276 3402 6328 3408
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5644 2774 5672 2994
rect 5644 2746 5856 2774
rect 5828 800 5856 2746
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6104 800 6132 2314
rect 6380 800 6408 4082
rect 6472 2446 6500 4966
rect 6564 3602 6592 7278
rect 6656 7274 6684 36586
rect 6736 36576 6788 36582
rect 6736 36518 6788 36524
rect 6748 35290 6776 36518
rect 7012 36168 7064 36174
rect 7012 36110 7064 36116
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 7024 34932 7052 36110
rect 7116 35834 7144 36722
rect 7208 36378 7236 37182
rect 7484 36854 7512 37198
rect 7760 36922 7788 39200
rect 7840 37120 7892 37126
rect 7840 37062 7892 37068
rect 7748 36916 7800 36922
rect 7748 36858 7800 36864
rect 7472 36848 7524 36854
rect 7472 36790 7524 36796
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7470 36272 7526 36281
rect 7470 36207 7526 36216
rect 7484 36174 7512 36207
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7104 35828 7156 35834
rect 7104 35770 7156 35776
rect 7484 35290 7512 36110
rect 7748 35488 7800 35494
rect 7748 35430 7800 35436
rect 7472 35284 7524 35290
rect 7472 35226 7524 35232
rect 7104 34944 7156 34950
rect 7024 34904 7104 34932
rect 7104 34886 7156 34892
rect 6920 33516 6972 33522
rect 6920 33458 6972 33464
rect 6932 32298 6960 33458
rect 6920 32292 6972 32298
rect 6920 32234 6972 32240
rect 6920 29844 6972 29850
rect 6920 29786 6972 29792
rect 6932 28762 6960 29786
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6748 25498 6776 28494
rect 6932 27606 6960 28698
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6932 25362 6960 25910
rect 6920 25356 6972 25362
rect 6920 25298 6972 25304
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20058 6776 20878
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6828 20324 6880 20330
rect 6828 20266 6880 20272
rect 6840 20074 6868 20266
rect 6840 20058 6960 20074
rect 6736 20052 6788 20058
rect 6840 20052 6972 20058
rect 6840 20046 6920 20052
rect 6736 19994 6788 20000
rect 6920 19994 6972 20000
rect 7024 19854 7052 20538
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7024 17134 7052 19790
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16114 6868 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6840 14482 6868 16050
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6932 12850 6960 13942
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7116 10198 7144 34886
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 7484 30598 7512 32166
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7484 29850 7512 30534
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7760 22094 7788 35430
rect 7668 22066 7788 22094
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7300 20466 7328 20946
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19854 7420 20334
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7392 17882 7420 19790
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17678 7420 17818
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17202 7420 17614
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 15026 7236 16458
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7300 14414 7328 16934
rect 7576 15162 7604 17070
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 12850 7236 14214
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 8566 7328 9386
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7668 7546 7696 22066
rect 7852 21486 7880 37062
rect 7932 36780 7984 36786
rect 7932 36722 7984 36728
rect 7944 36378 7972 36722
rect 7932 36372 7984 36378
rect 8128 36360 8156 39200
rect 8496 37262 8524 39200
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8864 36922 8892 39200
rect 9232 37618 9260 39200
rect 9232 37590 9352 37618
rect 8852 36916 8904 36922
rect 8852 36858 8904 36864
rect 8576 36780 8628 36786
rect 8576 36722 8628 36728
rect 8300 36372 8352 36378
rect 8128 36332 8300 36360
rect 7932 36314 7984 36320
rect 8300 36314 8352 36320
rect 8024 36168 8076 36174
rect 8024 36110 8076 36116
rect 8036 35894 8064 36110
rect 8036 35866 8156 35894
rect 8128 35494 8156 35866
rect 8588 35834 8616 36722
rect 9220 36168 9272 36174
rect 9220 36110 9272 36116
rect 8576 35828 8628 35834
rect 8576 35770 8628 35776
rect 9036 35692 9088 35698
rect 9036 35634 9088 35640
rect 8116 35488 8168 35494
rect 8116 35430 8168 35436
rect 8024 33312 8076 33318
rect 8024 33254 8076 33260
rect 8036 32434 8064 33254
rect 8024 32428 8076 32434
rect 8024 32370 8076 32376
rect 8036 30326 8064 32370
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 8036 29646 8064 30262
rect 8024 29640 8076 29646
rect 8024 29582 8076 29588
rect 8128 27334 8156 35430
rect 9048 34950 9076 35634
rect 9036 34944 9088 34950
rect 9036 34886 9088 34892
rect 9048 32774 9076 34886
rect 9232 34610 9260 36110
rect 9324 35834 9352 37590
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 9416 36718 9444 37198
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9312 35828 9364 35834
rect 9312 35770 9364 35776
rect 9600 35290 9628 39200
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 9496 34672 9548 34678
rect 9496 34614 9548 34620
rect 9220 34604 9272 34610
rect 9220 34546 9272 34552
rect 9508 33998 9536 34614
rect 9692 34542 9720 36722
rect 9876 36378 9904 39200
rect 10140 37256 10192 37262
rect 10140 37198 10192 37204
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 10152 35290 10180 37198
rect 10244 36378 10272 39200
rect 10612 37262 10640 39200
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 10416 37120 10468 37126
rect 10416 37062 10468 37068
rect 10232 36372 10284 36378
rect 10232 36314 10284 36320
rect 10232 36168 10284 36174
rect 10232 36110 10284 36116
rect 10244 35290 10272 36110
rect 10140 35284 10192 35290
rect 10140 35226 10192 35232
rect 10232 35284 10284 35290
rect 10232 35226 10284 35232
rect 9680 34536 9732 34542
rect 9680 34478 9732 34484
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9496 33992 9548 33998
rect 9496 33934 9548 33940
rect 9036 32768 9088 32774
rect 9036 32710 9088 32716
rect 9508 31754 9536 33934
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9508 31726 9628 31754
rect 9600 29578 9628 31726
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 8680 29102 8708 29514
rect 9600 29306 9628 29514
rect 9588 29300 9640 29306
rect 9588 29242 9640 29248
rect 8668 29096 8720 29102
rect 8668 29038 8720 29044
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8680 25974 8708 29038
rect 8668 25968 8720 25974
rect 8668 25910 8720 25916
rect 8680 25770 8708 25910
rect 8668 25764 8720 25770
rect 8668 25706 8720 25712
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7944 24954 7972 25162
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 9692 24886 9720 25094
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 8220 19718 8248 20266
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8220 17678 8248 19654
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7760 16794 7788 17070
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 8220 16454 8248 17614
rect 8496 17338 8524 17614
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14414 7788 14894
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7760 12986 7788 14350
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6656 6866 6684 7210
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 4622 6960 5510
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6656 3126 6684 4422
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6748 1714 6776 3402
rect 6656 1686 6776 1714
rect 6656 800 6684 1686
rect 6932 800 6960 4558
rect 7024 3942 7052 5578
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7208 4214 7236 4966
rect 7760 4554 7788 4966
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4282 7328 4422
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7668 4214 7696 4490
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 2854 7052 3334
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7208 800 7236 4150
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7472 3528 7524 3534
rect 7576 3505 7604 3946
rect 7472 3470 7524 3476
rect 7562 3496 7618 3505
rect 7484 800 7512 3470
rect 7562 3431 7618 3440
rect 7760 800 7788 4490
rect 7930 4176 7986 4185
rect 7930 4111 7986 4120
rect 7944 3670 7972 4111
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3126 7972 3334
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 8036 3058 8064 5510
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8312 4826 8340 5102
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8036 800 8064 2994
rect 8128 2446 8156 3878
rect 8312 3777 8340 4626
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4078 8432 4422
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8298 3768 8354 3777
rect 8298 3703 8354 3712
rect 8496 3534 8524 4966
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8298 3224 8354 3233
rect 8298 3159 8354 3168
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8312 800 8340 3159
rect 8390 3088 8446 3097
rect 8390 3023 8392 3032
rect 8444 3023 8446 3032
rect 8392 2994 8444 3000
rect 8588 800 8616 4082
rect 8772 2774 8800 11222
rect 9784 9654 9812 32506
rect 9876 28558 9904 34478
rect 10140 33924 10192 33930
rect 10140 33866 10192 33872
rect 10152 33658 10180 33866
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 10428 32502 10456 37062
rect 10980 36922 11008 39200
rect 10968 36916 11020 36922
rect 10968 36858 11020 36864
rect 10692 36780 10744 36786
rect 10692 36722 10744 36728
rect 10704 35834 10732 36722
rect 11348 36378 11376 39200
rect 11624 37194 11652 39200
rect 11612 37188 11664 37194
rect 11612 37130 11664 37136
rect 11992 36922 12020 39200
rect 12256 37732 12308 37738
rect 12256 37674 12308 37680
rect 12268 37466 12296 37674
rect 12256 37460 12308 37466
rect 12256 37402 12308 37408
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 11980 36916 12032 36922
rect 11980 36858 12032 36864
rect 11336 36372 11388 36378
rect 11336 36314 11388 36320
rect 11704 36168 11756 36174
rect 11704 36110 11756 36116
rect 12070 36136 12126 36145
rect 11716 35834 11744 36110
rect 12070 36071 12072 36080
rect 12124 36071 12126 36080
rect 12072 36042 12124 36048
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 10968 35692 11020 35698
rect 10968 35634 11020 35640
rect 11428 35692 11480 35698
rect 11428 35634 11480 35640
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10796 34542 10824 35022
rect 10980 35018 11008 35634
rect 11244 35624 11296 35630
rect 11244 35566 11296 35572
rect 10968 35012 11020 35018
rect 10968 34954 11020 34960
rect 11256 34542 11284 35566
rect 11440 34950 11468 35634
rect 11428 34944 11480 34950
rect 11428 34886 11480 34892
rect 10784 34536 10836 34542
rect 10784 34478 10836 34484
rect 11244 34536 11296 34542
rect 11244 34478 11296 34484
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10520 33318 10548 33390
rect 10508 33312 10560 33318
rect 10508 33254 10560 33260
rect 10416 32496 10468 32502
rect 10416 32438 10468 32444
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 10152 24818 10180 29514
rect 10796 27606 10824 34478
rect 11060 33856 11112 33862
rect 11060 33798 11112 33804
rect 11072 33658 11100 33798
rect 11060 33652 11112 33658
rect 11060 33594 11112 33600
rect 11072 33522 11100 33594
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10784 27600 10836 27606
rect 10784 27542 10836 27548
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 20806 9996 21286
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9968 19922 9996 20742
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 19786 9996 19858
rect 10152 19854 10180 24754
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 9968 14006 9996 19722
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10244 12442 10272 22714
rect 11256 22094 11284 34478
rect 11334 30288 11390 30297
rect 11334 30223 11336 30232
rect 11388 30223 11390 30232
rect 11336 30194 11388 30200
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 11348 29034 11376 29514
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 11440 24698 11468 34886
rect 12084 34746 12112 36042
rect 12176 35290 12204 37198
rect 12360 36360 12388 39200
rect 12728 36854 12756 39200
rect 13096 36922 13124 39200
rect 13176 37664 13228 37670
rect 13176 37606 13228 37612
rect 13188 37398 13216 37606
rect 13176 37392 13228 37398
rect 13176 37334 13228 37340
rect 13176 37188 13228 37194
rect 13176 37130 13228 37136
rect 13084 36916 13136 36922
rect 13084 36858 13136 36864
rect 13188 36854 13216 37130
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 13176 36848 13228 36854
rect 13176 36790 13228 36796
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 12440 36372 12492 36378
rect 12360 36332 12440 36360
rect 12440 36314 12492 36320
rect 12164 35284 12216 35290
rect 12164 35226 12216 35232
rect 12544 35154 12572 36722
rect 12728 35290 12756 36790
rect 13268 36644 13320 36650
rect 13268 36586 13320 36592
rect 12900 36236 12952 36242
rect 12900 36178 12952 36184
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 12532 35148 12584 35154
rect 12532 35090 12584 35096
rect 12912 34746 12940 36178
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 12900 34740 12952 34746
rect 12900 34682 12952 34688
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 11716 30410 11744 33594
rect 11716 30394 11928 30410
rect 11716 30388 11940 30394
rect 11716 30382 11888 30388
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11624 30122 11652 30262
rect 11612 30116 11664 30122
rect 11612 30058 11664 30064
rect 11520 29776 11572 29782
rect 11520 29718 11572 29724
rect 11532 29170 11560 29718
rect 11624 29578 11652 30058
rect 11716 30054 11744 30382
rect 11888 30330 11940 30336
rect 12992 30320 13044 30326
rect 12990 30288 12992 30297
rect 13044 30288 13046 30297
rect 11796 30252 11848 30258
rect 12990 30223 13046 30232
rect 11796 30194 11848 30200
rect 11704 30048 11756 30054
rect 11704 29990 11756 29996
rect 11716 29646 11744 29990
rect 11808 29714 11836 30194
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11704 29640 11756 29646
rect 11704 29582 11756 29588
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11900 29170 11928 29990
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 13096 26790 13124 29038
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13096 25498 13124 26726
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11532 24818 11560 25162
rect 11624 24818 11652 25230
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 13004 24954 13032 25162
rect 12992 24948 13044 24954
rect 12992 24890 13044 24896
rect 12624 24880 12676 24886
rect 12676 24828 12756 24834
rect 12624 24822 12756 24828
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 12532 24812 12584 24818
rect 12636 24806 12756 24822
rect 13096 24818 13124 25434
rect 12532 24754 12584 24760
rect 11440 24670 11560 24698
rect 11256 22066 11468 22094
rect 11440 21622 11468 22066
rect 11428 21616 11480 21622
rect 11428 21558 11480 21564
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20602 11100 20810
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11532 15162 11560 24670
rect 11624 24206 11652 24754
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12452 24410 12480 24686
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 12544 24070 12572 24754
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12268 19514 12296 20334
rect 12544 19854 12572 24006
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12544 19446 12572 19790
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12636 19310 12664 19722
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12636 17626 12664 19246
rect 12544 17598 12664 17626
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 17202 12480 17478
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12544 17134 12572 17598
rect 12728 17338 12756 24806
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13188 21690 13216 34954
rect 13280 31822 13308 36586
rect 13464 36378 13492 39200
rect 13740 37244 13768 39200
rect 13820 37256 13872 37262
rect 13740 37216 13820 37244
rect 13820 37198 13872 37204
rect 14004 37120 14056 37126
rect 14004 37062 14056 37068
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13452 36168 13504 36174
rect 13452 36110 13504 36116
rect 13912 36168 13964 36174
rect 13912 36110 13964 36116
rect 13360 35556 13412 35562
rect 13360 35498 13412 35504
rect 13268 31816 13320 31822
rect 13268 31758 13320 31764
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13096 19990 13124 20742
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12820 19242 12848 19654
rect 13096 19378 13124 19926
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12820 17202 12848 19178
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16590 12296 16934
rect 12544 16590 12572 17070
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 15434 12112 16390
rect 12544 15706 12572 16526
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10244 12238 10272 12378
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9784 9110 9812 9590
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8864 2990 8892 4694
rect 9048 4146 9076 4966
rect 9140 4622 9168 8842
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8956 3641 8984 4014
rect 8942 3632 8998 3641
rect 8942 3567 8998 3576
rect 9140 3074 9168 4558
rect 9048 3046 9168 3074
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8772 2746 8892 2774
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8772 2310 8800 2518
rect 8864 2446 8892 2746
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8956 1442 8984 2790
rect 9048 2514 9076 3046
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9140 2582 9168 2926
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9232 2514 9260 4966
rect 9416 3602 9444 5510
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3194 9352 3334
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9232 2394 9260 2450
rect 8864 1414 8984 1442
rect 9140 2366 9260 2394
rect 8864 800 8892 1414
rect 9140 800 9168 2366
rect 9416 800 9444 3538
rect 9600 3194 9628 8842
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8498 9812 8774
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9692 3058 9720 4966
rect 9876 4078 9904 7822
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9600 2922 9812 2938
rect 9588 2916 9812 2922
rect 9640 2910 9812 2916
rect 9588 2858 9640 2864
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9692 800 9720 2518
rect 9784 2038 9812 2910
rect 9876 2650 9904 4014
rect 10152 3058 10180 4422
rect 10336 3058 10364 12106
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 8974 10456 11018
rect 10612 9110 10640 15098
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9968 800 9996 2994
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10244 800 10272 2382
rect 10520 800 10548 3130
rect 10612 2446 10640 4966
rect 10704 2650 10732 12718
rect 10796 3942 10824 14486
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10888 3534 10916 11562
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 7886 11008 8366
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10796 800 10824 2858
rect 10980 2378 11008 5714
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 4622 11100 5510
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11072 800 11100 4558
rect 11164 3466 11192 11086
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 3534 11284 4422
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11348 3058 11376 12038
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11428 7812 11480 7818
rect 11428 7754 11480 7760
rect 11440 3942 11468 7754
rect 11532 7410 11560 8230
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11532 3233 11560 4966
rect 11624 3738 11652 14894
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11808 8022 11836 13806
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12176 12434 12204 12786
rect 12084 12406 12204 12434
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11992 11150 12020 11630
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4146 11928 4966
rect 11888 4140 11940 4146
rect 11716 4100 11888 4128
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11518 3224 11574 3233
rect 11518 3159 11574 3168
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11348 800 11376 2858
rect 11716 2774 11744 4100
rect 11888 4082 11940 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11992 3482 12020 4082
rect 12084 3738 12112 12406
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11624 2746 11744 2774
rect 11900 3454 12020 3482
rect 11624 800 11652 2746
rect 11900 800 11928 3454
rect 11978 3224 12034 3233
rect 11978 3159 12034 3168
rect 11992 2446 12020 3159
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12084 1766 12112 2246
rect 12072 1760 12124 1766
rect 12072 1702 12124 1708
rect 12176 800 12204 3878
rect 12268 3058 12296 8366
rect 12452 4026 12480 11834
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 10674 12572 11494
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12912 8566 12940 17546
rect 13372 17338 13400 35498
rect 13464 35494 13492 36110
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13464 13870 13492 35430
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 13556 32178 13584 34682
rect 13924 34610 13952 36110
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 13728 34536 13780 34542
rect 13728 34478 13780 34484
rect 13740 33862 13768 34478
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13740 32434 13768 33798
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13556 32150 13768 32178
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 13556 23798 13584 27542
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13648 14618 13676 31758
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13648 13802 13676 14554
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4146 12572 4966
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12452 3998 12572 4026
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12544 2938 12572 3998
rect 12636 3058 12664 7142
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 4826 12756 5510
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12714 3768 12770 3777
rect 12714 3703 12770 3712
rect 12728 3602 12756 3703
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12452 800 12480 2926
rect 12544 2910 12664 2938
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12544 1902 12572 2790
rect 12636 2446 12664 2910
rect 12820 2774 12848 4558
rect 13004 4146 13032 10406
rect 13096 4690 13124 13126
rect 13740 11354 13768 32150
rect 13924 12918 13952 34546
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 12728 2746 12848 2774
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12532 1896 12584 1902
rect 12532 1838 12584 1844
rect 12728 800 12756 2746
rect 13004 800 13032 3946
rect 13096 3534 13124 4626
rect 13372 4622 13400 4966
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13096 2854 13124 3470
rect 13372 2990 13400 4422
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13280 800 13308 2858
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13372 2650 13400 2790
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13464 800 13492 4558
rect 13556 3194 13584 11018
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9586 13860 9862
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 4146 13768 9318
rect 14016 7274 14044 37062
rect 14108 36922 14136 39200
rect 14096 36916 14148 36922
rect 14096 36858 14148 36864
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 14200 34610 14228 36110
rect 14292 35834 14320 36722
rect 14476 36378 14504 39200
rect 14844 37262 14872 39200
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 14832 36712 14884 36718
rect 14832 36654 14884 36660
rect 14924 36712 14976 36718
rect 14924 36654 14976 36660
rect 14464 36372 14516 36378
rect 14464 36314 14516 36320
rect 14844 35834 14872 36654
rect 14936 36310 14964 36654
rect 15120 36310 15148 37198
rect 15212 36922 15240 39200
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 14924 36304 14976 36310
rect 14924 36246 14976 36252
rect 15108 36304 15160 36310
rect 15108 36246 15160 36252
rect 15488 35834 15516 39200
rect 15856 37448 15884 39200
rect 15856 37420 15976 37448
rect 15844 37324 15896 37330
rect 15844 37266 15896 37272
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14832 35828 14884 35834
rect 14832 35770 14884 35776
rect 15476 35828 15528 35834
rect 15476 35770 15528 35776
rect 14464 35692 14516 35698
rect 14464 35634 14516 35640
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 14476 34950 14504 35634
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24818 14136 25094
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14108 24274 14136 24754
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14200 14006 14228 34546
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14384 30326 14412 32370
rect 14372 30320 14424 30326
rect 14372 30262 14424 30268
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14384 27062 14412 27270
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14372 25696 14424 25702
rect 14372 25638 14424 25644
rect 14384 25362 14412 25638
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14476 16590 14504 34886
rect 14936 34610 14964 35634
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 15752 35080 15804 35086
rect 15752 35022 15804 35028
rect 15120 34746 15148 35022
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 14844 30190 14872 32166
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14660 14346 14688 14758
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 9654 14136 13670
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9654 14320 9930
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3233 13676 3334
rect 13634 3224 13690 3233
rect 13544 3188 13596 3194
rect 13634 3159 13690 3168
rect 13544 3130 13596 3136
rect 13648 2854 13676 3159
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13740 800 13768 3878
rect 14016 2446 14044 4966
rect 14108 4622 14136 5510
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14108 3534 14136 3946
rect 14200 3602 14228 7278
rect 14292 5778 14320 9590
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14384 3720 14412 9522
rect 14476 3738 14504 13874
rect 14660 13870 14688 14282
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14660 13190 14688 13806
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14752 12434 14780 16458
rect 14936 14618 14964 34546
rect 15108 31748 15160 31754
rect 15108 31690 15160 31696
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14568 12406 14780 12434
rect 14292 3692 14412 3720
rect 14464 3732 14516 3738
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3126 14136 3334
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14016 800 14044 2382
rect 14200 2378 14228 3538
rect 14292 3126 14320 3692
rect 14464 3674 14516 3680
rect 14568 3618 14596 12406
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15028 11286 15056 11562
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 7002 14872 7210
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 15028 6254 15056 7686
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14384 3590 14596 3618
rect 14384 3194 14412 3590
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14554 3496 14610 3505
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14278 2408 14334 2417
rect 14188 2372 14240 2378
rect 14278 2343 14334 2352
rect 14188 2314 14240 2320
rect 14292 2310 14320 2343
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14384 2122 14412 2994
rect 14292 2094 14412 2122
rect 14292 800 14320 2094
rect 14476 1834 14504 3470
rect 14554 3431 14556 3440
rect 14608 3431 14610 3440
rect 14556 3402 14608 3408
rect 14660 3058 14688 5510
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14752 2774 14780 3878
rect 14568 2746 14780 2774
rect 14464 1828 14516 1834
rect 14464 1770 14516 1776
rect 14568 800 14596 2746
rect 14844 2446 14872 4966
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 3534 14964 4422
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 15028 3058 15056 6054
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15028 2530 15056 2994
rect 15120 2650 15148 31690
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15212 17882 15240 20402
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 7410 15240 16526
rect 15304 10266 15332 29650
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15396 3194 15424 28562
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15488 25770 15516 27270
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 15488 25362 15516 25706
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15488 15570 15516 19654
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15580 6390 15608 14010
rect 15764 13734 15792 35022
rect 15856 31754 15884 37266
rect 15948 37262 15976 37420
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 15948 35834 15976 36722
rect 16224 36378 16252 39200
rect 16592 36378 16620 39200
rect 16960 36854 16988 39200
rect 17236 36922 17264 39200
rect 17408 37324 17460 37330
rect 17408 37266 17460 37272
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 16948 36848 17000 36854
rect 16948 36790 17000 36796
rect 16212 36372 16264 36378
rect 16212 36314 16264 36320
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 15936 35828 15988 35834
rect 15936 35770 15988 35776
rect 16120 35692 16172 35698
rect 16120 35634 16172 35640
rect 16132 33862 16160 35634
rect 16500 35562 16528 36110
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16580 35624 16632 35630
rect 16580 35566 16632 35572
rect 16488 35556 16540 35562
rect 16488 35498 16540 35504
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 15856 31726 16068 31754
rect 15936 30320 15988 30326
rect 15936 30262 15988 30268
rect 15948 30054 15976 30262
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15856 26790 15884 26930
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15856 26586 15884 26726
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15856 20466 15884 26522
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15948 19854 15976 23462
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 16040 6866 16068 31726
rect 16132 14006 16160 33798
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16224 29850 16252 29990
rect 16212 29844 16264 29850
rect 16212 29786 16264 29792
rect 16224 29170 16252 29786
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 7206 16160 7346
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 7002 16160 7142
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15028 2502 15148 2530
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14844 800 14872 2382
rect 15120 800 15148 2502
rect 15488 2258 15516 4422
rect 15580 4078 15608 6326
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15672 2446 15700 5510
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15764 3058 15792 4966
rect 15856 3602 15884 6258
rect 16224 5914 16252 14282
rect 16592 11898 16620 35566
rect 16776 34950 16804 35634
rect 16764 34944 16816 34950
rect 16764 34886 16816 34892
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16500 6322 16528 6666
rect 16776 6390 16804 34886
rect 16960 34746 16988 36790
rect 17316 36644 17368 36650
rect 17316 36586 17368 36592
rect 17132 36168 17184 36174
rect 17132 36110 17184 36116
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 17144 33862 17172 36110
rect 17224 35216 17276 35222
rect 17224 35158 17276 35164
rect 17236 35086 17264 35158
rect 17224 35080 17276 35086
rect 17224 35022 17276 35028
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16224 4570 16252 5850
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16132 4542 16252 4570
rect 16132 4146 16160 4542
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 16132 3534 16160 3878
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16028 3392 16080 3398
rect 16026 3360 16028 3369
rect 16080 3360 16082 3369
rect 16026 3295 16082 3304
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15396 2230 15516 2258
rect 15396 800 15424 2230
rect 15672 800 15700 2382
rect 15948 800 15976 2926
rect 16132 2106 16160 3470
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 16224 800 16252 4422
rect 16394 4040 16450 4049
rect 16394 3975 16450 3984
rect 16302 3632 16358 3641
rect 16302 3567 16358 3576
rect 16316 2922 16344 3567
rect 16408 3126 16436 3975
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16396 3120 16448 3126
rect 16500 3097 16528 3538
rect 16396 3062 16448 3068
rect 16486 3088 16542 3097
rect 16486 3023 16542 3032
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16684 2446 16712 4966
rect 16868 3194 16896 26930
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 17052 12434 17080 25910
rect 17144 15162 17172 33798
rect 17328 31142 17356 36586
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17236 23322 17264 26794
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 16960 12406 17080 12434
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16672 2440 16724 2446
rect 16500 2400 16672 2428
rect 16500 800 16528 2400
rect 16672 2382 16724 2388
rect 16776 800 16804 2926
rect 16960 2650 16988 12406
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 17052 4486 17080 9930
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17144 9722 17172 9862
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17236 5114 17264 13874
rect 17420 10198 17448 37266
rect 17500 37256 17552 37262
rect 17500 37198 17552 37204
rect 17512 35290 17540 37198
rect 17604 36378 17632 39200
rect 17972 37262 18000 39200
rect 17960 37256 18012 37262
rect 17960 37198 18012 37204
rect 17592 36372 17644 36378
rect 17592 36314 17644 36320
rect 17868 35692 17920 35698
rect 17868 35634 17920 35640
rect 17880 35494 17908 35634
rect 17868 35488 17920 35494
rect 17868 35430 17920 35436
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17604 26858 17632 28358
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17604 23322 17632 23666
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17788 19922 17816 23122
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17696 17270 17724 18226
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17696 16590 17724 17206
rect 17788 17202 17816 19314
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 16658 17816 17138
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17788 16114 17816 16390
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17420 9654 17448 10134
rect 17512 9994 17540 10406
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17144 5086 17264 5114
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17052 4078 17080 4422
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17052 800 17080 3878
rect 17144 3738 17172 5086
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17236 3058 17264 4966
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17328 3534 17356 3946
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 3126 17448 3334
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17512 2650 17540 8298
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17604 2446 17632 4422
rect 17696 3466 17724 14962
rect 17880 13954 17908 35430
rect 17972 35290 18000 37198
rect 18052 37188 18104 37194
rect 18052 37130 18104 37136
rect 18064 36174 18092 37130
rect 18340 36922 18368 39200
rect 18328 36916 18380 36922
rect 18328 36858 18380 36864
rect 18604 36644 18656 36650
rect 18604 36586 18656 36592
rect 18052 36168 18104 36174
rect 18052 36110 18104 36116
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18064 34202 18092 36110
rect 18616 35290 18644 36586
rect 18708 36378 18736 39200
rect 19076 37262 19104 39200
rect 19064 37256 19116 37262
rect 19064 37198 19116 37204
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 18696 36372 18748 36378
rect 18696 36314 18748 36320
rect 18604 35284 18656 35290
rect 18604 35226 18656 35232
rect 18800 35222 18828 36722
rect 19076 35290 19104 37198
rect 19352 36922 19380 39200
rect 19720 39114 19748 39200
rect 19812 39114 19840 39222
rect 19720 39086 19840 39114
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 18788 35216 18840 35222
rect 18788 35158 18840 35164
rect 18420 35148 18472 35154
rect 18604 35148 18656 35154
rect 18472 35108 18604 35136
rect 18420 35090 18472 35096
rect 18604 35090 18656 35096
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 18340 33658 18368 34546
rect 19444 34490 19472 37062
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36922 20024 39222
rect 20074 39200 20130 40000
rect 20442 39200 20498 40000
rect 20810 39200 20866 40000
rect 21086 39200 21142 40000
rect 21454 39200 21510 40000
rect 21822 39200 21878 40000
rect 22190 39200 22246 40000
rect 22558 39200 22614 40000
rect 22926 39200 22982 40000
rect 23202 39200 23258 40000
rect 23570 39200 23626 40000
rect 23938 39200 23994 40000
rect 24306 39200 24362 40000
rect 24674 39200 24730 40000
rect 24950 39200 25006 40000
rect 25318 39200 25374 40000
rect 25686 39200 25742 40000
rect 26054 39200 26110 40000
rect 26422 39200 26478 40000
rect 26790 39200 26846 40000
rect 27066 39200 27122 40000
rect 27434 39200 27490 40000
rect 27802 39200 27858 40000
rect 28170 39200 28226 40000
rect 28538 39200 28594 40000
rect 28814 39200 28870 40000
rect 29182 39200 29238 40000
rect 29550 39200 29606 40000
rect 29656 39222 29868 39250
rect 20088 37262 20116 39200
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 20088 35290 20116 37198
rect 20456 37126 20484 39200
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 20444 37120 20496 37126
rect 20444 37062 20496 37068
rect 20260 36780 20312 36786
rect 20260 36722 20312 36728
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20180 35494 20208 36110
rect 20168 35488 20220 35494
rect 20168 35430 20220 35436
rect 20076 35284 20128 35290
rect 20076 35226 20128 35232
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19352 34462 19472 34490
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18604 33516 18656 33522
rect 18604 33458 18656 33464
rect 18616 33114 18644 33458
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 18604 33108 18656 33114
rect 18604 33050 18656 33056
rect 19260 32910 19288 33254
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18524 31754 18552 31962
rect 18524 31726 18644 31754
rect 18328 30116 18380 30122
rect 18328 30058 18380 30064
rect 18340 28694 18368 30058
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 18432 28558 18460 29990
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 27470 18460 28358
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17972 22098 18000 23054
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17972 20058 18000 22034
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17972 18426 18000 19790
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18064 18290 18092 18634
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15502 18552 15846
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17788 13926 17908 13954
rect 17788 10266 17816 13926
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 12918 17908 13806
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17788 3602 17816 4014
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17328 800 17356 2382
rect 17696 2258 17724 2994
rect 17604 2230 17724 2258
rect 17604 800 17632 2230
rect 17880 800 17908 3334
rect 17972 3126 18000 14826
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18432 6934 18460 7482
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18524 5914 18552 13806
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18064 3058 18092 4422
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18156 2378 18184 3878
rect 18340 3058 18368 4966
rect 18524 3534 18552 5850
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18616 3194 18644 31726
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 18708 27606 18736 30194
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18800 16522 18828 30602
rect 18892 24206 18920 32710
rect 19260 30326 19288 32846
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19352 27130 19380 34462
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 19444 33454 19472 34342
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19444 32774 19472 33390
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 19536 32910 19564 33322
rect 19524 32904 19576 32910
rect 19524 32846 19576 32852
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19444 30326 19472 32710
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19444 30190 19472 30262
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19444 30054 19472 30126
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19996 26994 20024 34342
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19444 23526 19472 24074
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18892 16114 18920 18634
rect 19444 18630 19472 23462
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 20180 22094 20208 35430
rect 20272 34542 20300 36722
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20088 22066 20208 22094
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19514 20024 19858
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19812 18698 19840 19314
rect 19904 18970 19932 19382
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19996 18698 20024 19450
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5914 18736 6054
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 18156 800 18184 2314
rect 18432 800 18460 2314
rect 18708 800 18736 2790
rect 18800 2582 18828 8366
rect 19352 8362 19380 14554
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19812 12170 19840 12582
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19444 11830 19472 12106
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20088 11898 20116 22066
rect 20168 19236 20220 19242
rect 20168 19178 20220 19184
rect 20180 16114 20208 19178
rect 20272 19174 20300 34478
rect 20364 22778 20392 37062
rect 20824 36922 20852 39200
rect 21100 37262 21128 39200
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 21088 37256 21140 37262
rect 21088 37198 21140 37204
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20548 36378 20576 36722
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20444 36100 20496 36106
rect 20444 36042 20496 36048
rect 20456 34542 20484 36042
rect 20732 35494 20760 36110
rect 20916 35834 20944 37198
rect 21468 36922 21496 39200
rect 21456 36916 21508 36922
rect 21456 36858 21508 36864
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21008 36378 21036 36722
rect 21088 36712 21140 36718
rect 21088 36654 21140 36660
rect 21180 36712 21232 36718
rect 21180 36654 21232 36660
rect 20996 36372 21048 36378
rect 20996 36314 21048 36320
rect 20904 35828 20956 35834
rect 20904 35770 20956 35776
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20536 35216 20588 35222
rect 20536 35158 20588 35164
rect 20444 34536 20496 34542
rect 20444 34478 20496 34484
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20456 17338 20484 34478
rect 20548 33930 20576 35158
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20548 25430 20576 32846
rect 20536 25424 20588 25430
rect 20536 25366 20588 25372
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20180 15706 20208 16050
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19444 11354 19472 11766
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20180 8498 20208 8774
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20364 8430 20392 15438
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11762 20484 12038
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 6390 19380 7210
rect 20180 6730 20208 7278
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18892 1902 18920 5646
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18984 3534 19012 4966
rect 19062 4176 19118 4185
rect 19168 4146 19196 6190
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19352 4298 19380 4966
rect 19260 4270 19380 4298
rect 19062 4111 19118 4120
rect 19156 4140 19208 4146
rect 19076 4078 19104 4111
rect 19156 4082 19208 4088
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19260 3890 19288 4270
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19168 3862 19288 3890
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18880 1896 18932 1902
rect 18880 1838 18932 1844
rect 18984 800 19012 3062
rect 19168 2378 19196 3862
rect 19352 3738 19380 4082
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 19260 800 19288 3470
rect 19444 3058 19472 6598
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19812 4078 19840 4150
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19812 3738 19840 4014
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3194 20024 6666
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20088 4622 20116 5510
rect 20076 4616 20128 4622
rect 20180 4593 20208 6666
rect 20076 4558 20128 4564
rect 20166 4584 20222 4593
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19890 2544 19946 2553
rect 19444 1170 19472 2518
rect 19890 2479 19946 2488
rect 19904 2446 19932 2479
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 2088 20024 2994
rect 19812 2060 20024 2088
rect 19444 1142 19564 1170
rect 19536 800 19564 1142
rect 19812 800 19840 2060
rect 20088 800 20116 4558
rect 20166 4519 20222 4528
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 3126 20208 4422
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 20272 2446 20300 8298
rect 20548 7274 20576 17138
rect 20732 12442 20760 35430
rect 21100 34950 21128 36654
rect 21192 35086 21220 36654
rect 21836 36378 21864 39200
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 21824 36372 21876 36378
rect 21824 36314 21876 36320
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20916 24410 20944 24550
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20996 23588 21048 23594
rect 20996 23530 21048 23536
rect 21008 23050 21036 23530
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 21008 22710 21036 22986
rect 20996 22704 21048 22710
rect 20996 22646 21048 22652
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 21008 22030 21036 22374
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21008 19378 21036 21966
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21100 18426 21128 34886
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21192 22098 21220 23054
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 20810 14512 20866 14521
rect 20810 14447 20812 14456
rect 20864 14447 20866 14456
rect 20812 14418 20864 14424
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20640 8498 20668 8842
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20640 7750 20668 8434
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20364 3670 20392 4014
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 20456 3534 20484 4966
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4282 20576 4422
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20640 4010 20668 7686
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20456 3058 20484 3470
rect 20548 3194 20576 3878
rect 20732 3738 20760 8298
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6798 20852 7142
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 4622 20944 5510
rect 21008 4826 21036 11018
rect 21088 7268 21140 7274
rect 21088 7210 21140 7216
rect 21100 6798 21128 7210
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20364 800 20392 2790
rect 20640 800 20668 3470
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20732 2922 20760 3334
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20916 800 20944 4558
rect 21192 3534 21220 4966
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21192 800 21220 2790
rect 21284 2650 21312 33798
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 21468 25974 21496 31826
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21928 22094 21956 37266
rect 22204 37194 22232 39200
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 22008 36168 22060 36174
rect 22008 36110 22060 36116
rect 22020 35494 22048 36110
rect 22204 35834 22232 37130
rect 22572 36922 22600 39200
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22560 36780 22612 36786
rect 22560 36722 22612 36728
rect 22192 35828 22244 35834
rect 22192 35770 22244 35776
rect 22572 35766 22600 36722
rect 22836 36032 22888 36038
rect 22836 35974 22888 35980
rect 22560 35760 22612 35766
rect 22560 35702 22612 35708
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 21836 22066 21956 22094
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21560 9110 21588 17750
rect 21836 12374 21864 22066
rect 22020 15094 22048 35430
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22296 30190 22324 30534
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22296 29646 22324 29990
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22112 25498 22140 25842
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22204 22982 22232 25094
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22204 22574 22232 22918
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22388 17882 22416 18702
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22296 12986 22324 13126
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 22480 11830 22508 34886
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22664 26234 22692 31078
rect 22744 30660 22796 30666
rect 22744 30602 22796 30608
rect 22756 30394 22784 30602
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22848 26234 22876 35974
rect 22940 35834 22968 39200
rect 23216 36786 23244 39200
rect 23296 37120 23348 37126
rect 23296 37062 23348 37068
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23308 36530 23336 37062
rect 23584 36922 23612 39200
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23676 36802 23704 37810
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23584 36774 23704 36802
rect 23124 36502 23336 36530
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 22928 35828 22980 35834
rect 22928 35770 22980 35776
rect 23020 35692 23072 35698
rect 23020 35634 23072 35640
rect 23032 34950 23060 35634
rect 23020 34944 23072 34950
rect 23020 34886 23072 34892
rect 23124 32570 23152 36502
rect 23296 36100 23348 36106
rect 23296 36042 23348 36048
rect 23308 34610 23336 36042
rect 23296 34604 23348 34610
rect 23296 34546 23348 34552
rect 23112 32564 23164 32570
rect 23112 32506 23164 32512
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22940 29306 22968 30194
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 23400 26234 23428 36518
rect 23492 35834 23520 36722
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 22664 26206 22784 26234
rect 22848 26206 22968 26234
rect 22756 22710 22784 26206
rect 22836 25424 22888 25430
rect 22836 25366 22888 25372
rect 22848 25226 22876 25366
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22940 15162 22968 26206
rect 23308 26206 23428 26234
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23124 25294 23152 25638
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23308 20074 23336 26206
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23400 24206 23428 25230
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23400 22098 23428 24142
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23400 21554 23428 22034
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23308 20046 23428 20074
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23124 19378 23152 19790
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23124 18970 23152 19314
rect 23216 19242 23244 19654
rect 23204 19236 23256 19242
rect 23204 19178 23256 19184
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23216 18834 23244 19178
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23308 18766 23336 19926
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23400 17610 23428 20046
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 17678 23520 18566
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23388 17604 23440 17610
rect 23388 17546 23440 17552
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 13530 22600 14962
rect 22940 14482 22968 15098
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11082 22048 11698
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21468 4622 21496 4966
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21468 800 21496 4558
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 3534 21588 4422
rect 21652 4282 21680 5238
rect 22204 4622 22232 5510
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 22204 4146 22232 4558
rect 22296 4282 22324 5102
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21744 800 21772 4082
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22020 800 22048 3878
rect 22296 3602 22324 4218
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22112 2650 22140 2994
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22296 2514 22324 3538
rect 22388 3534 22416 4422
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 22480 2514 22508 4966
rect 22558 4040 22614 4049
rect 22558 3975 22614 3984
rect 22572 3670 22600 3975
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22664 3058 22692 4966
rect 22756 4690 22784 14350
rect 23584 8634 23612 36774
rect 23664 36644 23716 36650
rect 23664 36586 23716 36592
rect 23676 36310 23704 36586
rect 23952 36378 23980 39200
rect 24320 37262 24348 39200
rect 24308 37256 24360 37262
rect 24308 37198 24360 37204
rect 24124 37188 24176 37194
rect 24124 37130 24176 37136
rect 24136 36854 24164 37130
rect 24124 36848 24176 36854
rect 24124 36790 24176 36796
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 23664 36304 23716 36310
rect 23664 36246 23716 36252
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 13938 23704 35974
rect 24320 35834 24348 37198
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24308 35828 24360 35834
rect 24308 35770 24360 35776
rect 24032 34468 24084 34474
rect 24032 34410 24084 34416
rect 24044 33862 24072 34410
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23768 20058 23796 21490
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23768 19446 23796 19994
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 24216 18896 24268 18902
rect 24216 18838 24268 18844
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23768 14550 23796 14758
rect 23952 14618 23980 14758
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23676 13530 23704 13874
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23768 12646 23796 13330
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23768 12170 23796 12582
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23584 8362 23612 8570
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23952 7886 23980 8230
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23204 7812 23256 7818
rect 23204 7754 23256 7760
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22664 2774 22692 2994
rect 22572 2746 22692 2774
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22480 2394 22508 2450
rect 22296 2366 22508 2394
rect 22296 800 22324 2366
rect 22572 800 22600 2746
rect 22848 800 22876 3878
rect 22940 3126 22968 3946
rect 23032 3602 23060 4422
rect 23216 4146 23244 7754
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23400 3913 23428 5034
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23664 3936 23716 3942
rect 23386 3904 23442 3913
rect 23664 3878 23716 3884
rect 23386 3839 23442 3848
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 23032 1766 23060 3538
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 23020 1760 23072 1766
rect 23020 1702 23072 1708
rect 23124 800 23152 3062
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23400 800 23428 2994
rect 23676 800 23704 3878
rect 23768 3534 23796 4966
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23860 3126 23888 4422
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 24044 2774 24072 8910
rect 24136 3126 24164 13194
rect 24228 9654 24256 18838
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24412 14618 24440 14894
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24412 14006 24440 14554
rect 24400 14000 24452 14006
rect 24400 13942 24452 13948
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 23860 2746 24072 2774
rect 23860 2310 23888 2746
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23952 800 23980 2382
rect 24228 800 24256 3470
rect 24412 2446 24440 4966
rect 24504 3670 24532 14962
rect 24596 11694 24624 37062
rect 24688 36938 24716 39200
rect 24964 36938 24992 39200
rect 25332 37262 25360 39200
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25504 37256 25556 37262
rect 25504 37198 25556 37204
rect 24688 36922 24900 36938
rect 24964 36922 25084 36938
rect 24688 36916 24912 36922
rect 24688 36910 24860 36916
rect 24964 36916 25096 36922
rect 24964 36910 25044 36916
rect 24860 36858 24912 36864
rect 25044 36858 25096 36864
rect 24860 36712 24912 36718
rect 24688 36660 24860 36666
rect 24688 36654 24912 36660
rect 24688 36638 24900 36654
rect 24688 36582 24716 36638
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 25332 36378 25360 37198
rect 25412 36780 25464 36786
rect 25412 36722 25464 36728
rect 25320 36372 25372 36378
rect 25320 36314 25372 36320
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24872 35494 24900 36110
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24688 8838 24716 26862
rect 24872 14550 24900 35430
rect 24964 34542 24992 36042
rect 25424 35494 25452 36722
rect 25412 35488 25464 35494
rect 25412 35430 25464 35436
rect 24952 34536 25004 34542
rect 24952 34478 25004 34484
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25332 32230 25360 32370
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24872 8906 24900 9318
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24872 8634 24900 8842
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24872 8430 24900 8570
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24964 6866 24992 30262
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25240 29170 25268 29514
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25240 28082 25268 29106
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25332 26234 25360 32166
rect 25240 26206 25360 26234
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 22642 25176 24006
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25044 20324 25096 20330
rect 25044 20266 25096 20272
rect 25056 19922 25084 20266
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24596 3126 24624 5510
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24688 4282 24716 4422
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24688 3942 24716 4218
rect 24780 4146 24808 5714
rect 24872 5642 24900 6666
rect 25056 5914 25084 8978
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24872 3398 24900 5034
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 25056 4622 25084 4966
rect 25148 4826 25176 9522
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24492 2916 24544 2922
rect 24492 2858 24544 2864
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24504 800 24532 2858
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 24780 800 24808 2314
rect 25056 800 25084 4558
rect 25240 2417 25268 26206
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25332 13938 25360 14282
rect 25424 14006 25452 35430
rect 25516 35018 25544 37198
rect 25700 37126 25728 39200
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 25688 37120 25740 37126
rect 25688 37062 25740 37068
rect 25504 35012 25556 35018
rect 25504 34954 25556 34960
rect 25608 29714 25636 37062
rect 26068 36666 26096 39200
rect 26436 36786 26464 39200
rect 26700 37800 26752 37806
rect 26700 37742 26752 37748
rect 26608 37188 26660 37194
rect 26608 37130 26660 37136
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 26068 36650 26372 36666
rect 26068 36644 26384 36650
rect 26068 36638 26332 36644
rect 26332 36586 26384 36592
rect 26332 36372 26384 36378
rect 26332 36314 26384 36320
rect 26344 36038 26372 36314
rect 26436 36310 26464 36722
rect 26620 36378 26648 37130
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26424 36304 26476 36310
rect 26424 36246 26476 36252
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 26332 36032 26384 36038
rect 26332 35974 26384 35980
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 26240 35012 26292 35018
rect 26240 34954 26292 34960
rect 26252 34610 26280 34954
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 26344 32570 26372 35634
rect 26424 34944 26476 34950
rect 26424 34886 26476 34892
rect 26332 32564 26384 32570
rect 26332 32506 26384 32512
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 26252 31822 26280 32370
rect 26332 32224 26384 32230
rect 26332 32166 26384 32172
rect 26344 32026 26372 32166
rect 26332 32020 26384 32026
rect 26332 31962 26384 31968
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 26436 30546 26464 34886
rect 26528 32026 26556 36110
rect 26712 35894 26740 37742
rect 26804 37126 26832 39200
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 26792 37120 26844 37126
rect 26792 37062 26844 37068
rect 26884 36780 26936 36786
rect 26884 36722 26936 36728
rect 26712 35866 26832 35894
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26344 30518 26464 30546
rect 25596 29708 25648 29714
rect 25596 29650 25648 29656
rect 25780 28484 25832 28490
rect 25780 28426 25832 28432
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 25700 24410 25728 25162
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18698 25728 19110
rect 25596 18692 25648 18698
rect 25596 18634 25648 18640
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25504 16176 25556 16182
rect 25504 16118 25556 16124
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25332 3466 25360 3878
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25424 3058 25452 5850
rect 25516 3126 25544 16118
rect 25608 9042 25636 18634
rect 25792 12986 25820 28426
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 26160 27606 26188 28018
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26252 27470 26280 28018
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 26240 27056 26292 27062
rect 26240 26998 26292 27004
rect 26252 24342 26280 26998
rect 26240 24336 26292 24342
rect 26240 24278 26292 24284
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 26068 22778 26096 22986
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 25872 21412 25924 21418
rect 25872 21354 25924 21360
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25700 5710 25728 6394
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25884 4690 25912 21354
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 26068 18834 26096 19858
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26160 19242 26188 19450
rect 26148 19236 26200 19242
rect 26148 19178 26200 19184
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26056 18828 26108 18834
rect 26056 18770 26108 18776
rect 26252 18766 26280 19110
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26252 15434 26280 18566
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 26344 14006 26372 30518
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 26436 28082 26464 28358
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26436 26042 26464 28018
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 26436 25226 26464 25978
rect 26424 25220 26476 25226
rect 26424 25162 26476 25168
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26436 19122 26464 22374
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26516 19168 26568 19174
rect 26436 19116 26516 19122
rect 26436 19110 26568 19116
rect 26436 19094 26556 19110
rect 26436 18902 26464 19094
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 25596 4072 25648 4078
rect 25596 4014 25648 4020
rect 25608 3602 25636 4014
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25226 2408 25282 2417
rect 25226 2343 25282 2352
rect 25332 800 25360 2858
rect 25700 2854 25728 3878
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 25700 1442 25728 2790
rect 25608 1414 25728 1442
rect 25608 800 25636 1414
rect 25884 800 25912 3674
rect 25976 3058 26004 7686
rect 26160 7546 26188 9114
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26160 7410 26188 7482
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 26068 4010 26096 5306
rect 26252 4758 26280 7278
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 26056 4004 26108 4010
rect 26056 3946 26108 3952
rect 26528 3534 26556 5850
rect 26620 5370 26648 21082
rect 26804 11626 26832 35866
rect 26896 35578 26924 36722
rect 26988 35834 27016 37198
rect 27080 36922 27108 39200
rect 27068 36916 27120 36922
rect 27068 36858 27120 36864
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27264 36378 27292 36722
rect 27252 36372 27304 36378
rect 27252 36314 27304 36320
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 26976 35828 27028 35834
rect 26976 35770 27028 35776
rect 26896 35550 27016 35578
rect 26988 35494 27016 35550
rect 26976 35488 27028 35494
rect 26976 35430 27028 35436
rect 26988 30326 27016 35430
rect 27080 30938 27108 36110
rect 27448 35766 27476 39200
rect 27816 37126 27844 39200
rect 28078 37224 28134 37233
rect 28078 37159 28134 37168
rect 27804 37120 27856 37126
rect 27804 37062 27856 37068
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 27436 35760 27488 35766
rect 27436 35702 27488 35708
rect 27528 35692 27580 35698
rect 27528 35634 27580 35640
rect 27540 34746 27568 35634
rect 27528 34740 27580 34746
rect 27528 34682 27580 34688
rect 28000 34678 28028 36110
rect 27988 34672 28040 34678
rect 27988 34614 28040 34620
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 27540 33522 27568 34546
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27816 32910 27844 33390
rect 27896 33312 27948 33318
rect 27896 33254 27948 33260
rect 27804 32904 27856 32910
rect 27804 32846 27856 32852
rect 27804 32496 27856 32502
rect 27804 32438 27856 32444
rect 27528 31952 27580 31958
rect 27528 31894 27580 31900
rect 27540 31822 27568 31894
rect 27528 31816 27580 31822
rect 27528 31758 27580 31764
rect 27068 30932 27120 30938
rect 27068 30874 27120 30880
rect 27540 30802 27568 31758
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27160 30660 27212 30666
rect 27160 30602 27212 30608
rect 26976 30320 27028 30326
rect 26976 30262 27028 30268
rect 27172 28082 27200 30602
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 27080 27470 27108 27814
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27172 25974 27200 28018
rect 27448 27674 27476 28018
rect 27436 27668 27488 27674
rect 27436 27610 27488 27616
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27264 22574 27292 22918
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27264 19990 27292 22510
rect 27252 19984 27304 19990
rect 27252 19926 27304 19932
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26988 19514 27016 19654
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27264 19446 27292 19790
rect 27344 19780 27396 19786
rect 27344 19722 27396 19728
rect 27356 19446 27384 19722
rect 27252 19440 27304 19446
rect 27252 19382 27304 19388
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 26792 11620 26844 11626
rect 26792 11562 26844 11568
rect 26804 11354 26832 11562
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26896 8566 26924 11018
rect 27172 10062 27200 11494
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 26884 8560 26936 8566
rect 26884 8502 26936 8508
rect 26700 8492 26752 8498
rect 26700 8434 26752 8440
rect 26712 5914 26740 8434
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26804 7002 26832 7210
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 26160 800 26188 3334
rect 26620 2774 26648 4966
rect 26700 4616 26752 4622
rect 26700 4558 26752 4564
rect 26712 4010 26740 4558
rect 26700 4004 26752 4010
rect 26700 3946 26752 3952
rect 26804 3534 26832 5510
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 26896 4690 26924 5238
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 26988 3942 27016 8842
rect 27264 7562 27292 15846
rect 27356 15638 27384 19382
rect 27344 15632 27396 15638
rect 27344 15574 27396 15580
rect 27816 11286 27844 32438
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 27816 10810 27844 11222
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27436 8832 27488 8838
rect 27436 8774 27488 8780
rect 27172 7534 27292 7562
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26620 2746 26740 2774
rect 26712 2446 26740 2746
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 26436 800 26464 2314
rect 26712 800 26740 2382
rect 26896 800 26924 3334
rect 27172 2553 27200 7534
rect 27252 6180 27304 6186
rect 27252 6122 27304 6128
rect 27264 2582 27292 6122
rect 27448 5302 27476 8774
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27632 6390 27660 6734
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27436 5296 27488 5302
rect 27436 5238 27488 5244
rect 27448 4826 27476 5238
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 27344 4548 27396 4554
rect 27344 4490 27396 4496
rect 27252 2576 27304 2582
rect 27158 2544 27214 2553
rect 27252 2518 27304 2524
rect 27158 2479 27214 2488
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27172 800 27200 2382
rect 27356 2378 27384 4490
rect 27540 4146 27568 4966
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27540 3738 27568 4082
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27816 3534 27844 7142
rect 27908 5409 27936 33254
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 28000 12102 28028 21422
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 28000 11218 28028 11766
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27988 9512 28040 9518
rect 27988 9454 28040 9460
rect 27894 5400 27950 5409
rect 27894 5335 27950 5344
rect 28000 5114 28028 9454
rect 27908 5086 28028 5114
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27344 2372 27396 2378
rect 27344 2314 27396 2320
rect 27448 800 27476 3062
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 27540 1970 27568 2858
rect 27528 1964 27580 1970
rect 27528 1906 27580 1912
rect 27724 800 27752 3334
rect 27908 2922 27936 5086
rect 27988 5024 28040 5030
rect 27988 4966 28040 4972
rect 28000 3126 28028 4966
rect 28092 4078 28120 37159
rect 28184 36922 28212 39200
rect 28552 37262 28580 39200
rect 28828 37618 28856 39200
rect 28828 37590 28948 37618
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28816 37256 28868 37262
rect 28816 37198 28868 37204
rect 28448 37188 28500 37194
rect 28448 37130 28500 37136
rect 28172 36916 28224 36922
rect 28172 36858 28224 36864
rect 28460 36242 28488 37130
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28644 36378 28672 36722
rect 28632 36372 28684 36378
rect 28632 36314 28684 36320
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 28736 35894 28764 37062
rect 28828 36378 28856 37198
rect 28816 36372 28868 36378
rect 28816 36314 28868 36320
rect 28816 36168 28868 36174
rect 28816 36110 28868 36116
rect 28644 35866 28764 35894
rect 28172 35488 28224 35494
rect 28172 35430 28224 35436
rect 28184 35222 28212 35430
rect 28172 35216 28224 35222
rect 28172 35158 28224 35164
rect 28448 35080 28500 35086
rect 28448 35022 28500 35028
rect 28460 33046 28488 35022
rect 28448 33040 28500 33046
rect 28448 32982 28500 32988
rect 28460 31822 28488 32982
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28172 25152 28224 25158
rect 28172 25094 28224 25100
rect 28184 24614 28212 25094
rect 28172 24608 28224 24614
rect 28172 24550 28224 24556
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 20534 28304 23054
rect 28264 20528 28316 20534
rect 28264 20470 28316 20476
rect 28276 19310 28304 20470
rect 28264 19304 28316 19310
rect 28264 19246 28316 19252
rect 28276 17542 28304 19246
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 28276 15706 28304 17478
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28356 12096 28408 12102
rect 28356 12038 28408 12044
rect 28368 11626 28396 12038
rect 28356 11620 28408 11626
rect 28356 11562 28408 11568
rect 28540 11552 28592 11558
rect 28540 11494 28592 11500
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28460 9654 28488 11154
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 28552 9586 28580 11494
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28172 6656 28224 6662
rect 28172 6598 28224 6604
rect 28184 4146 28212 6598
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 28172 4004 28224 4010
rect 28172 3946 28224 3952
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 27896 2916 27948 2922
rect 27896 2858 27948 2864
rect 28092 2774 28120 2994
rect 28000 2746 28120 2774
rect 28000 800 28028 2746
rect 28184 2394 28212 3946
rect 28276 2446 28304 4422
rect 28368 4010 28396 7686
rect 28644 7546 28672 35866
rect 28828 35290 28856 36110
rect 28920 35834 28948 37590
rect 29092 37460 29144 37466
rect 29092 37402 29144 37408
rect 29104 35894 29132 37402
rect 29196 36922 29224 39200
rect 29564 39114 29592 39200
rect 29656 39114 29684 39222
rect 29564 39086 29684 39114
rect 29552 37256 29604 37262
rect 29552 37198 29604 37204
rect 29184 36916 29236 36922
rect 29184 36858 29236 36864
rect 29276 36780 29328 36786
rect 29276 36722 29328 36728
rect 29288 36310 29316 36722
rect 29276 36304 29328 36310
rect 29276 36246 29328 36252
rect 29368 36304 29420 36310
rect 29368 36246 29420 36252
rect 29380 36145 29408 36246
rect 29366 36136 29422 36145
rect 29366 36071 29422 36080
rect 29104 35866 29316 35894
rect 28908 35828 28960 35834
rect 28908 35770 28960 35776
rect 28816 35284 28868 35290
rect 28816 35226 28868 35232
rect 28908 35216 28960 35222
rect 28908 35158 28960 35164
rect 28724 34060 28776 34066
rect 28724 34002 28776 34008
rect 28736 8786 28764 34002
rect 28920 26234 28948 35158
rect 29000 34944 29052 34950
rect 29000 34886 29052 34892
rect 29012 28626 29040 34886
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 29196 32026 29224 33458
rect 29184 32020 29236 32026
rect 29184 31962 29236 31968
rect 29000 28620 29052 28626
rect 29000 28562 29052 28568
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 28828 26206 28948 26234
rect 28828 8922 28856 26206
rect 29012 25226 29040 28426
rect 29000 25220 29052 25226
rect 29000 25162 29052 25168
rect 29012 20534 29040 25162
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29012 15162 29040 16050
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 29196 15094 29224 15506
rect 29184 15088 29236 15094
rect 29184 15030 29236 15036
rect 28908 12844 28960 12850
rect 28908 12786 28960 12792
rect 28920 11898 28948 12786
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 28828 8894 28948 8922
rect 28736 8758 28856 8786
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28828 5030 28856 8758
rect 28920 5250 28948 8894
rect 29000 7812 29052 7818
rect 29000 7754 29052 7760
rect 29012 7274 29040 7754
rect 29000 7268 29052 7274
rect 29000 7210 29052 7216
rect 29288 5370 29316 35866
rect 29564 35562 29592 37198
rect 29840 37126 29868 39222
rect 29918 39200 29974 40000
rect 30286 39200 30342 40000
rect 30562 39200 30618 40000
rect 30930 39200 30986 40000
rect 31298 39200 31354 40000
rect 31666 39200 31722 40000
rect 32034 39200 32090 40000
rect 32402 39200 32458 40000
rect 32678 39200 32734 40000
rect 33046 39200 33102 40000
rect 33414 39200 33470 40000
rect 33782 39200 33838 40000
rect 34150 39200 34206 40000
rect 34426 39200 34482 40000
rect 34794 39200 34850 40000
rect 35162 39200 35218 40000
rect 35530 39200 35586 40000
rect 35898 39200 35954 40000
rect 36266 39200 36322 40000
rect 36542 39200 36598 40000
rect 36910 39200 36966 40000
rect 37016 39222 37228 39250
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29748 35834 29776 37062
rect 29932 36922 29960 39200
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29552 35556 29604 35562
rect 29552 35498 29604 35504
rect 29460 35488 29512 35494
rect 29460 35430 29512 35436
rect 29472 35154 29500 35430
rect 29460 35148 29512 35154
rect 29460 35090 29512 35096
rect 30024 33658 30052 36722
rect 30194 36272 30250 36281
rect 30194 36207 30250 36216
rect 30208 36174 30236 36207
rect 30196 36168 30248 36174
rect 30196 36110 30248 36116
rect 30300 35834 30328 39200
rect 30576 37262 30604 39200
rect 30656 37324 30708 37330
rect 30656 37266 30708 37272
rect 30564 37256 30616 37262
rect 30564 37198 30616 37204
rect 30472 36100 30524 36106
rect 30472 36042 30524 36048
rect 30288 35828 30340 35834
rect 30288 35770 30340 35776
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 30012 33652 30064 33658
rect 30012 33594 30064 33600
rect 30104 32020 30156 32026
rect 30104 31962 30156 31968
rect 29920 24132 29972 24138
rect 29920 24074 29972 24080
rect 29932 23526 29960 24074
rect 29920 23520 29972 23526
rect 29920 23462 29972 23468
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29460 14884 29512 14890
rect 29460 14826 29512 14832
rect 29472 14618 29500 14826
rect 29460 14612 29512 14618
rect 29460 14554 29512 14560
rect 29564 12434 29592 21830
rect 29472 12406 29592 12434
rect 29368 7336 29420 7342
rect 29368 7278 29420 7284
rect 29276 5364 29328 5370
rect 29276 5306 29328 5312
rect 28920 5222 29040 5250
rect 29288 5234 29316 5306
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28356 4004 28408 4010
rect 28356 3946 28408 3952
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 28356 3460 28408 3466
rect 28356 3402 28408 3408
rect 28368 3126 28396 3402
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 28356 3120 28408 3126
rect 28356 3062 28408 3068
rect 28092 2378 28212 2394
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28080 2372 28212 2378
rect 28132 2366 28212 2372
rect 28080 2314 28132 2320
rect 28172 2304 28224 2310
rect 28460 2258 28488 3334
rect 28172 2246 28224 2252
rect 28184 1902 28212 2246
rect 28276 2230 28488 2258
rect 28172 1896 28224 1902
rect 28172 1838 28224 1844
rect 28276 800 28304 2230
rect 28552 800 28580 3878
rect 28644 3534 28672 4558
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 28736 3058 28764 4966
rect 29012 4282 29040 5222
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29276 4480 29328 4486
rect 29276 4422 29328 4428
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 28828 3670 28856 4082
rect 29288 4078 29316 4422
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 29184 4004 29236 4010
rect 29184 3946 29236 3952
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 28816 3664 28868 3670
rect 28816 3606 28868 3612
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28828 800 28856 3062
rect 29012 2446 29040 3878
rect 29196 3670 29224 3946
rect 29184 3664 29236 3670
rect 29184 3606 29236 3612
rect 29288 3466 29316 4014
rect 29276 3460 29328 3466
rect 29276 3402 29328 3408
rect 29380 3058 29408 7278
rect 29472 3534 29500 12406
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29552 4004 29604 4010
rect 29552 3946 29604 3952
rect 29564 3738 29592 3946
rect 29552 3732 29604 3738
rect 29552 3674 29604 3680
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 29104 800 29132 2382
rect 29564 2088 29592 3538
rect 29656 2514 29684 6054
rect 29840 5914 29868 6190
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 29736 5568 29788 5574
rect 29736 5510 29788 5516
rect 29748 3126 29776 5510
rect 29828 3936 29880 3942
rect 29828 3878 29880 3884
rect 29840 3602 29868 3878
rect 29828 3596 29880 3602
rect 29828 3538 29880 3544
rect 29736 3120 29788 3126
rect 29736 3062 29788 3068
rect 29932 2514 29960 23462
rect 30116 8090 30144 31962
rect 30288 30116 30340 30122
rect 30288 30058 30340 30064
rect 30300 29170 30328 30058
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30300 27946 30328 29106
rect 30288 27940 30340 27946
rect 30288 27882 30340 27888
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30208 19514 30236 19858
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 30392 16250 30420 34886
rect 30484 21894 30512 36042
rect 30576 35766 30604 37198
rect 30564 35760 30616 35766
rect 30564 35702 30616 35708
rect 30564 35080 30616 35086
rect 30564 35022 30616 35028
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30576 16250 30604 35022
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30576 15162 30604 16050
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30104 8084 30156 8090
rect 30104 8026 30156 8032
rect 30012 7812 30064 7818
rect 30012 7754 30064 7760
rect 30024 6866 30052 7754
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 30012 6656 30064 6662
rect 30012 6598 30064 6604
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30024 3602 30052 6598
rect 30104 6180 30156 6186
rect 30104 6122 30156 6128
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 29644 2508 29696 2514
rect 29644 2450 29696 2456
rect 29920 2508 29972 2514
rect 29920 2450 29972 2456
rect 29380 2060 29592 2088
rect 29380 800 29408 2060
rect 29656 800 29684 2450
rect 30024 2394 30052 3538
rect 30116 2446 30144 6122
rect 30472 6112 30524 6118
rect 30472 6054 30524 6060
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30392 4570 30420 5102
rect 30208 4542 30420 4570
rect 30208 3670 30236 4542
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30300 3913 30328 4082
rect 30286 3904 30342 3913
rect 30286 3839 30342 3848
rect 30196 3664 30248 3670
rect 30196 3606 30248 3612
rect 30392 2774 30420 4422
rect 30484 3058 30512 6054
rect 30576 4554 30604 6598
rect 30668 5914 30696 37266
rect 30944 36922 30972 39200
rect 31208 37256 31260 37262
rect 31208 37198 31260 37204
rect 31220 37126 31248 37198
rect 31208 37120 31260 37126
rect 31208 37062 31260 37068
rect 30932 36916 30984 36922
rect 30932 36858 30984 36864
rect 31116 36848 31168 36854
rect 31116 36790 31168 36796
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 30932 36100 30984 36106
rect 30932 36042 30984 36048
rect 30748 30048 30800 30054
rect 30748 29990 30800 29996
rect 30760 25974 30788 29990
rect 30840 28484 30892 28490
rect 30840 28426 30892 28432
rect 30852 28218 30880 28426
rect 30840 28212 30892 28218
rect 30840 28154 30892 28160
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30852 27334 30880 27406
rect 30840 27328 30892 27334
rect 30840 27270 30892 27276
rect 30852 26586 30880 27270
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 30852 26042 30880 26522
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 30748 25968 30800 25974
rect 30748 25910 30800 25916
rect 30944 25498 30972 36042
rect 31036 34950 31064 36722
rect 31128 36242 31156 36790
rect 31116 36236 31168 36242
rect 31116 36178 31168 36184
rect 31220 35834 31248 37062
rect 31312 36378 31340 39200
rect 31484 37732 31536 37738
rect 31484 37674 31536 37680
rect 31300 36372 31352 36378
rect 31300 36314 31352 36320
rect 31208 35828 31260 35834
rect 31208 35770 31260 35776
rect 31300 35692 31352 35698
rect 31300 35634 31352 35640
rect 31024 34944 31076 34950
rect 31024 34886 31076 34892
rect 31312 34202 31340 35634
rect 31300 34196 31352 34202
rect 31300 34138 31352 34144
rect 31496 34134 31524 37674
rect 31576 37664 31628 37670
rect 31576 37606 31628 37612
rect 31484 34128 31536 34134
rect 31484 34070 31536 34076
rect 31484 33992 31536 33998
rect 31484 33934 31536 33940
rect 31496 32570 31524 33934
rect 31484 32564 31536 32570
rect 31484 32506 31536 32512
rect 31392 29572 31444 29578
rect 31392 29514 31444 29520
rect 31404 29034 31432 29514
rect 31392 29028 31444 29034
rect 31392 28970 31444 28976
rect 31404 28150 31432 28970
rect 31392 28144 31444 28150
rect 31392 28086 31444 28092
rect 31404 27402 31432 28086
rect 31392 27396 31444 27402
rect 31392 27338 31444 27344
rect 30932 25492 30984 25498
rect 30932 25434 30984 25440
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30668 5710 30696 5850
rect 30656 5704 30708 5710
rect 30656 5646 30708 5652
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30564 4548 30616 4554
rect 30564 4490 30616 4496
rect 30564 4140 30616 4146
rect 30668 4128 30696 5510
rect 30760 4146 30788 9862
rect 30616 4100 30696 4128
rect 30748 4140 30800 4146
rect 30564 4082 30616 4088
rect 30748 4082 30800 4088
rect 30576 3398 30604 4082
rect 30564 3392 30616 3398
rect 30564 3334 30616 3340
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30208 2746 30420 2774
rect 29932 2366 30052 2394
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 29932 800 29960 2366
rect 30208 800 30236 2746
rect 30484 800 30512 2994
rect 30760 800 30788 3334
rect 30852 3058 30880 24074
rect 31024 21616 31076 21622
rect 31024 21558 31076 21564
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30944 19378 30972 19654
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 31036 12442 31064 21558
rect 31024 12436 31076 12442
rect 31024 12378 31076 12384
rect 31116 12164 31168 12170
rect 31116 12106 31168 12112
rect 31128 11898 31156 12106
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31208 11620 31260 11626
rect 31208 11562 31260 11568
rect 31024 9444 31076 9450
rect 31024 9386 31076 9392
rect 30932 6112 30984 6118
rect 30932 6054 30984 6060
rect 30944 5574 30972 6054
rect 30932 5568 30984 5574
rect 30932 5510 30984 5516
rect 30932 5364 30984 5370
rect 30932 5306 30984 5312
rect 30944 3534 30972 5306
rect 31036 4622 31064 9386
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 31128 4706 31156 5510
rect 31220 4826 31248 11562
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 31128 4678 31248 4706
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 31128 4214 31156 4558
rect 31116 4208 31168 4214
rect 31116 4150 31168 4156
rect 31220 3584 31248 4678
rect 31312 3738 31340 25094
rect 31404 24206 31432 25298
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31404 23798 31432 24142
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 31404 23186 31432 23734
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31404 22166 31432 23122
rect 31392 22160 31444 22166
rect 31392 22102 31444 22108
rect 31392 16584 31444 16590
rect 31392 16526 31444 16532
rect 31404 15706 31432 16526
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31496 14006 31524 15302
rect 31484 14000 31536 14006
rect 31484 13942 31536 13948
rect 31588 6866 31616 37606
rect 31680 37244 31708 39200
rect 31760 37256 31812 37262
rect 31680 37216 31760 37244
rect 31760 37198 31812 37204
rect 32048 36922 32076 39200
rect 32036 36916 32088 36922
rect 32036 36858 32088 36864
rect 31944 36780 31996 36786
rect 31944 36722 31996 36728
rect 31668 36168 31720 36174
rect 31668 36110 31720 36116
rect 31680 35086 31708 36110
rect 31668 35080 31720 35086
rect 31668 35022 31720 35028
rect 31956 34950 31984 36722
rect 32416 35562 32444 39200
rect 32496 37324 32548 37330
rect 32496 37266 32548 37272
rect 32404 35556 32456 35562
rect 32404 35498 32456 35504
rect 31944 34944 31996 34950
rect 31944 34886 31996 34892
rect 31668 34128 31720 34134
rect 31668 34070 31720 34076
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 31392 6112 31444 6118
rect 31392 6054 31444 6060
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31220 3556 31340 3584
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 31036 800 31064 3334
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 2038 31156 2246
rect 31116 2032 31168 2038
rect 31116 1974 31168 1980
rect 31312 800 31340 3556
rect 31404 3466 31432 6054
rect 31680 5914 31708 34070
rect 31760 28076 31812 28082
rect 31760 28018 31812 28024
rect 31772 27538 31800 28018
rect 31760 27532 31812 27538
rect 31760 27474 31812 27480
rect 31852 23724 31904 23730
rect 31852 23666 31904 23672
rect 31864 23526 31892 23666
rect 31852 23520 31904 23526
rect 31852 23462 31904 23468
rect 31864 16574 31892 23462
rect 31956 16658 31984 34886
rect 32404 30320 32456 30326
rect 32404 30262 32456 30268
rect 32220 30252 32272 30258
rect 32220 30194 32272 30200
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 32140 29714 32168 30126
rect 32128 29708 32180 29714
rect 32128 29650 32180 29656
rect 32232 29646 32260 30194
rect 32312 29776 32364 29782
rect 32312 29718 32364 29724
rect 32220 29640 32272 29646
rect 32220 29582 32272 29588
rect 32220 21684 32272 21690
rect 32220 21626 32272 21632
rect 32128 17264 32180 17270
rect 32128 17206 32180 17212
rect 31944 16652 31996 16658
rect 31944 16594 31996 16600
rect 31772 16546 31892 16574
rect 31668 5908 31720 5914
rect 31668 5850 31720 5856
rect 31484 5296 31536 5302
rect 31484 5238 31536 5244
rect 31496 4486 31524 5238
rect 31680 5234 31708 5850
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 31576 4548 31628 4554
rect 31576 4490 31628 4496
rect 31484 4480 31536 4486
rect 31484 4422 31536 4428
rect 31392 3460 31444 3466
rect 31392 3402 31444 3408
rect 31588 800 31616 4490
rect 31772 3618 31800 16546
rect 32036 11552 32088 11558
rect 32036 11494 32088 11500
rect 31944 9376 31996 9382
rect 31944 9318 31996 9324
rect 31852 5568 31904 5574
rect 31852 5510 31904 5516
rect 31864 5234 31892 5510
rect 31956 5250 31984 9318
rect 32048 5370 32076 11494
rect 32140 8566 32168 17206
rect 32128 8560 32180 8566
rect 32128 8502 32180 8508
rect 32128 8424 32180 8430
rect 32128 8366 32180 8372
rect 32140 7818 32168 8366
rect 32232 7954 32260 21626
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 32140 6866 32168 7754
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 32036 5364 32088 5370
rect 32036 5306 32088 5312
rect 31852 5228 31904 5234
rect 31956 5222 32168 5250
rect 31852 5170 31904 5176
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31726 3590 31800 3618
rect 31726 3346 31754 3590
rect 31726 3318 31800 3346
rect 31772 2514 31800 3318
rect 31760 2508 31812 2514
rect 31760 2450 31812 2456
rect 31864 800 31892 3878
rect 31956 3602 31984 4966
rect 32140 4146 32168 5222
rect 32232 4706 32260 6598
rect 32324 4826 32352 29718
rect 32416 29646 32444 30262
rect 32404 29640 32456 29646
rect 32404 29582 32456 29588
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32416 27470 32444 27814
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32508 26234 32536 37266
rect 32692 37244 32720 39200
rect 32772 37256 32824 37262
rect 32692 37216 32772 37244
rect 32772 37198 32824 37204
rect 33060 36938 33088 39200
rect 33060 36922 33180 36938
rect 33060 36916 33192 36922
rect 33060 36910 33140 36916
rect 33140 36858 33192 36864
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 33152 35894 33180 36722
rect 33232 36100 33284 36106
rect 33232 36042 33284 36048
rect 33060 35866 33180 35894
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 32968 34950 32996 35634
rect 32956 34944 33008 34950
rect 32956 34886 33008 34892
rect 32864 34536 32916 34542
rect 32864 34478 32916 34484
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32784 32366 32812 32846
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 32876 32026 32904 34478
rect 32864 32020 32916 32026
rect 32864 31962 32916 31968
rect 32864 30864 32916 30870
rect 32864 30806 32916 30812
rect 32588 30660 32640 30666
rect 32588 30602 32640 30608
rect 32600 30394 32628 30602
rect 32588 30388 32640 30394
rect 32588 30330 32640 30336
rect 32876 29850 32904 30806
rect 32968 30326 32996 34886
rect 33060 34542 33088 35866
rect 33140 35012 33192 35018
rect 33140 34954 33192 34960
rect 33048 34536 33100 34542
rect 33048 34478 33100 34484
rect 33152 34202 33180 34954
rect 33140 34196 33192 34202
rect 33140 34138 33192 34144
rect 33048 31340 33100 31346
rect 33048 31282 33100 31288
rect 33060 30938 33088 31282
rect 33048 30932 33100 30938
rect 33048 30874 33100 30880
rect 32956 30320 33008 30326
rect 32956 30262 33008 30268
rect 32864 29844 32916 29850
rect 32864 29786 32916 29792
rect 32588 29640 32640 29646
rect 32588 29582 32640 29588
rect 32600 28082 32628 29582
rect 32588 28076 32640 28082
rect 32588 28018 32640 28024
rect 32600 27334 32628 28018
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32600 27130 32628 27270
rect 32588 27124 32640 27130
rect 32588 27066 32640 27072
rect 32508 26206 32628 26234
rect 32600 15706 32628 26206
rect 33244 22778 33272 36042
rect 33428 35834 33456 39200
rect 33796 37262 33824 39200
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 33416 35828 33468 35834
rect 33416 35770 33468 35776
rect 33520 35290 33548 37198
rect 34164 36922 34192 39200
rect 34336 37188 34388 37194
rect 34336 37130 34388 37136
rect 34152 36916 34204 36922
rect 34152 36858 34204 36864
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 33968 36100 34020 36106
rect 33968 36042 34020 36048
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 33876 35692 33928 35698
rect 33876 35634 33928 35640
rect 33508 35284 33560 35290
rect 33508 35226 33560 35232
rect 33600 34944 33652 34950
rect 33600 34886 33652 34892
rect 33508 33992 33560 33998
rect 33508 33934 33560 33940
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 33324 30320 33376 30326
rect 33324 30262 33376 30268
rect 33232 22772 33284 22778
rect 33232 22714 33284 22720
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 32968 22438 32996 22578
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32404 12776 32456 12782
rect 32404 12718 32456 12724
rect 32416 11830 32444 12718
rect 32404 11824 32456 11830
rect 32404 11766 32456 11772
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32416 5370 32444 7822
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32404 5364 32456 5370
rect 32404 5306 32456 5312
rect 32312 4820 32364 4826
rect 32312 4762 32364 4768
rect 32232 4678 32352 4706
rect 32220 4208 32272 4214
rect 32220 4150 32272 4156
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32232 4010 32260 4150
rect 32324 4146 32352 4678
rect 32404 4276 32456 4282
rect 32404 4218 32456 4224
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32416 4010 32444 4218
rect 32220 4004 32272 4010
rect 32220 3946 32272 3952
rect 32404 4004 32456 4010
rect 32404 3946 32456 3952
rect 32220 3732 32272 3738
rect 32220 3674 32272 3680
rect 31944 3596 31996 3602
rect 31944 3538 31996 3544
rect 32232 2446 32260 3674
rect 32600 3058 32628 6598
rect 32692 5914 32720 8434
rect 32864 6112 32916 6118
rect 32864 6054 32916 6060
rect 32680 5908 32732 5914
rect 32680 5850 32732 5856
rect 32772 5296 32824 5302
rect 32772 5238 32824 5244
rect 32784 4214 32812 5238
rect 32876 5234 32904 6054
rect 32864 5228 32916 5234
rect 32864 5170 32916 5176
rect 32772 4208 32824 4214
rect 32772 4150 32824 4156
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 32220 2440 32272 2446
rect 32140 2400 32220 2428
rect 32140 800 32168 2400
rect 32220 2382 32272 2388
rect 32416 800 32444 2994
rect 32692 800 32720 3334
rect 32876 2774 32904 5170
rect 32968 3058 32996 22374
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33244 19514 33272 19790
rect 33232 19508 33284 19514
rect 33232 19450 33284 19456
rect 33244 19378 33272 19450
rect 33232 19372 33284 19378
rect 33232 19314 33284 19320
rect 33048 9716 33100 9722
rect 33048 9658 33100 9664
rect 33060 8974 33088 9658
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 33336 8566 33364 30262
rect 33428 30258 33456 31078
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 33520 26234 33548 33934
rect 33428 26206 33548 26234
rect 33324 8560 33376 8566
rect 33324 8502 33376 8508
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 33046 3496 33102 3505
rect 33046 3431 33048 3440
rect 33100 3431 33102 3440
rect 33048 3402 33100 3408
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 32876 2746 32996 2774
rect 32968 800 32996 2746
rect 33244 800 33272 5510
rect 33336 2990 33364 6598
rect 33428 4826 33456 26206
rect 33612 11286 33640 34886
rect 33704 34542 33732 35634
rect 33692 34536 33744 34542
rect 33692 34478 33744 34484
rect 33704 17202 33732 34478
rect 33888 33862 33916 35634
rect 33876 33856 33928 33862
rect 33876 33798 33928 33804
rect 33888 29782 33916 33798
rect 33876 29776 33928 29782
rect 33876 29718 33928 29724
rect 33784 24132 33836 24138
rect 33784 24074 33836 24080
rect 33796 23118 33824 24074
rect 33980 23526 34008 36042
rect 34256 34950 34284 36722
rect 34244 34944 34296 34950
rect 34244 34886 34296 34892
rect 34348 26234 34376 37130
rect 34440 36378 34468 39200
rect 34808 37210 34836 39200
rect 35176 37754 35204 39200
rect 35176 37726 35388 37754
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34808 37182 34928 37210
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 34520 36780 34572 36786
rect 34520 36722 34572 36728
rect 34428 36372 34480 36378
rect 34428 36314 34480 36320
rect 34532 35222 34560 36722
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 34520 35216 34572 35222
rect 34520 35158 34572 35164
rect 34428 34536 34480 34542
rect 34428 34478 34480 34484
rect 34256 26206 34376 26234
rect 33968 23520 34020 23526
rect 33968 23462 34020 23468
rect 33784 23112 33836 23118
rect 33784 23054 33836 23060
rect 33796 22574 33824 23054
rect 33784 22568 33836 22574
rect 33784 22510 33836 22516
rect 33692 17196 33744 17202
rect 33692 17138 33744 17144
rect 33796 12782 33824 22510
rect 34256 17270 34284 26206
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 34348 19514 34376 19654
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 34244 17264 34296 17270
rect 34244 17206 34296 17212
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34164 16250 34192 17070
rect 34152 16244 34204 16250
rect 34152 16186 34204 16192
rect 33784 12776 33836 12782
rect 33784 12718 33836 12724
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33600 11280 33652 11286
rect 33600 11222 33652 11228
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33508 6112 33560 6118
rect 33508 6054 33560 6060
rect 33520 5216 33548 6054
rect 33612 5370 33640 8434
rect 33784 6996 33836 7002
rect 33784 6938 33836 6944
rect 33796 5914 33824 6938
rect 33784 5908 33836 5914
rect 33704 5868 33784 5896
rect 33600 5364 33652 5370
rect 33600 5306 33652 5312
rect 33520 5188 33640 5216
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 33520 4826 33548 5034
rect 33416 4820 33468 4826
rect 33416 4762 33468 4768
rect 33508 4820 33560 4826
rect 33508 4762 33560 4768
rect 33324 2984 33376 2990
rect 33324 2926 33376 2932
rect 33612 2922 33640 5188
rect 33704 4622 33732 5868
rect 33784 5850 33836 5856
rect 33784 5092 33836 5098
rect 33784 5034 33836 5040
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33796 4486 33824 5034
rect 33784 4480 33836 4486
rect 33784 4422 33836 4428
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33796 3058 33824 3878
rect 33888 3534 33916 12582
rect 34336 7200 34388 7206
rect 34336 7142 34388 7148
rect 33968 6656 34020 6662
rect 33968 6598 34020 6604
rect 33980 5234 34008 6598
rect 34060 6112 34112 6118
rect 34060 6054 34112 6060
rect 34072 5710 34100 6054
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 33968 5228 34020 5234
rect 33968 5170 34020 5176
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 33600 2916 33652 2922
rect 33600 2858 33652 2864
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33520 800 33548 2790
rect 33612 2774 33640 2858
rect 33980 2774 34008 5170
rect 33612 2746 33732 2774
rect 33704 2446 33732 2746
rect 33796 2746 34008 2774
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33796 800 33824 2746
rect 33968 2304 34020 2310
rect 33968 2246 34020 2252
rect 33980 1834 34008 2246
rect 33968 1828 34020 1834
rect 33968 1770 34020 1776
rect 34072 800 34100 5646
rect 34152 4480 34204 4486
rect 34152 4422 34204 4428
rect 34164 4146 34192 4422
rect 34152 4140 34204 4146
rect 34152 4082 34204 4088
rect 34348 4010 34376 7142
rect 34440 5370 34468 34478
rect 34716 33998 34744 36110
rect 34704 33992 34756 33998
rect 34704 33934 34756 33940
rect 34808 26234 34836 37062
rect 34900 36854 34928 37182
rect 35360 36922 35388 37726
rect 35544 37618 35572 39200
rect 35806 39128 35862 39137
rect 35806 39063 35862 39072
rect 35544 37590 35664 37618
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 35348 36916 35400 36922
rect 35348 36858 35400 36864
rect 34888 36848 34940 36854
rect 34888 36790 34940 36796
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35452 36378 35480 37198
rect 35532 37120 35584 37126
rect 35532 37062 35584 37068
rect 35440 36372 35492 36378
rect 35440 36314 35492 36320
rect 35348 35692 35400 35698
rect 35348 35634 35400 35640
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35360 33318 35388 35634
rect 35348 33312 35400 33318
rect 35348 33254 35400 33260
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35348 32428 35400 32434
rect 35348 32370 35400 32376
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35360 31482 35388 32370
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35440 27396 35492 27402
rect 35440 27338 35492 27344
rect 35452 26994 35480 27338
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34624 26206 34836 26234
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 9178 34560 23462
rect 34624 17882 34652 26206
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35544 21146 35572 37062
rect 35636 35834 35664 37590
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35728 36854 35756 37198
rect 35716 36848 35768 36854
rect 35716 36790 35768 36796
rect 35714 35864 35770 35873
rect 35624 35828 35676 35834
rect 35714 35799 35770 35808
rect 35624 35770 35676 35776
rect 35624 35692 35676 35698
rect 35624 35634 35676 35640
rect 35636 34066 35664 35634
rect 35624 34060 35676 34066
rect 35624 34002 35676 34008
rect 35728 33998 35756 35799
rect 35820 35290 35848 39063
rect 35912 37262 35940 39200
rect 35992 37392 36044 37398
rect 35992 37334 36044 37340
rect 36280 37346 36308 39200
rect 35900 37256 35952 37262
rect 35900 37198 35952 37204
rect 35808 35284 35860 35290
rect 35808 35226 35860 35232
rect 35900 35080 35952 35086
rect 35900 35022 35952 35028
rect 35808 34400 35860 34406
rect 35808 34342 35860 34348
rect 35820 34241 35848 34342
rect 35806 34232 35862 34241
rect 35806 34167 35862 34176
rect 35912 34134 35940 35022
rect 35900 34128 35952 34134
rect 35900 34070 35952 34076
rect 35716 33992 35768 33998
rect 35716 33934 35768 33940
rect 35728 33658 35756 33934
rect 35716 33652 35768 33658
rect 35716 33594 35768 33600
rect 35912 31346 35940 34070
rect 35900 31340 35952 31346
rect 35900 31282 35952 31288
rect 35912 30938 35940 31282
rect 35900 30932 35952 30938
rect 35900 30874 35952 30880
rect 35912 28490 35940 30874
rect 35900 28484 35952 28490
rect 35900 28426 35952 28432
rect 35912 27538 35940 28426
rect 35900 27532 35952 27538
rect 35900 27474 35952 27480
rect 35912 26994 35940 27474
rect 35900 26988 35952 26994
rect 35900 26930 35952 26936
rect 35900 22704 35952 22710
rect 35900 22646 35952 22652
rect 35532 21140 35584 21146
rect 35532 21082 35584 21088
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35912 19718 35940 22646
rect 35900 19712 35952 19718
rect 35900 19654 35952 19660
rect 35912 19514 35940 19654
rect 35900 19508 35952 19514
rect 35900 19450 35952 19456
rect 34704 19440 34756 19446
rect 34704 19382 34756 19388
rect 34716 18970 34744 19382
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34612 17876 34664 17882
rect 34612 17818 34664 17824
rect 34808 15706 34836 19314
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 35360 15706 35388 15982
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 35348 15700 35400 15706
rect 35348 15642 35400 15648
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34808 14521 34836 15438
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34794 14512 34850 14521
rect 34716 14470 34794 14498
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34428 5364 34480 5370
rect 34428 5306 34480 5312
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34336 4004 34388 4010
rect 34336 3946 34388 3952
rect 34244 3936 34296 3942
rect 34244 3878 34296 3884
rect 34256 3738 34284 3878
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 34336 3392 34388 3398
rect 34336 3334 34388 3340
rect 34348 800 34376 3334
rect 34440 3126 34468 4014
rect 34532 3534 34560 6598
rect 34520 3528 34572 3534
rect 34520 3470 34572 3476
rect 34428 3120 34480 3126
rect 34428 3062 34480 3068
rect 34624 2446 34652 7142
rect 34716 2650 34744 14470
rect 34794 14447 34850 14456
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35348 11076 35400 11082
rect 35348 11018 35400 11024
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34796 8900 34848 8906
rect 34796 8842 34848 8848
rect 34808 5914 34836 8842
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34796 5908 34848 5914
rect 34796 5850 34848 5856
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35164 4548 35216 4554
rect 35164 4490 35216 4496
rect 35176 4049 35204 4490
rect 35162 4040 35218 4049
rect 35360 4026 35388 11018
rect 36004 10810 36032 37334
rect 36280 37318 36400 37346
rect 36266 37224 36322 37233
rect 36266 37159 36322 37168
rect 36280 37126 36308 37159
rect 36268 37120 36320 37126
rect 36268 37062 36320 37068
rect 36372 36922 36400 37318
rect 36360 36916 36412 36922
rect 36360 36858 36412 36864
rect 36268 36780 36320 36786
rect 36268 36722 36320 36728
rect 36280 34542 36308 36722
rect 36360 35692 36412 35698
rect 36360 35634 36412 35640
rect 36268 34536 36320 34542
rect 36268 34478 36320 34484
rect 36372 33318 36400 35634
rect 36556 35562 36584 39200
rect 36924 39114 36952 39200
rect 37016 39114 37044 39222
rect 36924 39086 37044 39114
rect 36634 37496 36690 37505
rect 36634 37431 36690 37440
rect 36544 35556 36596 35562
rect 36544 35498 36596 35504
rect 36452 35012 36504 35018
rect 36452 34954 36504 34960
rect 36360 33312 36412 33318
rect 36360 33254 36412 33260
rect 36268 32972 36320 32978
rect 36268 32914 36320 32920
rect 36176 31680 36228 31686
rect 36176 31622 36228 31628
rect 36188 31414 36216 31622
rect 36176 31408 36228 31414
rect 36176 31350 36228 31356
rect 36084 27872 36136 27878
rect 36084 27814 36136 27820
rect 36096 25294 36124 27814
rect 36280 26234 36308 32914
rect 36188 26206 36308 26234
rect 36084 25288 36136 25294
rect 36084 25230 36136 25236
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 36096 21010 36124 22374
rect 36084 21004 36136 21010
rect 36084 20946 36136 20952
rect 35992 10804 36044 10810
rect 35992 10746 36044 10752
rect 35808 8900 35860 8906
rect 35808 8842 35860 8848
rect 35820 8786 35848 8842
rect 35820 8758 36124 8786
rect 35820 8566 35848 8758
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35532 7744 35584 7750
rect 35532 7686 35584 7692
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35452 5710 35480 6734
rect 35544 6390 35572 7686
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35532 5840 35584 5846
rect 35532 5782 35584 5788
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 35438 5400 35494 5409
rect 35438 5335 35494 5344
rect 35452 5302 35480 5335
rect 35440 5296 35492 5302
rect 35440 5238 35492 5244
rect 35544 4146 35572 5782
rect 35636 4185 35664 6258
rect 35622 4176 35678 4185
rect 35532 4140 35584 4146
rect 35622 4111 35678 4120
rect 35532 4082 35584 4088
rect 35360 3998 35572 4026
rect 35162 3975 35218 3984
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 34808 2530 34836 3470
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34808 2502 34928 2530
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34624 800 34652 2382
rect 34900 800 34928 2502
rect 35360 1986 35388 3878
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 35176 1958 35388 1986
rect 35176 800 35204 1958
rect 35452 800 35480 3062
rect 35544 3058 35572 3998
rect 35624 4004 35676 4010
rect 35624 3946 35676 3952
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35636 2854 35664 3946
rect 35728 3126 35756 7822
rect 35900 7200 35952 7206
rect 35900 7142 35952 7148
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35820 5642 35848 6598
rect 35808 5636 35860 5642
rect 35808 5578 35860 5584
rect 35716 3120 35768 3126
rect 35716 3062 35768 3068
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 35624 2848 35676 2854
rect 35624 2790 35676 2796
rect 35728 800 35756 2858
rect 35912 2514 35940 7142
rect 35992 6112 36044 6118
rect 35992 6054 36044 6060
rect 36004 4758 36032 6054
rect 36096 5914 36124 8758
rect 36188 8090 36216 26206
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36176 8084 36228 8090
rect 36176 8026 36228 8032
rect 36176 7336 36228 7342
rect 36176 7278 36228 7284
rect 36188 6322 36216 7278
rect 36176 6316 36228 6322
rect 36176 6258 36228 6264
rect 36084 5908 36136 5914
rect 36084 5850 36136 5856
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 35992 4752 36044 4758
rect 35992 4694 36044 4700
rect 36096 4622 36124 5510
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 35992 4480 36044 4486
rect 35992 4422 36044 4428
rect 35900 2508 35952 2514
rect 35900 2450 35952 2456
rect 36004 800 36032 4422
rect 36280 4214 36308 8298
rect 36268 4208 36320 4214
rect 36268 4150 36320 4156
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 36188 2106 36216 2382
rect 36176 2100 36228 2106
rect 36176 2042 36228 2048
rect 36280 800 36308 4150
rect 36372 2922 36400 33254
rect 36464 31686 36492 34954
rect 36648 34746 36676 37431
rect 37200 37244 37228 39222
rect 37278 39200 37334 40000
rect 37646 39200 37702 40000
rect 38014 39200 38070 40000
rect 38290 39200 38346 40000
rect 38658 39200 38714 40000
rect 39026 39200 39082 40000
rect 39394 39200 39450 40000
rect 39762 39200 39818 40000
rect 37292 37618 37320 39200
rect 37292 37590 37412 37618
rect 37280 37256 37332 37262
rect 37200 37216 37280 37244
rect 37280 37198 37332 37204
rect 37292 35834 37320 37198
rect 37280 35828 37332 35834
rect 37280 35770 37332 35776
rect 37384 35562 37412 37590
rect 37556 36712 37608 36718
rect 37556 36654 37608 36660
rect 37568 36242 37596 36654
rect 37556 36236 37608 36242
rect 37556 36178 37608 36184
rect 37372 35556 37424 35562
rect 37372 35498 37424 35504
rect 37280 35080 37332 35086
rect 37280 35022 37332 35028
rect 37292 34746 37320 35022
rect 36636 34740 36688 34746
rect 36636 34682 36688 34688
rect 37280 34740 37332 34746
rect 37280 34682 37332 34688
rect 37188 34672 37240 34678
rect 37188 34614 37240 34620
rect 37096 34536 37148 34542
rect 37096 34478 37148 34484
rect 36636 33992 36688 33998
rect 36556 33952 36636 33980
rect 36556 32774 36584 33952
rect 36636 33934 36688 33940
rect 37108 32978 37136 34478
rect 37200 34202 37228 34614
rect 37556 34604 37608 34610
rect 37556 34546 37608 34552
rect 37188 34196 37240 34202
rect 37188 34138 37240 34144
rect 37096 32972 37148 32978
rect 37096 32914 37148 32920
rect 36544 32768 36596 32774
rect 36544 32710 36596 32716
rect 36452 31680 36504 31686
rect 36452 31622 36504 31628
rect 36464 31346 36492 31622
rect 36452 31340 36504 31346
rect 36452 31282 36504 31288
rect 36556 15162 36584 32710
rect 37568 27606 37596 34546
rect 37660 34202 37688 39200
rect 38028 36854 38056 39200
rect 38016 36848 38068 36854
rect 38016 36790 38068 36796
rect 37924 35692 37976 35698
rect 37924 35634 37976 35640
rect 37832 35556 37884 35562
rect 37832 35498 37884 35504
rect 37648 34196 37700 34202
rect 37648 34138 37700 34144
rect 37556 27600 37608 27606
rect 37556 27542 37608 27548
rect 37188 26784 37240 26790
rect 37188 26726 37240 26732
rect 36636 23656 36688 23662
rect 36636 23598 36688 23604
rect 36648 22710 36676 23598
rect 37096 22772 37148 22778
rect 37096 22714 37148 22720
rect 36636 22704 36688 22710
rect 36636 22646 36688 22652
rect 37108 21962 37136 22714
rect 37096 21956 37148 21962
rect 37096 21898 37148 21904
rect 37096 20936 37148 20942
rect 37096 20878 37148 20884
rect 36636 15428 36688 15434
rect 36636 15370 36688 15376
rect 36544 15156 36596 15162
rect 36544 15098 36596 15104
rect 36452 8832 36504 8838
rect 36452 8774 36504 8780
rect 36464 5234 36492 8774
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36452 5228 36504 5234
rect 36452 5170 36504 5176
rect 36556 3534 36584 7686
rect 36648 5710 36676 15370
rect 36728 10464 36780 10470
rect 36728 10406 36780 10412
rect 36740 6866 36768 10406
rect 37004 9988 37056 9994
rect 37004 9930 37056 9936
rect 36728 6860 36780 6866
rect 36728 6802 36780 6808
rect 36728 6316 36780 6322
rect 36728 6258 36780 6264
rect 36636 5704 36688 5710
rect 36636 5646 36688 5652
rect 36740 3942 36768 6258
rect 36820 5024 36872 5030
rect 36820 4966 36872 4972
rect 36728 3936 36780 3942
rect 36728 3878 36780 3884
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36360 2916 36412 2922
rect 36360 2858 36412 2864
rect 36464 2582 36492 2994
rect 36452 2576 36504 2582
rect 36452 2518 36504 2524
rect 36544 2508 36596 2514
rect 36544 2450 36596 2456
rect 36556 800 36584 2450
rect 36832 800 36860 4966
rect 37016 4758 37044 9930
rect 37108 5710 37136 20878
rect 37200 15502 37228 26726
rect 37568 26234 37596 27542
rect 37568 26206 37780 26234
rect 37752 23866 37780 26206
rect 37740 23860 37792 23866
rect 37740 23802 37792 23808
rect 37556 23724 37608 23730
rect 37556 23666 37608 23672
rect 37568 23118 37596 23666
rect 37556 23112 37608 23118
rect 37556 23054 37608 23060
rect 37568 20346 37596 23054
rect 37648 22976 37700 22982
rect 37648 22918 37700 22924
rect 37660 22642 37688 22918
rect 37648 22636 37700 22642
rect 37648 22578 37700 22584
rect 37660 20482 37688 22578
rect 37740 21888 37792 21894
rect 37740 21830 37792 21836
rect 37752 20602 37780 21830
rect 37740 20596 37792 20602
rect 37740 20538 37792 20544
rect 37660 20454 37780 20482
rect 37568 20318 37688 20346
rect 37372 18896 37424 18902
rect 37372 18838 37424 18844
rect 37280 18420 37332 18426
rect 37280 18362 37332 18368
rect 37188 15496 37240 15502
rect 37188 15438 37240 15444
rect 37292 14498 37320 18362
rect 37384 15162 37412 18838
rect 37556 17060 37608 17066
rect 37556 17002 37608 17008
rect 37464 16448 37516 16454
rect 37464 16390 37516 16396
rect 37476 16182 37504 16390
rect 37464 16176 37516 16182
rect 37464 16118 37516 16124
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 37568 14498 37596 17002
rect 37292 14470 37412 14498
rect 37280 14408 37332 14414
rect 37280 14350 37332 14356
rect 37292 14249 37320 14350
rect 37278 14240 37334 14249
rect 37278 14175 37334 14184
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 37292 11082 37320 14010
rect 37280 11076 37332 11082
rect 37280 11018 37332 11024
rect 37384 10810 37412 14470
rect 37476 14470 37596 14498
rect 37372 10804 37424 10810
rect 37372 10746 37424 10752
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 37188 7404 37240 7410
rect 37188 7346 37240 7352
rect 37200 6066 37228 7346
rect 37292 6186 37320 10610
rect 37476 9382 37504 14470
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37568 13326 37596 14350
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 37464 9376 37516 9382
rect 37464 9318 37516 9324
rect 37464 8356 37516 8362
rect 37464 8298 37516 8304
rect 37372 6792 37424 6798
rect 37372 6734 37424 6740
rect 37384 6322 37412 6734
rect 37372 6316 37424 6322
rect 37372 6258 37424 6264
rect 37280 6180 37332 6186
rect 37280 6122 37332 6128
rect 37200 6038 37320 6066
rect 37096 5704 37148 5710
rect 37096 5646 37148 5652
rect 37004 4752 37056 4758
rect 37004 4694 37056 4700
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 37096 4004 37148 4010
rect 37096 3946 37148 3952
rect 37108 800 37136 3946
rect 37200 2553 37228 4558
rect 37186 2544 37242 2553
rect 37292 2514 37320 6038
rect 37372 4548 37424 4554
rect 37372 4490 37424 4496
rect 37384 4010 37412 4490
rect 37372 4004 37424 4010
rect 37372 3946 37424 3952
rect 37476 3058 37504 8298
rect 37556 5568 37608 5574
rect 37556 5510 37608 5516
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37476 2774 37504 2994
rect 37384 2746 37504 2774
rect 37568 2774 37596 5510
rect 37660 3602 37688 20318
rect 37752 14074 37780 20454
rect 37740 14068 37792 14074
rect 37740 14010 37792 14016
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37752 13258 37780 13874
rect 37740 13252 37792 13258
rect 37740 13194 37792 13200
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 37752 6458 37780 9522
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37844 6390 37872 35498
rect 37936 33658 37964 35634
rect 38028 34746 38056 36790
rect 38200 36644 38252 36650
rect 38200 36586 38252 36592
rect 38016 34740 38068 34746
rect 38016 34682 38068 34688
rect 38016 33992 38068 33998
rect 38016 33934 38068 33940
rect 37924 33652 37976 33658
rect 37924 33594 37976 33600
rect 38028 32230 38056 33934
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38120 32502 38148 32846
rect 38108 32496 38160 32502
rect 38106 32464 38108 32473
rect 38160 32464 38162 32473
rect 38106 32399 38162 32408
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 37924 30592 37976 30598
rect 37924 30534 37976 30540
rect 37936 29850 37964 30534
rect 37924 29844 37976 29850
rect 37924 29786 37976 29792
rect 38028 26234 38056 32166
rect 38108 31340 38160 31346
rect 38108 31282 38160 31288
rect 38120 30841 38148 31282
rect 38212 31090 38240 36586
rect 38304 35290 38332 39200
rect 38384 37188 38436 37194
rect 38384 37130 38436 37136
rect 38292 35284 38344 35290
rect 38292 35226 38344 35232
rect 38212 31062 38332 31090
rect 38106 30832 38162 30841
rect 38106 30767 38162 30776
rect 38108 29640 38160 29646
rect 38108 29582 38160 29588
rect 38120 29209 38148 29582
rect 38106 29200 38162 29209
rect 38106 29135 38162 29144
rect 38108 28076 38160 28082
rect 38108 28018 38160 28024
rect 38120 27577 38148 28018
rect 38106 27568 38162 27577
rect 38106 27503 38162 27512
rect 38028 26206 38240 26234
rect 38106 25800 38162 25809
rect 38106 25735 38108 25744
rect 38160 25735 38162 25744
rect 38108 25706 38160 25712
rect 38014 24168 38070 24177
rect 38014 24103 38016 24112
rect 38068 24103 38070 24112
rect 38016 24074 38068 24080
rect 38106 22536 38162 22545
rect 38106 22471 38162 22480
rect 38120 22030 38148 22471
rect 38108 22024 38160 22030
rect 38108 21966 38160 21972
rect 38106 20904 38162 20913
rect 38106 20839 38162 20848
rect 38120 20466 38148 20839
rect 38108 20460 38160 20466
rect 38108 20402 38160 20408
rect 38106 19136 38162 19145
rect 38106 19071 38162 19080
rect 38120 18766 38148 19071
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 37924 18624 37976 18630
rect 37924 18566 37976 18572
rect 37936 16574 37964 18566
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 38120 17513 38148 17614
rect 38106 17504 38162 17513
rect 38106 17439 38162 17448
rect 37936 16546 38056 16574
rect 38028 16250 38056 16546
rect 38016 16244 38068 16250
rect 38016 16186 38068 16192
rect 38014 15872 38070 15881
rect 38014 15807 38070 15816
rect 38028 15502 38056 15807
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 38028 15162 38056 15438
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 38108 12640 38160 12646
rect 38108 12582 38160 12588
rect 38120 12481 38148 12582
rect 38106 12472 38162 12481
rect 38106 12407 38162 12416
rect 37924 12096 37976 12102
rect 37924 12038 37976 12044
rect 37936 11354 37964 12038
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 38108 11144 38160 11150
rect 38108 11086 38160 11092
rect 38120 10849 38148 11086
rect 38106 10840 38162 10849
rect 38106 10775 38162 10784
rect 38106 9208 38162 9217
rect 38106 9143 38162 9152
rect 38120 8974 38148 9143
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 37924 8424 37976 8430
rect 37924 8366 37976 8372
rect 37832 6384 37884 6390
rect 37832 6326 37884 6332
rect 37740 6112 37792 6118
rect 37740 6054 37792 6060
rect 37752 5778 37780 6054
rect 37740 5772 37792 5778
rect 37740 5714 37792 5720
rect 37844 5370 37872 6326
rect 37832 5364 37884 5370
rect 37832 5306 37884 5312
rect 37936 4554 37964 8366
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 38120 7585 38148 7822
rect 38106 7576 38162 7585
rect 38106 7511 38162 7520
rect 38108 7200 38160 7206
rect 38108 7142 38160 7148
rect 38014 5808 38070 5817
rect 38014 5743 38070 5752
rect 38028 5642 38056 5743
rect 38016 5636 38068 5642
rect 38016 5578 38068 5584
rect 38120 5234 38148 7142
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 37648 3596 37700 3602
rect 37648 3538 37700 3544
rect 37568 2746 37688 2774
rect 37186 2479 37242 2488
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37384 800 37412 2746
rect 37660 800 37688 2746
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 37936 800 37964 2382
rect 38120 921 38148 5170
rect 38212 4010 38240 26206
rect 38304 8634 38332 31062
rect 38292 8628 38344 8634
rect 38292 8570 38344 8576
rect 38304 7478 38332 8570
rect 38292 7472 38344 7478
rect 38292 7414 38344 7420
rect 38396 4146 38424 37130
rect 38568 36168 38620 36174
rect 38568 36110 38620 36116
rect 38476 33924 38528 33930
rect 38476 33866 38528 33872
rect 38488 22778 38516 33866
rect 38476 22772 38528 22778
rect 38476 22714 38528 22720
rect 38580 19310 38608 36110
rect 38672 33658 38700 39200
rect 38844 36100 38896 36106
rect 38844 36042 38896 36048
rect 38752 35080 38804 35086
rect 38752 35022 38804 35028
rect 38660 33652 38712 33658
rect 38660 33594 38712 33600
rect 38764 33538 38792 35022
rect 38672 33510 38792 33538
rect 38568 19304 38620 19310
rect 38568 19246 38620 19252
rect 38476 15020 38528 15026
rect 38476 14962 38528 14968
rect 38488 6798 38516 14962
rect 38672 14006 38700 33510
rect 38752 33448 38804 33454
rect 38752 33390 38804 33396
rect 38764 16182 38792 33390
rect 38856 23594 38884 36042
rect 39040 35698 39068 39200
rect 39028 35692 39080 35698
rect 39028 35634 39080 35640
rect 39408 34542 39436 39200
rect 39776 34678 39804 39200
rect 39764 34672 39816 34678
rect 39764 34614 39816 34620
rect 39396 34536 39448 34542
rect 39396 34478 39448 34484
rect 38844 23588 38896 23594
rect 38844 23530 38896 23536
rect 38844 19372 38896 19378
rect 38844 19314 38896 19320
rect 38752 16176 38804 16182
rect 38752 16118 38804 16124
rect 38660 14000 38712 14006
rect 38660 13942 38712 13948
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 38200 4004 38252 4010
rect 38200 3946 38252 3952
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 38106 912 38162 921
rect 38106 847 38162 856
rect 38212 800 38240 3470
rect 38396 3466 38424 4082
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38488 800 38516 6598
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 38764 800 38792 2926
rect 38856 2514 38884 19314
rect 39580 6316 39632 6322
rect 39580 6258 39632 6264
rect 39304 5840 39356 5846
rect 39304 5782 39356 5788
rect 39028 3936 39080 3942
rect 39028 3878 39080 3884
rect 38844 2508 38896 2514
rect 38844 2450 38896 2456
rect 39040 800 39068 3878
rect 39316 800 39344 5782
rect 39592 800 39620 6258
rect 39856 6248 39908 6254
rect 39856 6190 39908 6196
rect 39868 800 39896 6190
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
<< via2 >>
rect 1582 29960 1638 30016
rect 3146 9968 3202 10024
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4434 3440 4490 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5078 4004 5134 4040
rect 5078 3984 5080 4004
rect 5080 3984 5132 4004
rect 5132 3984 5134 4004
rect 5538 3304 5594 3360
rect 6274 3460 6330 3496
rect 6274 3440 6276 3460
rect 6276 3440 6328 3460
rect 6328 3440 6330 3460
rect 7470 36216 7526 36272
rect 7562 3440 7618 3496
rect 7930 4120 7986 4176
rect 8298 3712 8354 3768
rect 8298 3168 8354 3224
rect 8390 3052 8446 3088
rect 8390 3032 8392 3052
rect 8392 3032 8444 3052
rect 8444 3032 8446 3052
rect 12070 36100 12126 36136
rect 12070 36080 12072 36100
rect 12072 36080 12124 36100
rect 12124 36080 12126 36100
rect 11334 30252 11390 30288
rect 11334 30232 11336 30252
rect 11336 30232 11388 30252
rect 11388 30232 11390 30252
rect 12990 30268 12992 30288
rect 12992 30268 13044 30288
rect 13044 30268 13046 30288
rect 12990 30232 13046 30268
rect 8942 3576 8998 3632
rect 11518 3168 11574 3224
rect 11978 3168 12034 3224
rect 12714 3712 12770 3768
rect 13634 3168 13690 3224
rect 14278 2352 14334 2408
rect 14554 3460 14610 3496
rect 14554 3440 14556 3460
rect 14556 3440 14608 3460
rect 14608 3440 14610 3460
rect 16026 3340 16028 3360
rect 16028 3340 16080 3360
rect 16080 3340 16082 3360
rect 16026 3304 16082 3340
rect 16394 3984 16450 4040
rect 16302 3576 16358 3632
rect 16486 3032 16542 3088
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19062 4120 19118 4176
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19890 2488 19946 2544
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20166 4528 20222 4584
rect 20810 14476 20866 14512
rect 20810 14456 20812 14476
rect 20812 14456 20864 14476
rect 20864 14456 20866 14476
rect 22558 3984 22614 4040
rect 23386 3848 23442 3904
rect 25226 2352 25282 2408
rect 28078 37168 28134 37224
rect 27158 2488 27214 2544
rect 27894 5344 27950 5400
rect 29366 36080 29422 36136
rect 30194 36216 30250 36272
rect 30286 3848 30342 3904
rect 33046 3460 33102 3496
rect 33046 3440 33048 3460
rect 33048 3440 33100 3460
rect 33100 3440 33102 3460
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35806 39072 35862 39128
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35714 35808 35770 35864
rect 35806 34176 35862 34232
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34794 14456 34850 14512
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35162 3984 35218 4040
rect 36266 37168 36322 37224
rect 36634 37440 36690 37496
rect 35438 5344 35494 5400
rect 35622 4120 35678 4176
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37278 14184 37334 14240
rect 37186 2488 37242 2544
rect 38106 32444 38108 32464
rect 38108 32444 38160 32464
rect 38160 32444 38162 32464
rect 38106 32408 38162 32444
rect 38106 30776 38162 30832
rect 38106 29144 38162 29200
rect 38106 27512 38162 27568
rect 38106 25764 38162 25800
rect 38106 25744 38108 25764
rect 38108 25744 38160 25764
rect 38160 25744 38162 25764
rect 38014 24132 38070 24168
rect 38014 24112 38016 24132
rect 38016 24112 38068 24132
rect 38068 24112 38070 24132
rect 38106 22480 38162 22536
rect 38106 20848 38162 20904
rect 38106 19080 38162 19136
rect 38106 17448 38162 17504
rect 38014 15816 38070 15872
rect 38106 12416 38162 12472
rect 38106 10784 38162 10840
rect 38106 9152 38162 9208
rect 38106 7520 38162 7576
rect 38014 5752 38070 5808
rect 38106 856 38162 912
<< metal3 >>
rect 35801 39130 35867 39133
rect 39200 39130 40000 39160
rect 35801 39128 40000 39130
rect 35801 39072 35806 39128
rect 35862 39072 40000 39128
rect 35801 39070 40000 39072
rect 35801 39067 35867 39070
rect 39200 39040 40000 39070
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 36629 37498 36695 37501
rect 39200 37498 40000 37528
rect 36629 37496 40000 37498
rect 36629 37440 36634 37496
rect 36690 37440 40000 37496
rect 36629 37438 40000 37440
rect 36629 37435 36695 37438
rect 39200 37408 40000 37438
rect 28073 37226 28139 37229
rect 36261 37226 36327 37229
rect 28073 37224 36327 37226
rect 28073 37168 28078 37224
rect 28134 37168 36266 37224
rect 36322 37168 36327 37224
rect 28073 37166 36327 37168
rect 28073 37163 28139 37166
rect 36261 37163 36327 37166
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 7465 36274 7531 36277
rect 30189 36274 30255 36277
rect 7465 36272 30255 36274
rect 7465 36216 7470 36272
rect 7526 36216 30194 36272
rect 30250 36216 30255 36272
rect 7465 36214 30255 36216
rect 7465 36211 7531 36214
rect 30189 36211 30255 36214
rect 12065 36138 12131 36141
rect 29361 36138 29427 36141
rect 12065 36136 29427 36138
rect 12065 36080 12070 36136
rect 12126 36080 29366 36136
rect 29422 36080 29427 36136
rect 12065 36078 29427 36080
rect 12065 36075 12131 36078
rect 29361 36075 29427 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 35709 35866 35775 35869
rect 39200 35866 40000 35896
rect 35709 35864 40000 35866
rect 35709 35808 35714 35864
rect 35770 35808 40000 35864
rect 35709 35806 40000 35808
rect 35709 35803 35775 35806
rect 39200 35776 40000 35806
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 35801 34234 35867 34237
rect 39200 34234 40000 34264
rect 35801 34232 40000 34234
rect 35801 34176 35806 34232
rect 35862 34176 40000 34232
rect 35801 34174 40000 34176
rect 35801 34171 35867 34174
rect 39200 34144 40000 34174
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 38101 32466 38167 32469
rect 39200 32466 40000 32496
rect 38101 32464 40000 32466
rect 38101 32408 38106 32464
rect 38162 32408 40000 32464
rect 38101 32406 40000 32408
rect 38101 32403 38167 32406
rect 39200 32376 40000 32406
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 38101 30834 38167 30837
rect 39200 30834 40000 30864
rect 38101 30832 40000 30834
rect 38101 30776 38106 30832
rect 38162 30776 40000 30832
rect 38101 30774 40000 30776
rect 38101 30771 38167 30774
rect 39200 30744 40000 30774
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 11329 30290 11395 30293
rect 12985 30290 13051 30293
rect 11329 30288 13051 30290
rect 11329 30232 11334 30288
rect 11390 30232 12990 30288
rect 13046 30232 13051 30288
rect 11329 30230 13051 30232
rect 11329 30227 11395 30230
rect 12985 30227 13051 30230
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 38101 29202 38167 29205
rect 39200 29202 40000 29232
rect 38101 29200 40000 29202
rect 38101 29144 38106 29200
rect 38162 29144 40000 29200
rect 38101 29142 40000 29144
rect 38101 29139 38167 29142
rect 39200 29112 40000 29142
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 38101 27570 38167 27573
rect 39200 27570 40000 27600
rect 38101 27568 40000 27570
rect 38101 27512 38106 27568
rect 38162 27512 40000 27568
rect 38101 27510 40000 27512
rect 38101 27507 38167 27510
rect 39200 27480 40000 27510
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 38101 25802 38167 25805
rect 39200 25802 40000 25832
rect 38101 25800 40000 25802
rect 38101 25744 38106 25800
rect 38162 25744 40000 25800
rect 38101 25742 40000 25744
rect 38101 25739 38167 25742
rect 39200 25712 40000 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 38009 24170 38075 24173
rect 39200 24170 40000 24200
rect 38009 24168 40000 24170
rect 38009 24112 38014 24168
rect 38070 24112 40000 24168
rect 38009 24110 40000 24112
rect 38009 24107 38075 24110
rect 39200 24080 40000 24110
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 38101 22538 38167 22541
rect 39200 22538 40000 22568
rect 38101 22536 40000 22538
rect 38101 22480 38106 22536
rect 38162 22480 40000 22536
rect 38101 22478 40000 22480
rect 38101 22475 38167 22478
rect 39200 22448 40000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 38101 20906 38167 20909
rect 39200 20906 40000 20936
rect 38101 20904 40000 20906
rect 38101 20848 38106 20904
rect 38162 20848 40000 20904
rect 38101 20846 40000 20848
rect 38101 20843 38167 20846
rect 39200 20816 40000 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 38101 19138 38167 19141
rect 39200 19138 40000 19168
rect 38101 19136 40000 19138
rect 38101 19080 38106 19136
rect 38162 19080 40000 19136
rect 38101 19078 40000 19080
rect 38101 19075 38167 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 39200 19048 40000 19078
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 38101 17506 38167 17509
rect 39200 17506 40000 17536
rect 38101 17504 40000 17506
rect 38101 17448 38106 17504
rect 38162 17448 40000 17504
rect 38101 17446 40000 17448
rect 38101 17443 38167 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 39200 17416 40000 17446
rect 19568 17375 19888 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 38009 15874 38075 15877
rect 39200 15874 40000 15904
rect 38009 15872 40000 15874
rect 38009 15816 38014 15872
rect 38070 15816 40000 15872
rect 38009 15814 40000 15816
rect 38009 15811 38075 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 39200 15784 40000 15814
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 20805 14514 20871 14517
rect 34789 14514 34855 14517
rect 20805 14512 34855 14514
rect 20805 14456 20810 14512
rect 20866 14456 34794 14512
rect 34850 14456 34855 14512
rect 20805 14454 34855 14456
rect 20805 14451 20871 14454
rect 34789 14451 34855 14454
rect 37273 14242 37339 14245
rect 39200 14242 40000 14272
rect 37273 14240 40000 14242
rect 37273 14184 37278 14240
rect 37334 14184 40000 14240
rect 37273 14182 40000 14184
rect 37273 14179 37339 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 39200 14152 40000 14182
rect 19568 14111 19888 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 38101 12474 38167 12477
rect 39200 12474 40000 12504
rect 38101 12472 40000 12474
rect 38101 12416 38106 12472
rect 38162 12416 40000 12472
rect 38101 12414 40000 12416
rect 38101 12411 38167 12414
rect 39200 12384 40000 12414
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 38101 10842 38167 10845
rect 39200 10842 40000 10872
rect 38101 10840 40000 10842
rect 38101 10784 38106 10840
rect 38162 10784 40000 10840
rect 38101 10782 40000 10784
rect 38101 10779 38167 10782
rect 39200 10752 40000 10782
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 0 10026 800 10056
rect 3141 10026 3207 10029
rect 0 10024 3207 10026
rect 0 9968 3146 10024
rect 3202 9968 3207 10024
rect 0 9966 3207 9968
rect 0 9936 800 9966
rect 3141 9963 3207 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 38101 9210 38167 9213
rect 39200 9210 40000 9240
rect 38101 9208 40000 9210
rect 38101 9152 38106 9208
rect 38162 9152 40000 9208
rect 38101 9150 40000 9152
rect 38101 9147 38167 9150
rect 39200 9120 40000 9150
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 38101 7578 38167 7581
rect 39200 7578 40000 7608
rect 38101 7576 40000 7578
rect 38101 7520 38106 7576
rect 38162 7520 40000 7576
rect 38101 7518 40000 7520
rect 38101 7515 38167 7518
rect 39200 7488 40000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 38009 5810 38075 5813
rect 39200 5810 40000 5840
rect 38009 5808 40000 5810
rect 38009 5752 38014 5808
rect 38070 5752 40000 5808
rect 38009 5750 40000 5752
rect 38009 5747 38075 5750
rect 39200 5720 40000 5750
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 27889 5402 27955 5405
rect 35433 5402 35499 5405
rect 27889 5400 35499 5402
rect 27889 5344 27894 5400
rect 27950 5344 35438 5400
rect 35494 5344 35499 5400
rect 27889 5342 35499 5344
rect 27889 5339 27955 5342
rect 35433 5339 35499 5342
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 20161 4586 20227 4589
rect 20118 4584 20227 4586
rect 20118 4528 20166 4584
rect 20222 4528 20227 4584
rect 20118 4523 20227 4528
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 7925 4178 7991 4181
rect 19057 4178 19123 4181
rect 20118 4178 20178 4523
rect 7925 4176 20178 4178
rect 7925 4120 7930 4176
rect 7986 4120 19062 4176
rect 19118 4120 20178 4176
rect 7925 4118 20178 4120
rect 35617 4178 35683 4181
rect 39200 4178 40000 4208
rect 35617 4176 40000 4178
rect 35617 4120 35622 4176
rect 35678 4120 40000 4176
rect 35617 4118 40000 4120
rect 7925 4115 7991 4118
rect 19057 4115 19123 4118
rect 35617 4115 35683 4118
rect 39200 4088 40000 4118
rect 5073 4042 5139 4045
rect 16389 4042 16455 4045
rect 5073 4040 16455 4042
rect 5073 3984 5078 4040
rect 5134 3984 16394 4040
rect 16450 3984 16455 4040
rect 5073 3982 16455 3984
rect 5073 3979 5139 3982
rect 16389 3979 16455 3982
rect 22553 4042 22619 4045
rect 35157 4042 35223 4045
rect 22553 4040 35223 4042
rect 22553 3984 22558 4040
rect 22614 3984 35162 4040
rect 35218 3984 35223 4040
rect 22553 3982 35223 3984
rect 22553 3979 22619 3982
rect 35157 3979 35223 3982
rect 23381 3906 23447 3909
rect 30281 3906 30347 3909
rect 23381 3904 30347 3906
rect 23381 3848 23386 3904
rect 23442 3848 30286 3904
rect 30342 3848 30347 3904
rect 23381 3846 30347 3848
rect 23381 3843 23447 3846
rect 30281 3843 30347 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 8293 3770 8359 3773
rect 12709 3770 12775 3773
rect 8293 3768 12775 3770
rect 8293 3712 8298 3768
rect 8354 3712 12714 3768
rect 12770 3712 12775 3768
rect 8293 3710 12775 3712
rect 8293 3707 8359 3710
rect 12709 3707 12775 3710
rect 8937 3634 9003 3637
rect 16297 3634 16363 3637
rect 8937 3632 16363 3634
rect 8937 3576 8942 3632
rect 8998 3576 16302 3632
rect 16358 3576 16363 3632
rect 8937 3574 16363 3576
rect 8937 3571 9003 3574
rect 16297 3571 16363 3574
rect 4429 3498 4495 3501
rect 6269 3498 6335 3501
rect 4429 3496 6335 3498
rect 4429 3440 4434 3496
rect 4490 3440 6274 3496
rect 6330 3440 6335 3496
rect 4429 3438 6335 3440
rect 4429 3435 4495 3438
rect 6269 3435 6335 3438
rect 7557 3498 7623 3501
rect 14549 3498 14615 3501
rect 33041 3498 33107 3501
rect 7557 3496 14615 3498
rect 7557 3440 7562 3496
rect 7618 3440 14554 3496
rect 14610 3440 14615 3496
rect 7557 3438 14615 3440
rect 7557 3435 7623 3438
rect 14549 3435 14615 3438
rect 16254 3496 33107 3498
rect 16254 3440 33046 3496
rect 33102 3440 33107 3496
rect 16254 3438 33107 3440
rect 5533 3362 5599 3365
rect 16021 3362 16087 3365
rect 5533 3360 16087 3362
rect 5533 3304 5538 3360
rect 5594 3304 16026 3360
rect 16082 3304 16087 3360
rect 5533 3302 16087 3304
rect 5533 3299 5599 3302
rect 16021 3299 16087 3302
rect 8293 3226 8359 3229
rect 11513 3226 11579 3229
rect 11973 3226 12039 3229
rect 8293 3224 12039 3226
rect 8293 3168 8298 3224
rect 8354 3168 11518 3224
rect 11574 3168 11978 3224
rect 12034 3168 12039 3224
rect 8293 3166 12039 3168
rect 8293 3163 8359 3166
rect 11513 3163 11579 3166
rect 11973 3163 12039 3166
rect 13629 3226 13695 3229
rect 16254 3226 16314 3438
rect 33041 3435 33107 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 13629 3224 16314 3226
rect 13629 3168 13634 3224
rect 13690 3168 16314 3224
rect 13629 3166 16314 3168
rect 13629 3163 13695 3166
rect 8385 3090 8451 3093
rect 16481 3090 16547 3093
rect 8385 3088 16547 3090
rect 8385 3032 8390 3088
rect 8446 3032 16486 3088
rect 16542 3032 16547 3088
rect 8385 3030 16547 3032
rect 8385 3027 8451 3030
rect 16481 3027 16547 3030
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 19885 2546 19951 2549
rect 27153 2546 27219 2549
rect 19885 2544 27219 2546
rect 19885 2488 19890 2544
rect 19946 2488 27158 2544
rect 27214 2488 27219 2544
rect 19885 2486 27219 2488
rect 19885 2483 19951 2486
rect 27153 2483 27219 2486
rect 37181 2546 37247 2549
rect 39200 2546 40000 2576
rect 37181 2544 40000 2546
rect 37181 2488 37186 2544
rect 37242 2488 40000 2544
rect 37181 2486 40000 2488
rect 37181 2483 37247 2486
rect 39200 2456 40000 2486
rect 14273 2410 14339 2413
rect 25221 2410 25287 2413
rect 14273 2408 25287 2410
rect 14273 2352 14278 2408
rect 14334 2352 25226 2408
rect 25282 2352 25287 2408
rect 14273 2350 25287 2352
rect 14273 2347 14339 2350
rect 25221 2347 25287 2350
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 38101 914 38167 917
rect 39200 914 40000 944
rect 38101 912 40000 914
rect 38101 856 38106 912
rect 38162 856 40000 912
rect 38101 854 40000 856
rect 38101 851 38167 854
rect 39200 824 40000 854
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1644511149
transform -1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B
timestamp 1644511149
transform 1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__B
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__B
timestamp 1644511149
transform -1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1644511149
transform -1 0 24564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1644511149
transform -1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1644511149
transform -1 0 23368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__B
timestamp 1644511149
transform -1 0 32568 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__B
timestamp 1644511149
transform -1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A_N
timestamp 1644511149
transform -1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B
timestamp 1644511149
transform -1 0 21712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A_N
timestamp 1644511149
transform 1 0 24472 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A_N
timestamp 1644511149
transform -1 0 29716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__B
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A_N
timestamp 1644511149
transform 1 0 24840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B
timestamp 1644511149
transform 1 0 23368 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B
timestamp 1644511149
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__B
timestamp 1644511149
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1644511149
transform -1 0 26496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B
timestamp 1644511149
transform -1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1644511149
transform -1 0 26496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__B
timestamp 1644511149
transform -1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1644511149
transform -1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 1644511149
transform -1 0 27140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__B
timestamp 1644511149
transform 1 0 27876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B
timestamp 1644511149
transform -1 0 27968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B
timestamp 1644511149
transform -1 0 31280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A_N
timestamp 1644511149
transform 1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__B
timestamp 1644511149
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1644511149
transform -1 0 34224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B
timestamp 1644511149
transform -1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B
timestamp 1644511149
transform -1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1644511149
transform -1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A_N
timestamp 1644511149
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__B
timestamp 1644511149
transform -1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1644511149
transform -1 0 36708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B
timestamp 1644511149
transform 1 0 35052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A_N
timestamp 1644511149
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1644511149
transform -1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__S
timestamp 1644511149
transform 1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1644511149
transform 1 0 3956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A0
timestamp 1644511149
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A0
timestamp 1644511149
transform -1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A0
timestamp 1644511149
transform -1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A0
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A0
timestamp 1644511149
transform -1 0 30176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A0
timestamp 1644511149
transform -1 0 32384 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A0
timestamp 1644511149
transform -1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1644511149
transform 1 0 12880 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1644511149
transform -1 0 34224 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A0
timestamp 1644511149
transform -1 0 13524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__S
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A0
timestamp 1644511149
transform -1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A0
timestamp 1644511149
transform -1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A0
timestamp 1644511149
transform -1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__S
timestamp 1644511149
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A0
timestamp 1644511149
transform -1 0 38180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A_N
timestamp 1644511149
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1644511149
transform -1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A0
timestamp 1644511149
transform -1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__S
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1644511149
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1644511149
transform -1 0 23920 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1644511149
transform -1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A0
timestamp 1644511149
transform -1 0 26680 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A0
timestamp 1644511149
transform -1 0 29072 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__B
timestamp 1644511149
transform -1 0 22448 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A0
timestamp 1644511149
transform 1 0 31464 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__B
timestamp 1644511149
transform -1 0 29716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A0
timestamp 1644511149
transform 1 0 33396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__S
timestamp 1644511149
transform -1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__S
timestamp 1644511149
transform -1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S
timestamp 1644511149
transform -1 0 23000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A_N
timestamp 1644511149
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1644511149
transform -1 0 3956 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1644511149
transform 1 0 11040 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A_N
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__B
timestamp 1644511149
transform 1 0 23552 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__B
timestamp 1644511149
transform -1 0 27876 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__B1
timestamp 1644511149
transform -1 0 31004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__B1
timestamp 1644511149
transform 1 0 31464 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1644511149
transform 1 0 26496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1644511149
transform -1 0 5888 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__B
timestamp 1644511149
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__B
timestamp 1644511149
transform -1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B
timestamp 1644511149
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1644511149
transform -1 0 4968 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__B
timestamp 1644511149
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1644511149
transform 1 0 7084 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__B
timestamp 1644511149
transform -1 0 30176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1644511149
transform -1 0 8188 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1644511149
transform -1 0 31372 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__B
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1644511149
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1644511149
transform 1 0 32936 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1644511149
transform 1 0 15640 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__B
timestamp 1644511149
transform -1 0 14812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1644511149
transform -1 0 15272 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__B
timestamp 1644511149
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1644511149
transform 1 0 14444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__B
timestamp 1644511149
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1644511149
transform -1 0 17112 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1644511149
transform -1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__B
timestamp 1644511149
transform -1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1644511149
transform -1 0 18124 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1644511149
transform 1 0 19688 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__B
timestamp 1644511149
transform -1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1644511149
transform 1 0 20700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1644511149
transform 1 0 11592 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1644511149
transform 1 0 13432 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1644511149
transform -1 0 15824 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1644511149
transform -1 0 16560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__B
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__B
timestamp 1644511149
transform -1 0 25760 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__B
timestamp 1644511149
transform -1 0 27600 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__B
timestamp 1644511149
transform -1 0 29900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1644511149
transform -1 0 24748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1644511149
transform 1 0 28244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1644511149
transform -1 0 35512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__B1
timestamp 1644511149
transform 1 0 33396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1644511149
transform 1 0 31464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__B1
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1644511149
transform 1 0 25668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__B1
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1644511149
transform 1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__B1_N
timestamp 1644511149
transform 1 0 9108 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__C1
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__B1
timestamp 1644511149
transform -1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1644511149
transform -1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1644511149
transform 1 0 6164 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1644511149
transform 1 0 5888 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1644511149
transform 1 0 5428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A
timestamp 1644511149
transform 1 0 7360 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__B1
timestamp 1644511149
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__A
timestamp 1644511149
transform 1 0 16008 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__B1
timestamp 1644511149
transform 1 0 19964 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__A
timestamp 1644511149
transform -1 0 23644 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__B1
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1644511149
transform 1 0 29624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1644511149
transform 1 0 27600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1644511149
transform -1 0 27784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1644511149
transform -1 0 23828 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1644511149
transform 1 0 16744 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1644511149
transform 1 0 15364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1644511149
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1644511149
transform 1 0 10488 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1644511149
transform 1 0 8372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1644511149
transform 1 0 3864 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1644511149
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1644511149
transform -1 0 8924 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1644511149
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1644511149
transform 1 0 4140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1644511149
transform 1 0 11224 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1644511149
transform 1 0 10488 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1644511149
transform 1 0 13524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1644511149
transform 1 0 17480 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1644511149
transform 1 0 35604 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1644511149
transform 1 0 33764 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1644511149
transform 1 0 35144 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__A
timestamp 1644511149
transform 1 0 2024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A
timestamp 1644511149
transform -1 0 29440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__A
timestamp 1644511149
transform 1 0 31188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A
timestamp 1644511149
transform -1 0 36156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__A
timestamp 1644511149
transform 1 0 36432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__A
timestamp 1644511149
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1644511149
transform -1 0 28796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1644511149
transform -1 0 38180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A
timestamp 1644511149
transform -1 0 38180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A
timestamp 1644511149
transform -1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__A
timestamp 1644511149
transform -1 0 37628 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__A
timestamp 1644511149
transform 1 0 37444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1644511149
transform -1 0 37628 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__A
timestamp 1644511149
transform 1 0 35880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1644511149
transform 1 0 10856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1644511149
transform -1 0 28336 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 33028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 33856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 34684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 35144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 36340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 34132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 33304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 36800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 28152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 28704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 28796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 29072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 29716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 30544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 32108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 34868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 25116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 32936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 34868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 36248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 37628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 36616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 35696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 35696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 27600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 28152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform -1 0 31096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 31648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 29992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 32292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 30728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 32752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 19688 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 20516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 21160 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 24380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 12420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 9476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 18308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 19044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 20516 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 21344 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 22172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1644511149
transform -1 0 23092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1644511149
transform -1 0 24656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1644511149
transform -1 0 23828 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1644511149
transform -1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1644511149
transform -1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1644511149
transform -1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1644511149
transform -1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1644511149
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1644511149
transform -1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1644511149
transform -1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1644511149
transform -1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1644511149
transform -1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1644511149
transform -1 0 1748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1644511149
transform -1 0 12328 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1644511149
transform -1 0 15180 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1644511149
transform -1 0 12880 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1644511149
transform -1 0 16100 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1644511149
transform -1 0 18584 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1644511149
transform -1 0 17664 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1644511149
transform -1 0 17020 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1644511149
transform -1 0 18216 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1644511149
transform -1 0 19412 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1644511149
transform -1 0 20148 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1644511149
transform -1 0 2300 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1644511149
transform -1 0 23828 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1644511149
transform -1 0 22632 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1644511149
transform -1 0 23920 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1644511149
transform -1 0 24472 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1644511149
transform -1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1644511149
transform -1 0 26036 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1644511149
transform -1 0 28980 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1644511149
transform -1 0 29716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1644511149
transform -1 0 31372 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1644511149
transform -1 0 29992 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1644511149
transform -1 0 2668 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1644511149
transform -1 0 34132 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1644511149
transform -1 0 33672 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1644511149
transform -1 0 35604 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1644511149
transform -1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1644511149
transform -1 0 38180 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1644511149
transform -1 0 37444 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1644511149
transform -1 0 37444 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1644511149
transform -1 0 37444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1644511149
transform -1 0 4692 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1644511149
transform -1 0 5244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1644511149
transform -1 0 6348 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1644511149
transform -1 0 6900 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1644511149
transform -1 0 10212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1644511149
transform -1 0 11684 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1644511149
transform -1 0 10028 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1644511149
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1644511149
transform -1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1644511149
transform -1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1644511149
transform -1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1644511149
transform -1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1644511149
transform -1 0 8096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1644511149
transform -1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1644511149
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1644511149
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1644511149
transform -1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1644511149
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1644511149
transform -1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1644511149
transform -1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1644511149
transform -1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1644511149
transform -1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1644511149
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1644511149
transform -1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1644511149
transform -1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1644511149
transform -1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1644511149
transform -1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1644511149
transform -1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1644511149
transform -1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1644511149
transform -1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1644511149
transform -1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1644511149
transform -1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1644511149
transform -1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1644511149
transform -1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1644511149
transform -1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1644511149
transform -1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1644511149
transform -1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1644511149
transform -1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input146_A
timestamp 1644511149
transform -1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input147_A
timestamp 1644511149
transform -1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input148_A
timestamp 1644511149
transform -1 0 37536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input149_A
timestamp 1644511149
transform -1 0 37536 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input150_A
timestamp 1644511149
transform -1 0 37536 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input151_A
timestamp 1644511149
transform -1 0 37536 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input152_A
timestamp 1644511149
transform -1 0 37444 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input153_A
timestamp 1644511149
transform -1 0 38180 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input154_A
timestamp 1644511149
transform -1 0 37536 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input155_A
timestamp 1644511149
transform -1 0 36800 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input156_A
timestamp 1644511149
transform -1 0 36800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input157_A
timestamp 1644511149
transform -1 0 36248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input158_A
timestamp 1644511149
transform -1 0 37444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input159_A
timestamp 1644511149
transform -1 0 38180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input160_A
timestamp 1644511149
transform -1 0 34868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input161_A
timestamp 1644511149
transform -1 0 37536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input162_A
timestamp 1644511149
transform -1 0 36892 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input163_A
timestamp 1644511149
transform -1 0 37536 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1644511149
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1644511149
transform -1 0 27048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output185_A
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output198_A
timestamp 1644511149
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output199_A
timestamp 1644511149
transform 1 0 16100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output204_A
timestamp 1644511149
transform -1 0 13432 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output209_A
timestamp 1644511149
transform -1 0 18768 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1644511149
transform 1 0 19872 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output223_A
timestamp 1644511149
transform 1 0 30820 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output224_A
timestamp 1644511149
transform 1 0 3036 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output225_A
timestamp 1644511149
transform 1 0 31924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1644511149
transform 1 0 32936 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1644511149
transform 1 0 34040 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output228_A
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output229_A
timestamp 1644511149
transform 1 0 35236 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1644511149
transform -1 0 36248 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1644511149
transform -1 0 34868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1644511149
transform -1 0 36892 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output233_A
timestamp 1644511149
transform -1 0 4508 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output242_A
timestamp 1644511149
transform -1 0 12972 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output243_A
timestamp 1644511149
transform 1 0 13892 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output244_A
timestamp 1644511149
transform 1 0 14536 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output245_A
timestamp 1644511149
transform 1 0 15916 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output246_A
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output247_A
timestamp 1644511149
transform -1 0 18216 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output248_A
timestamp 1644511149
transform 1 0 20424 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output249_A
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output252_A
timestamp 1644511149
transform 1 0 21896 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output253_A
timestamp 1644511149
transform 1 0 22816 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output254_A
timestamp 1644511149
transform -1 0 25024 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output255_A
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output256_A
timestamp 1644511149
transform -1 0 27140 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output261_A
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output262_A
timestamp 1644511149
transform -1 0 3772 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output263_A
timestamp 1644511149
transform -1 0 33856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output264_A
timestamp 1644511149
transform 1 0 33856 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output265_A
timestamp 1644511149
transform -1 0 34868 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output266_A
timestamp 1644511149
transform 1 0 35236 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output267_A
timestamp 1644511149
transform 1 0 35236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output268_A
timestamp 1644511149
transform 1 0 37444 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output270_A
timestamp 1644511149
transform -1 0 36340 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output271_A
timestamp 1644511149
transform -1 0 5060 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output272_A
timestamp 1644511149
transform -1 0 5612 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output273_A
timestamp 1644511149
transform -1 0 7452 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output274_A
timestamp 1644511149
transform -1 0 8004 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output275_A
timestamp 1644511149
transform -1 0 9292 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output276_A
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output277_A
timestamp 1644511149
transform -1 0 12236 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1644511149
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1644511149
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1644511149
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1644511149
transform 1 0 15640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1644511149
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1644511149
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_263
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_271
timestamp 1644511149
transform 1 0 26036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_348
timestamp 1644511149
transform 1 0 33120 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_42
timestamp 1644511149
transform 1 0 4968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_48
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1644511149
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1644511149
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 1644511149
transform 1 0 15088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1644511149
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_173
timestamp 1644511149
transform 1 0 17020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1644511149
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_207
timestamp 1644511149
transform 1 0 20148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_252
timestamp 1644511149
transform 1 0 24288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1644511149
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_313
timestamp 1644511149
transform 1 0 29900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_319
timestamp 1644511149
transform 1 0 30452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1644511149
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_351
timestamp 1644511149
transform 1 0 33396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_359
timestamp 1644511149
transform 1 0 34132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1644511149
transform 1 0 34684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1644511149
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1644511149
transform 1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_115
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_150
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1644511149
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_267
timestamp 1644511149
transform 1 0 25668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1644511149
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1644511149
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1644511149
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_324
timestamp 1644511149
transform 1 0 30912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1644511149
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_340
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_348
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_373
timestamp 1644511149
transform 1 0 35420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_385
timestamp 1644511149
transform 1 0 36524 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_61
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1644511149
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1644511149
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1644511149
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_203
timestamp 1644511149
transform 1 0 19780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_236
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_241
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_245
timestamp 1644511149
transform 1 0 23644 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_250
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_284
timestamp 1644511149
transform 1 0 27232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_291
timestamp 1644511149
transform 1 0 27876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1644511149
transform 1 0 28980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_313
timestamp 1644511149
transform 1 0 29900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_321
timestamp 1644511149
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_341
timestamp 1644511149
transform 1 0 32476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_348
timestamp 1644511149
transform 1 0 33120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_356
timestamp 1644511149
transform 1 0 33856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_375
timestamp 1644511149
transform 1 0 35604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_397
timestamp 1644511149
transform 1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 1644511149
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_37
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_45
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1644511149
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_68
timestamp 1644511149
transform 1 0 7360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1644511149
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_100
timestamp 1644511149
transform 1 0 10304 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_108
timestamp 1644511149
transform 1 0 11040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1644511149
transform 1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1644511149
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_123
timestamp 1644511149
transform 1 0 12420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1644511149
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_144
timestamp 1644511149
transform 1 0 14352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1644511149
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1644511149
transform 1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_164
timestamp 1644511149
transform 1 0 16192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 1644511149
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1644511149
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1644511149
transform 1 0 21160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_225
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_238
timestamp 1644511149
transform 1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1644511149
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_264
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1644511149
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1644511149
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_311
timestamp 1644511149
transform 1 0 29716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_317
timestamp 1644511149
transform 1 0 30268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_329
timestamp 1644511149
transform 1 0 31372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_341
timestamp 1644511149
transform 1 0 32476 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_353
timestamp 1644511149
transform 1 0 33580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_373
timestamp 1644511149
transform 1 0 35420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_379
timestamp 1644511149
transform 1 0 35972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_384
timestamp 1644511149
transform 1 0 36432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1644511149
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_5
timestamp 1644511149
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1644511149
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_59
timestamp 1644511149
transform 1 0 6532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1644511149
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_68
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_76
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1644511149
transform 1 0 8648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1644511149
transform 1 0 10304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1644511149
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1644511149
transform 1 0 12420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 1644511149
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1644511149
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_141
timestamp 1644511149
transform 1 0 14076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_147
timestamp 1644511149
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_150
timestamp 1644511149
transform 1 0 14904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1644511149
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_171
timestamp 1644511149
transform 1 0 16836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1644511149
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_192
timestamp 1644511149
transform 1 0 18768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_201
timestamp 1644511149
transform 1 0 19596 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_211
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_215
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1644511149
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_227
timestamp 1644511149
transform 1 0 21988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_239
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_247
timestamp 1644511149
transform 1 0 23828 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_253
timestamp 1644511149
transform 1 0 24380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_269
timestamp 1644511149
transform 1 0 25852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1644511149
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_285
timestamp 1644511149
transform 1 0 27324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_288
timestamp 1644511149
transform 1 0 27600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_294
timestamp 1644511149
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1644511149
transform 1 0 28520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1644511149
transform 1 0 28796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_308
timestamp 1644511149
transform 1 0 29440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1644511149
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_321
timestamp 1644511149
transform 1 0 30636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1644511149
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_340
timestamp 1644511149
transform 1 0 32384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_346
timestamp 1644511149
transform 1 0 32936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_350
timestamp 1644511149
transform 1 0 33304 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_359
timestamp 1644511149
transform 1 0 34132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_369
timestamp 1644511149
transform 1 0 35052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_377
timestamp 1644511149
transform 1 0 35788 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_383
timestamp 1644511149
transform 1 0 36340 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1644511149
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_5
timestamp 1644511149
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1644511149
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1644511149
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1644511149
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1644511149
transform 1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_62
timestamp 1644511149
transform 1 0 6808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_73
timestamp 1644511149
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1644511149
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_91 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1644511149
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1644511149
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_149
timestamp 1644511149
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1644511149
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_211
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_220
timestamp 1644511149
transform 1 0 21344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_226
timestamp 1644511149
transform 1 0 21896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1644511149
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_256
timestamp 1644511149
transform 1 0 24656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_260
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_263
timestamp 1644511149
transform 1 0 25300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1644511149
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1644511149
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_294
timestamp 1644511149
transform 1 0 28152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_317
timestamp 1644511149
transform 1 0 30268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_329
timestamp 1644511149
transform 1 0 31372 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_337
timestamp 1644511149
transform 1 0 32108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_343
timestamp 1644511149
transform 1 0 32660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_346
timestamp 1644511149
transform 1 0 32936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1644511149
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1644511149
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_368
timestamp 1644511149
transform 1 0 34960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_372
timestamp 1644511149
transform 1 0 35328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_376
timestamp 1644511149
transform 1 0 35696 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_382
timestamp 1644511149
transform 1 0 36248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_387
timestamp 1644511149
transform 1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1644511149
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_5
timestamp 1644511149
transform 1 0 1564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_17
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1644511149
transform 1 0 3220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1644511149
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1644511149
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1644511149
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1644511149
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1644511149
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_180
timestamp 1644511149
transform 1 0 17664 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_192
timestamp 1644511149
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_204
timestamp 1644511149
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1644511149
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_311
timestamp 1644511149
transform 1 0 29716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1644511149
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_326
timestamp 1644511149
transform 1 0 31096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1644511149
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_339
timestamp 1644511149
transform 1 0 32292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_347
timestamp 1644511149
transform 1 0 33028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_355
timestamp 1644511149
transform 1 0 33764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_367
timestamp 1644511149
transform 1 0 34868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_374
timestamp 1644511149
transform 1 0 35512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_381
timestamp 1644511149
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1644511149
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_401
timestamp 1644511149
transform 1 0 37996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_46
timestamp 1644511149
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1644511149
transform 1 0 6440 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1644511149
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_67
timestamp 1644511149
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_151
timestamp 1644511149
transform 1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 1644511149
transform 1 0 16192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_174
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1644511149
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1644511149
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1644511149
transform 1 0 19596 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1644511149
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_214
timestamp 1644511149
transform 1 0 20792 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_217
timestamp 1644511149
transform 1 0 21068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_229
timestamp 1644511149
transform 1 0 22172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_241
timestamp 1644511149
transform 1 0 23276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1644511149
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_261
timestamp 1644511149
transform 1 0 25116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_273
timestamp 1644511149
transform 1 0 26220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_285
timestamp 1644511149
transform 1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_291
timestamp 1644511149
transform 1 0 27876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_297
timestamp 1644511149
transform 1 0 28428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1644511149
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_314
timestamp 1644511149
transform 1 0 29992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_322
timestamp 1644511149
transform 1 0 30728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_328
timestamp 1644511149
transform 1 0 31280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_338
timestamp 1644511149
transform 1 0 32200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_344
timestamp 1644511149
transform 1 0 32752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_350
timestamp 1644511149
transform 1 0 33304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_356
timestamp 1644511149
transform 1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_367
timestamp 1644511149
transform 1 0 34868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_379
timestamp 1644511149
transform 1 0 35972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_382
timestamp 1644511149
transform 1 0 36248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_388
timestamp 1644511149
transform 1 0 36800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1644511149
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1644511149
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1644511149
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_92
timestamp 1644511149
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1644511149
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_116
timestamp 1644511149
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_128
timestamp 1644511149
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_140
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_158
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_284
timestamp 1644511149
transform 1 0 27232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_290
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1644511149
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_301
timestamp 1644511149
transform 1 0 28796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_313
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_325
timestamp 1644511149
transform 1 0 31004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1644511149
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1644511149
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_365
timestamp 1644511149
transform 1 0 34684 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_376
timestamp 1644511149
transform 1 0 35696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_382
timestamp 1644511149
transform 1 0 36248 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1644511149
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_401
timestamp 1644511149
transform 1 0 37996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1644511149
transform 1 0 11868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_129
timestamp 1644511149
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1644511149
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_211
timestamp 1644511149
transform 1 0 20516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_223
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_235
timestamp 1644511149
transform 1 0 22724 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_273
timestamp 1644511149
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_285
timestamp 1644511149
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_297
timestamp 1644511149
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1644511149
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_317
timestamp 1644511149
transform 1 0 30268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1644511149
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_342
timestamp 1644511149
transform 1 0 32568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_354
timestamp 1644511149
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1644511149
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_370
timestamp 1644511149
transform 1 0 35144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_376
timestamp 1644511149
transform 1 0 35696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_386
timestamp 1644511149
transform 1 0 36616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_394
timestamp 1644511149
transform 1 0 37352 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1644511149
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_22
timestamp 1644511149
transform 1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_35
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1644511149
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1644511149
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1644511149
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1644511149
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1644511149
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_97
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1644511149
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_119
timestamp 1644511149
transform 1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp 1644511149
transform 1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1644511149
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1644511149
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp 1644511149
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1644511149
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_254
timestamp 1644511149
transform 1 0 24472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_260
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_266
timestamp 1644511149
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1644511149
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_345
timestamp 1644511149
transform 1 0 32844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1644511149
transform 1 0 33672 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_366
timestamp 1644511149
transform 1 0 34776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_374
timestamp 1644511149
transform 1 0 35512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_377
timestamp 1644511149
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_383
timestamp 1644511149
transform 1 0 36340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_397
timestamp 1644511149
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1644511149
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_31
timestamp 1644511149
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_39
timestamp 1644511149
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1644511149
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1644511149
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_103
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1644511149
transform 1 0 11684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_127
timestamp 1644511149
transform 1 0 12788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1644511149
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1644511149
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_261
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_272
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_278
timestamp 1644511149
transform 1 0 26680 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_290
timestamp 1644511149
transform 1 0 27784 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1644511149
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_374
timestamp 1644511149
transform 1 0 35512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_381
timestamp 1644511149
transform 1 0 36156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_387
timestamp 1644511149
transform 1 0 36708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_393
timestamp 1644511149
transform 1 0 37260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_396
timestamp 1644511149
transform 1 0 37536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1644511149
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1644511149
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_146
timestamp 1644511149
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1644511149
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1644511149
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_177
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_201
timestamp 1644511149
transform 1 0 19596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1644511149
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1644511149
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_301
timestamp 1644511149
transform 1 0 28796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_306
timestamp 1644511149
transform 1 0 29256 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1644511149
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_49
timestamp 1644511149
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1644511149
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1644511149
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_157
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_175
timestamp 1644511149
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1644511149
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1644511149
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1644511149
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1644511149
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1644511149
transform 1 0 13524 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1644511149
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1644511149
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_179
timestamp 1644511149
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_191
timestamp 1644511149
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1644511149
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_289
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_292
timestamp 1644511149
transform 1 0 27968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_304
timestamp 1644511149
transform 1 0 29072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_316
timestamp 1644511149
transform 1 0 30176 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1644511149
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_381
timestamp 1644511149
transform 1 0 36156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1644511149
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_397
timestamp 1644511149
transform 1 0 37628 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1644511149
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1644511149
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1644511149
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_185
timestamp 1644511149
transform 1 0 18124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1644511149
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1644511149
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1644511149
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_283
timestamp 1644511149
transform 1 0 27140 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1644511149
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1644511149
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1644511149
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_29
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_41
timestamp 1644511149
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1644511149
transform 1 0 10028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1644511149
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_131
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_143
timestamp 1644511149
transform 1 0 14260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_155
timestamp 1644511149
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1644511149
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_202
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1644511149
transform 1 0 24748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1644511149
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_289
timestamp 1644511149
transform 1 0 27692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_299
timestamp 1644511149
transform 1 0 28612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_311
timestamp 1644511149
transform 1 0 29716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_315
timestamp 1644511149
transform 1 0 30084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_322
timestamp 1644511149
transform 1 0 30728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1644511149
transform 1 0 4508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_49
timestamp 1644511149
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_61
timestamp 1644511149
transform 1 0 6716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1644511149
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1644511149
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_100
timestamp 1644511149
transform 1 0 10304 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_112
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_124
timestamp 1644511149
transform 1 0 12512 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1644511149
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_216
timestamp 1644511149
transform 1 0 20976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_228
timestamp 1644511149
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_240
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_293
timestamp 1644511149
transform 1 0 28060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1644511149
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_331
timestamp 1644511149
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_343
timestamp 1644511149
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1644511149
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1644511149
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_85
timestamp 1644511149
transform 1 0 8924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_97
timestamp 1644511149
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1644511149
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_133
timestamp 1644511149
transform 1 0 13340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_145
timestamp 1644511149
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1644511149
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1644511149
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_204
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1644511149
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_247
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_259
timestamp 1644511149
transform 1 0 24932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1644511149
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_347
timestamp 1644511149
transform 1 0 33028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_354
timestamp 1644511149
transform 1 0 33672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_360
timestamp 1644511149
transform 1 0 34224 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_372
timestamp 1644511149
transform 1 0 35328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1644511149
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_399
timestamp 1644511149
transform 1 0 37812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1644511149
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_147
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_159
timestamp 1644511149
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_183
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_232
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_255
timestamp 1644511149
transform 1 0 24564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_267
timestamp 1644511149
transform 1 0 25668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_279
timestamp 1644511149
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_397
timestamp 1644511149
transform 1 0 37628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1644511149
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1644511149
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1644511149
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_177
timestamp 1644511149
transform 1 0 17388 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1644511149
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_255
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_263
timestamp 1644511149
transform 1 0 25300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1644511149
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_325
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_401
timestamp 1644511149
transform 1 0 37996 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1644511149
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_145
timestamp 1644511149
transform 1 0 14444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1644511149
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_229
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1644511149
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_255
timestamp 1644511149
transform 1 0 24564 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_267
timestamp 1644511149
transform 1 0 25668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_279
timestamp 1644511149
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_291
timestamp 1644511149
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1644511149
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_311
timestamp 1644511149
transform 1 0 29716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_323
timestamp 1644511149
transform 1 0 30820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_335
timestamp 1644511149
transform 1 0 31924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_347
timestamp 1644511149
transform 1 0 33028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1644511149
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_385
timestamp 1644511149
transform 1 0 36524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_72
timestamp 1644511149
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_84
timestamp 1644511149
transform 1 0 8832 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_96
timestamp 1644511149
transform 1 0 9936 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_177
timestamp 1644511149
transform 1 0 17388 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1644511149
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_239
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_242
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_248
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_260
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1644511149
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_291
timestamp 1644511149
transform 1 0 27876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_301
timestamp 1644511149
transform 1 0 28796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_311
timestamp 1644511149
transform 1 0 29716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_323
timestamp 1644511149
transform 1 0 30820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1644511149
transform 1 0 36064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_397
timestamp 1644511149
transform 1 0 37628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1644511149
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_35
timestamp 1644511149
transform 1 0 4324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_47
timestamp 1644511149
transform 1 0 5428 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_59
timestamp 1644511149
transform 1 0 6532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_71
timestamp 1644511149
transform 1 0 7636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1644511149
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1644511149
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_124
timestamp 1644511149
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1644511149
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1644511149
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1644511149
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_290
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1644511149
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_313
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_322
timestamp 1644511149
transform 1 0 30728 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_336
timestamp 1644511149
transform 1 0 32016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_342
timestamp 1644511149
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1644511149
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1644511149
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_368
timestamp 1644511149
transform 1 0 34960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_374
timestamp 1644511149
transform 1 0 35512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_382
timestamp 1644511149
transform 1 0 36248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_386
timestamp 1644511149
transform 1 0 36616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1644511149
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_398
timestamp 1644511149
transform 1 0 37720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1644511149
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_195
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_207
timestamp 1644511149
transform 1 0 20148 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_323
timestamp 1644511149
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_353
timestamp 1644511149
transform 1 0 33580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_366
timestamp 1644511149
transform 1 0 34776 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_378
timestamp 1644511149
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1644511149
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_401
timestamp 1644511149
transform 1 0 37996 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1644511149
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_67
timestamp 1644511149
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1644511149
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1644511149
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1644511149
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_183
timestamp 1644511149
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1644511149
transform 1 0 32292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1644511149
transform 1 0 33396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_397
timestamp 1644511149
transform 1 0 37628 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1644511149
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_65
timestamp 1644511149
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1644511149
transform 1 0 8004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_128
timestamp 1644511149
transform 1 0 12880 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_134
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_146
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_360
timestamp 1644511149
transform 1 0 34224 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_372
timestamp 1644511149
transform 1 0 35328 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 1644511149
transform 1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_34
timestamp 1644511149
transform 1 0 4232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_46
timestamp 1644511149
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_58
timestamp 1644511149
transform 1 0 6440 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_70
timestamp 1644511149
transform 1 0 7544 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_89
timestamp 1644511149
transform 1 0 9292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_95
timestamp 1644511149
transform 1 0 9844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_107
timestamp 1644511149
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_119
timestamp 1644511149
transform 1 0 12052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1644511149
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_255
timestamp 1644511149
transform 1 0 24564 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_267
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_279
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_291
timestamp 1644511149
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1644511149
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_397
timestamp 1644511149
transform 1 0 37628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_177
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_183
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_195
timestamp 1644511149
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_207
timestamp 1644511149
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1644511149
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_206
timestamp 1644511149
transform 1 0 20056 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_230
timestamp 1644511149
transform 1 0 22264 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_269
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_367
timestamp 1644511149
transform 1 0 34868 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_379
timestamp 1644511149
transform 1 0 35972 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_391
timestamp 1644511149
transform 1 0 37076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1644511149
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_140
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_152
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_312
timestamp 1644511149
transform 1 0 29808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_353
timestamp 1644511149
transform 1 0 33580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_363
timestamp 1644511149
transform 1 0 34500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_398
timestamp 1644511149
transform 1 0 37720 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1644511149
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_37
timestamp 1644511149
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_49
timestamp 1644511149
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1644511149
transform 1 0 6716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_69
timestamp 1644511149
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1644511149
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_100
timestamp 1644511149
transform 1 0 10304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_112
timestamp 1644511149
transform 1 0 11408 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1644511149
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_229
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_242
timestamp 1644511149
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_285
timestamp 1644511149
transform 1 0 27324 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1644511149
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_319
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_326
timestamp 1644511149
transform 1 0 31096 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_332
timestamp 1644511149
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_344
timestamp 1644511149
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1644511149
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_66
timestamp 1644511149
transform 1 0 7176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_78
timestamp 1644511149
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_90
timestamp 1644511149
transform 1 0 9384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1644511149
transform 1 0 11684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1644511149
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_299
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_323
timestamp 1644511149
transform 1 0 30820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_396
timestamp 1644511149
transform 1 0 37536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1644511149
transform 1 0 38180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_63
timestamp 1644511149
transform 1 0 6900 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_69
timestamp 1644511149
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1644511149
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1644511149
transform 1 0 12420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1644511149
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_400
timestamp 1644511149
transform 1 0 37904 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1644511149
transform 1 0 38456 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1644511149
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_26
timestamp 1644511149
transform 1 0 3496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1644511149
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1644511149
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_246
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1644511149
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp 1644511149
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1644511149
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_60
timestamp 1644511149
transform 1 0 6624 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_72
timestamp 1644511149
transform 1 0 7728 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_219
timestamp 1644511149
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_231
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1644511149
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_316
timestamp 1644511149
transform 1 0 30176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_329
timestamp 1644511149
transform 1 0 31372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_341
timestamp 1644511149
transform 1 0 32476 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1644511149
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_393
timestamp 1644511149
transform 1 0 37260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_396
timestamp 1644511149
transform 1 0 37536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_230
timestamp 1644511149
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_345
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_358
timestamp 1644511149
transform 1 0 34040 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_366
timestamp 1644511149
transform 1 0 34776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_371
timestamp 1644511149
transform 1 0 35236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1644511149
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_401
timestamp 1644511149
transform 1 0 37996 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_173
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1644511149
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1644511149
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_215
timestamp 1644511149
transform 1 0 20884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_220
timestamp 1644511149
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1644511149
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_284
timestamp 1644511149
transform 1 0 27232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_290
timestamp 1644511149
transform 1 0 27784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1644511149
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_337
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_348
timestamp 1644511149
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_397
timestamp 1644511149
transform 1 0 37628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_192
timestamp 1644511149
transform 1 0 18768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_198
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1644511149
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_316
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_324
timestamp 1644511149
transform 1 0 30912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_339
timestamp 1644511149
transform 1 0 32292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_351
timestamp 1644511149
transform 1 0 33396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_363
timestamp 1644511149
transform 1 0 34500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_375
timestamp 1644511149
transform 1 0 35604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1644511149
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_402
timestamp 1644511149
transform 1 0 38088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1644511149
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_128
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_259
timestamp 1644511149
transform 1 0 24932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1644511149
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1644511149
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_329
timestamp 1644511149
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_341
timestamp 1644511149
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1644511149
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1644511149
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1644511149
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_73
timestamp 1644511149
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_77
timestamp 1644511149
transform 1 0 8188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_94
timestamp 1644511149
transform 1 0 9752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_102
timestamp 1644511149
transform 1 0 10488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_122
timestamp 1644511149
transform 1 0 12328 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_130
timestamp 1644511149
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_61
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1644511149
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1644511149
transform 1 0 9292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_129
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_157
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_169
timestamp 1644511149
transform 1 0 16652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1644511149
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1644511149
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_334
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_340
timestamp 1644511149
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_352
timestamp 1644511149
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_11
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1644511149
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_35
timestamp 1644511149
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1644511149
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_77
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_153
timestamp 1644511149
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1644511149
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_241
timestamp 1644511149
transform 1 0 23276 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_247
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_285
timestamp 1644511149
transform 1 0 27324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_309
timestamp 1644511149
transform 1 0 29532 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1644511149
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_399
timestamp 1644511149
transform 1 0 37812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_35
timestamp 1644511149
transform 1 0 4324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_47
timestamp 1644511149
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_59
timestamp 1644511149
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_71
timestamp 1644511149
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1644511149
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_357
timestamp 1644511149
transform 1 0 33948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_377
timestamp 1644511149
transform 1 0 35788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1644511149
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_35
timestamp 1644511149
transform 1 0 4324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_48
timestamp 1644511149
transform 1 0 5520 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1644511149
transform 1 0 6072 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1644511149
transform 1 0 7176 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1644511149
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_169
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_286
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_298
timestamp 1644511149
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1644511149
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_336
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_373
timestamp 1644511149
transform 1 0 35420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_397
timestamp 1644511149
transform 1 0 37628 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1644511149
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_269
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_299
timestamp 1644511149
transform 1 0 28612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_341
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_353
timestamp 1644511149
transform 1 0 33580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_365
timestamp 1644511149
transform 1 0 34684 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_377
timestamp 1644511149
transform 1 0 35788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1644511149
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_57
timestamp 1644511149
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_181
timestamp 1644511149
transform 1 0 17756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_278
timestamp 1644511149
transform 1 0 26680 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1644511149
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_317
timestamp 1644511149
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_324
timestamp 1644511149
transform 1 0 30912 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_336
timestamp 1644511149
transform 1 0 32016 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_348
timestamp 1644511149
transform 1 0 33120 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_98
timestamp 1644511149
transform 1 0 10120 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1644511149
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_117
timestamp 1644511149
transform 1 0 11868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1644511149
transform 1 0 12420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_135
timestamp 1644511149
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_147
timestamp 1644511149
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1644511149
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_239
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_245
timestamp 1644511149
transform 1 0 23644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_257
timestamp 1644511149
transform 1 0 24748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_269
timestamp 1644511149
transform 1 0 25852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1644511149
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_93
timestamp 1644511149
transform 1 0 9660 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_99
timestamp 1644511149
transform 1 0 10212 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_107
timestamp 1644511149
transform 1 0 10948 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_112
timestamp 1644511149
transform 1 0 11408 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_124
timestamp 1644511149
transform 1 0 12512 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_266
timestamp 1644511149
transform 1 0 25576 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_278
timestamp 1644511149
transform 1 0 26680 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_290
timestamp 1644511149
transform 1 0 27784 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1644511149
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_344
timestamp 1644511149
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_393
timestamp 1644511149
transform 1 0 37260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_396
timestamp 1644511149
transform 1 0 37536 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_13
timestamp 1644511149
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_25
timestamp 1644511149
transform 1 0 3404 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_33
timestamp 1644511149
transform 1 0 4140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_41
timestamp 1644511149
transform 1 0 4876 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1644511149
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_64
timestamp 1644511149
transform 1 0 6992 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_76
timestamp 1644511149
transform 1 0 8096 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_88
timestamp 1644511149
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_100
timestamp 1644511149
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_118
timestamp 1644511149
transform 1 0 11960 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_124
timestamp 1644511149
transform 1 0 12512 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_132
timestamp 1644511149
transform 1 0 13248 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_150
timestamp 1644511149
transform 1 0 14904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_154
timestamp 1644511149
transform 1 0 15272 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_158
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_179
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_185
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1644511149
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1644511149
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_236
timestamp 1644511149
transform 1 0 22816 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_248
timestamp 1644511149
transform 1 0 23920 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_260
timestamp 1644511149
transform 1 0 25024 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1644511149
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_345
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_357
timestamp 1644511149
transform 1 0 33948 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_369
timestamp 1644511149
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_381
timestamp 1644511149
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1644511149
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_31
timestamp 1644511149
transform 1 0 3956 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_39
timestamp 1644511149
transform 1 0 4692 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_43
timestamp 1644511149
transform 1 0 5060 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_49
timestamp 1644511149
transform 1 0 5612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_61
timestamp 1644511149
transform 1 0 6716 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_73
timestamp 1644511149
transform 1 0 7820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1644511149
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1644511149
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_255
timestamp 1644511149
transform 1 0 24564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_267
timestamp 1644511149
transform 1 0 25668 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_275
timestamp 1644511149
transform 1 0 26404 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_291
timestamp 1644511149
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1644511149
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_341
timestamp 1644511149
transform 1 0 32476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_348
timestamp 1644511149
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_369
timestamp 1644511149
transform 1 0 35052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1644511149
transform 1 0 35328 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1644511149
transform 1 0 36432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_396
timestamp 1644511149
transform 1 0 37536 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_404
timestamp 1644511149
transform 1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_368
timestamp 1644511149
transform 1 0 34960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_396
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1644511149
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_268
timestamp 1644511149
transform 1 0 25760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_285
timestamp 1644511149
transform 1 0 27324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_288
timestamp 1644511149
transform 1 0 27600 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_297
timestamp 1644511149
transform 1 0 28428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1644511149
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_64
timestamp 1644511149
transform 1 0 6992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1644511149
transform 1 0 7544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1644511149
transform 1 0 8648 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1644511149
transform 1 0 9752 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1644511149
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_133
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1644511149
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1644511149
transform 1 0 25392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_346
timestamp 1644511149
transform 1 0 32936 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_370
timestamp 1644511149
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1644511149
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1644511149
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_397
timestamp 1644511149
transform 1 0 37628 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1644511149
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_201
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_207
timestamp 1644511149
transform 1 0 20148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_219
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_231
timestamp 1644511149
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_293
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1644511149
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1644511149
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_383
timestamp 1644511149
transform 1 0 36340 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_97
timestamp 1644511149
transform 1 0 10028 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp 1644511149
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1644511149
transform 1 0 12420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_135
timestamp 1644511149
transform 1 0 13524 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_147
timestamp 1644511149
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1644511149
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_187
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_194
timestamp 1644511149
transform 1 0 18952 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_206
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1644511149
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_320
timestamp 1644511149
transform 1 0 30544 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_369
timestamp 1644511149
transform 1 0 35052 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_379
timestamp 1644511149
transform 1 0 35972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_382
timestamp 1644511149
transform 1 0 36248 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1644511149
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_395
timestamp 1644511149
transform 1 0 37444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1644511149
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_106
timestamp 1644511149
transform 1 0 10856 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_112
timestamp 1644511149
transform 1 0 11408 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_124
timestamp 1644511149
transform 1 0 12512 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_163
timestamp 1644511149
transform 1 0 16100 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_171
timestamp 1644511149
transform 1 0 16836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_175
timestamp 1644511149
transform 1 0 17204 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_183
timestamp 1644511149
transform 1 0 17940 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1644511149
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1644511149
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_241
timestamp 1644511149
transform 1 0 23276 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 1644511149
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_327
timestamp 1644511149
transform 1 0 31188 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_355
timestamp 1644511149
transform 1 0 33764 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_358
timestamp 1644511149
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_367
timestamp 1644511149
transform 1 0 34868 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_373
timestamp 1644511149
transform 1 0 35420 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_379
timestamp 1644511149
transform 1 0 35972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_386
timestamp 1644511149
transform 1 0 36616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_394
timestamp 1644511149
transform 1 0 37352 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_402
timestamp 1644511149
transform 1 0 38088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1644511149
transform 1 0 38456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_17
timestamp 1644511149
transform 1 0 2668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_23
timestamp 1644511149
transform 1 0 3220 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_29
timestamp 1644511149
transform 1 0 3772 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_35
timestamp 1644511149
transform 1 0 4324 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1644511149
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_59
timestamp 1644511149
transform 1 0 6532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_71
timestamp 1644511149
transform 1 0 7636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_83
timestamp 1644511149
transform 1 0 8740 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_89
timestamp 1644511149
transform 1 0 9292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_95
timestamp 1644511149
transform 1 0 9844 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_103
timestamp 1644511149
transform 1 0 10580 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_106
timestamp 1644511149
transform 1 0 10856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_115
timestamp 1644511149
transform 1 0 11684 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_121
timestamp 1644511149
transform 1 0 12236 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_129
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_141
timestamp 1644511149
transform 1 0 14076 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_145
timestamp 1644511149
transform 1 0 14444 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_148
timestamp 1644511149
transform 1 0 14720 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_154
timestamp 1644511149
transform 1 0 15272 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_160
timestamp 1644511149
transform 1 0 15824 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_173
timestamp 1644511149
transform 1 0 17020 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_177
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1644511149
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 1644511149
transform 1 0 19504 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_206
timestamp 1644511149
transform 1 0 20056 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_212
timestamp 1644511149
transform 1 0 20608 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_229
timestamp 1644511149
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_232
timestamp 1644511149
transform 1 0 22448 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_242
timestamp 1644511149
transform 1 0 23368 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_252
timestamp 1644511149
transform 1 0 24288 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_345
timestamp 1644511149
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_348
timestamp 1644511149
transform 1 0 33120 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_356
timestamp 1644511149
transform 1 0 33856 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_364
timestamp 1644511149
transform 1 0 34592 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1644511149
transform 1 0 34868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_380
timestamp 1644511149
transform 1 0 36064 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_395
timestamp 1644511149
transform 1 0 37444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1644511149
transform 1 0 38180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_13
timestamp 1644511149
transform 1 0 2300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1644511149
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_31
timestamp 1644511149
transform 1 0 3956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_37
timestamp 1644511149
transform 1 0 4508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_43
timestamp 1644511149
transform 1 0 5060 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_49
timestamp 1644511149
transform 1 0 5612 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_57
timestamp 1644511149
transform 1 0 6348 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_63
timestamp 1644511149
transform 1 0 6900 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_69
timestamp 1644511149
transform 1 0 7452 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_75
timestamp 1644511149
transform 1 0 8004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_87
timestamp 1644511149
transform 1 0 9108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_104
timestamp 1644511149
transform 1 0 10672 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_110
timestamp 1644511149
transform 1 0 11224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_116
timestamp 1644511149
transform 1 0 11776 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_122
timestamp 1644511149
transform 1 0 12328 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1644511149
transform 1 0 12880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_134
timestamp 1644511149
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_147
timestamp 1644511149
transform 1 0 14628 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_151
timestamp 1644511149
transform 1 0 14996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_155
timestamp 1644511149
transform 1 0 15364 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_162
timestamp 1644511149
transform 1 0 16008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_168
timestamp 1644511149
transform 1 0 16560 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1644511149
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_180
timestamp 1644511149
transform 1 0 17664 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_186
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_199
timestamp 1644511149
transform 1 0 19412 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_207
timestamp 1644511149
transform 1 0 20148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_213
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_219
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_235
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1644511149
transform 1 0 27600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_300
timestamp 1644511149
transform 1 0 28704 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_322
timestamp 1644511149
transform 1 0 30728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_331
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_337
timestamp 1644511149
transform 1 0 32108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_348
timestamp 1644511149
transform 1 0 33120 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_354
timestamp 1644511149
transform 1 0 33672 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_367
timestamp 1644511149
transform 1 0 34868 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_375
timestamp 1644511149
transform 1 0 35604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_395
timestamp 1644511149
transform 1 0 37444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_13
timestamp 1644511149
transform 1 0 2300 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_20
timestamp 1644511149
transform 1 0 2944 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_33
timestamp 1644511149
transform 1 0 4140 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_45
timestamp 1644511149
transform 1 0 5244 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_49
timestamp 1644511149
transform 1 0 5612 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1644511149
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_61
timestamp 1644511149
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_67
timestamp 1644511149
transform 1 0 7268 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_77
timestamp 1644511149
transform 1 0 8188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_84
timestamp 1644511149
transform 1 0 8832 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_92
timestamp 1644511149
transform 1 0 9568 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_97
timestamp 1644511149
transform 1 0 10028 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1644511149
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_116
timestamp 1644511149
transform 1 0 11776 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_120
timestamp 1644511149
transform 1 0 12144 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_124
timestamp 1644511149
transform 1 0 12512 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_130
timestamp 1644511149
transform 1 0 13064 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_136
timestamp 1644511149
transform 1 0 13616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_145
timestamp 1644511149
transform 1 0 14444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_152
timestamp 1644511149
transform 1 0 15088 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_156
timestamp 1644511149
transform 1 0 15456 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_172
timestamp 1644511149
transform 1 0 16928 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_179
timestamp 1644511149
transform 1 0 17572 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_185
timestamp 1644511149
transform 1 0 18124 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_196
timestamp 1644511149
transform 1 0 19136 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_203
timestamp 1644511149
transform 1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_209
timestamp 1644511149
transform 1 0 20332 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1644511149
transform 1 0 22632 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_242
timestamp 1644511149
transform 1 0 23368 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1644511149
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_254
timestamp 1644511149
transform 1 0 24472 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_266
timestamp 1644511149
transform 1 0 25576 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_272
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_283
timestamp 1644511149
transform 1 0 27140 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_297
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_303
timestamp 1644511149
transform 1 0 28980 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_314
timestamp 1644511149
transform 1 0 29992 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_322
timestamp 1644511149
transform 1 0 30728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_326
timestamp 1644511149
transform 1 0 31096 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_341
timestamp 1644511149
transform 1 0 32476 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_346
timestamp 1644511149
transform 1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_354
timestamp 1644511149
transform 1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1644511149
transform 1 0 34408 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_366
timestamp 1644511149
transform 1 0 34776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_371
timestamp 1644511149
transform 1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_379
timestamp 1644511149
transform 1 0 35972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_383
timestamp 1644511149
transform 1 0 36340 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1644511149
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_395
timestamp 1644511149
transform 1 0 37444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_35
timestamp 1644511149
transform 1 0 4324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_39
timestamp 1644511149
transform 1 0 4692 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_42
timestamp 1644511149
transform 1 0 4968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_49
timestamp 1644511149
transform 1 0 5612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_58
timestamp 1644511149
transform 1 0 6440 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_70
timestamp 1644511149
transform 1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_89
timestamp 1644511149
transform 1 0 9292 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_95
timestamp 1644511149
transform 1 0 9844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_100
timestamp 1644511149
transform 1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_108
timestamp 1644511149
transform 1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_116
timestamp 1644511149
transform 1 0 11776 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_122
timestamp 1644511149
transform 1 0 12328 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_127
timestamp 1644511149
transform 1 0 12788 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_145
timestamp 1644511149
transform 1 0 14444 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1644511149
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_159
timestamp 1644511149
transform 1 0 15732 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_164
timestamp 1644511149
transform 1 0 16192 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_173
timestamp 1644511149
transform 1 0 17020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_179
timestamp 1644511149
transform 1 0 17572 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_184
timestamp 1644511149
transform 1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1644511149
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_201
timestamp 1644511149
transform 1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_208
timestamp 1644511149
transform 1 0 20240 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_215
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1644511149
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1644511149
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_264
timestamp 1644511149
transform 1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_268
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_271
timestamp 1644511149
transform 1 0 26036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_278
timestamp 1644511149
transform 1 0 26680 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_285
timestamp 1644511149
transform 1 0 27324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_291
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1644511149
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_311
timestamp 1644511149
transform 1 0 29716 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_315
timestamp 1644511149
transform 1 0 30084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_320
timestamp 1644511149
transform 1 0 30544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_328
timestamp 1644511149
transform 1 0 31280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_336
timestamp 1644511149
transform 1 0 32016 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_344
timestamp 1644511149
transform 1 0 32752 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_354
timestamp 1644511149
transform 1 0 33672 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_369
timestamp 1644511149
transform 1 0 35052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_375
timestamp 1644511149
transform 1 0 35604 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_11
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_35
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_61
timestamp 1644511149
transform 1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_77
timestamp 1644511149
transform 1 0 8188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_85
timestamp 1644511149
transform 1 0 8924 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_103
timestamp 1644511149
transform 1 0 10580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_115
timestamp 1644511149
transform 1 0 11684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_123
timestamp 1644511149
transform 1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1644511149
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_139
timestamp 1644511149
transform 1 0 13892 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_147
timestamp 1644511149
transform 1 0 14628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_153
timestamp 1644511149
transform 1 0 15180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_157
timestamp 1644511149
transform 1 0 15548 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1644511149
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_177
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1644511149
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_211
timestamp 1644511149
transform 1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1644511149
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_253
timestamp 1644511149
transform 1 0 24380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_269
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_285
timestamp 1644511149
transform 1 0 27324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1644511149
transform 1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_324
timestamp 1644511149
transform 1 0 30912 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_341
timestamp 1644511149
transform 1 0 32476 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_347
timestamp 1644511149
transform 1 0 33028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_352
timestamp 1644511149
transform 1 0 33488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_364
timestamp 1644511149
transform 1 0 34592 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_370
timestamp 1644511149
transform 1 0 35144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_375
timestamp 1644511149
transform 1 0 35604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_387
timestamp 1644511149
transform 1 0 36708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1644511149
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1644511149
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_13
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1644511149
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_52
timestamp 1644511149
transform 1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_67
timestamp 1644511149
transform 1 0 7268 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_75
timestamp 1644511149
transform 1 0 8004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_95
timestamp 1644511149
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_103
timestamp 1644511149
transform 1 0 10580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1644511149
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_123
timestamp 1644511149
transform 1 0 12420 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_149
timestamp 1644511149
transform 1 0 14812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_157
timestamp 1644511149
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_163
timestamp 1644511149
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1644511149
transform 1 0 17940 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_190
timestamp 1644511149
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_201
timestamp 1644511149
transform 1 0 19596 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_211
timestamp 1644511149
transform 1 0 20516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 1644511149
transform 1 0 21252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1644511149
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_241
timestamp 1644511149
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1644511149
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_257
timestamp 1644511149
transform 1 0 24748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_263
timestamp 1644511149
transform 1 0 25300 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_268
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1644511149
transform 1 0 26496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_285
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1644511149
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1644511149
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_313
timestamp 1644511149
transform 1 0 29900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1644511149
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 1644511149
transform 1 0 34132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_369
timestamp 1644511149
transform 1 0 35052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1644511149
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1644511149
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_397
timestamp 1644511149
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _193_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _194_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _195_
timestamp 1644511149
transform 1 0 9200 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1644511149
transform -1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _197_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1644511149
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _199_
timestamp 1644511149
transform 1 0 12052 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1644511149
transform -1 0 12420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _201_
timestamp 1644511149
transform 1 0 14444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1644511149
transform -1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _203_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27876 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _204_
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _205_
timestamp 1644511149
transform -1 0 23828 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _206_
timestamp 1644511149
transform 1 0 25944 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _207_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _208_
timestamp 1644511149
transform 1 0 22356 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _209_
timestamp 1644511149
transform -1 0 23184 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _210_
timestamp 1644511149
transform -1 0 32016 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1644511149
transform -1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _212_
timestamp 1644511149
transform 1 0 20332 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1644511149
transform 1 0 19320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _214_
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1644511149
transform -1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _216_
timestamp 1644511149
transform 1 0 25668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _218_
timestamp 1644511149
transform -1 0 29900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _220_
timestamp 1644511149
transform -1 0 24472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1644511149
transform -1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _222_
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _223_
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _224_
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1644511149
transform -1 0 25944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _226_
timestamp 1644511149
transform 1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1644511149
transform -1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _228_
timestamp 1644511149
transform 1 0 6532 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1644511149
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _230_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _231_
timestamp 1644511149
transform -1 0 27692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1644511149
transform -1 0 28704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _233_
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1644511149
transform -1 0 29256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _235_
timestamp 1644511149
transform 1 0 27968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1644511149
transform -1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _237_
timestamp 1644511149
transform -1 0 32200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1644511149
transform -1 0 33120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _239_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1644511149
transform -1 0 33672 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _241_
timestamp 1644511149
transform 1 0 14260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1644511149
transform -1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _243_
timestamp 1644511149
transform 1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1644511149
transform -1 0 35696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _245_
timestamp 1644511149
transform 1 0 16652 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1644511149
transform -1 0 36156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _247_
timestamp 1644511149
transform 1 0 35604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _248_
timestamp 1644511149
transform 1 0 36984 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_4  _249_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1644511149
transform 1 0 2668 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _251_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 3312 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _253_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _254_
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1644511149
transform -1 0 3496 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1644511149
transform 1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _258_
timestamp 1644511149
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1644511149
transform 1 0 6164 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp 1644511149
transform 1 0 5888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _261_
timestamp 1644511149
transform 1 0 32200 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _263_
timestamp 1644511149
transform -1 0 30544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _265_
timestamp 1644511149
transform -1 0 31280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _266_
timestamp 1644511149
transform -1 0 31648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _267_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _268_
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _269_
timestamp 1644511149
transform -1 0 32752 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_4  _270_
timestamp 1644511149
transform -1 0 32844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1644511149
transform 1 0 12236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _272_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _273_
timestamp 1644511149
transform -1 0 33672 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _274_
timestamp 1644511149
transform -1 0 13248 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _275_
timestamp 1644511149
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _277_
timestamp 1644511149
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1644511149
transform -1 0 16560 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _279_
timestamp 1644511149
transform -1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _281_
timestamp 1644511149
transform -1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _283_
timestamp 1644511149
transform -1 0 36892 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _284_
timestamp 1644511149
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1644511149
transform -1 0 20240 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1644511149
transform -1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _288_
timestamp 1644511149
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _289_
timestamp 1644511149
transform 1 0 22172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _290_
timestamp 1644511149
transform -1 0 10764 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _291_
timestamp 1644511149
transform 1 0 23552 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _292_
timestamp 1644511149
transform -1 0 11684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _293_
timestamp 1644511149
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp 1644511149
transform -1 0 13156 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _295_
timestamp 1644511149
transform 1 0 24748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _296_
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1644511149
transform 1 0 27048 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1644511149
transform -1 0 27324 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1644511149
transform 1 0 28612 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _301_
timestamp 1644511149
transform 1 0 22816 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1644511149
transform -1 0 28244 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1644511149
transform 1 0 31280 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _305_
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _306_
timestamp 1644511149
transform 1 0 30452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1644511149
transform 1 0 33948 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _308_
timestamp 1644511149
transform -1 0 34224 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1644511149
transform -1 0 19780 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _310_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1644511149
transform -1 0 20976 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _312_
timestamp 1644511149
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1644511149
transform -1 0 22632 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1644511149
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1644511149
transform -1 0 23828 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _316_
timestamp 1644511149
transform -1 0 35788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_4  _317_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 2668 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _319_
timestamp 1644511149
transform -1 0 30728 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _320_
timestamp 1644511149
transform -1 0 26036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_4  _321_
timestamp 1644511149
transform -1 0 32568 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _323_
timestamp 1644511149
transform -1 0 18216 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform -1 0 19780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _325_
timestamp 1644511149
transform 1 0 23736 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1644511149
transform -1 0 27784 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _327_
timestamp 1644511149
transform -1 0 28796 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _328_
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _329_
timestamp 1644511149
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _330_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27324 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _331_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22264 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _332_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20240 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _333_
timestamp 1644511149
transform -1 0 12880 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _334_
timestamp 1644511149
transform -1 0 13156 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _335_
timestamp 1644511149
transform -1 0 7728 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _336_
timestamp 1644511149
transform -1 0 7176 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _337_
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _338_
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _339_
timestamp 1644511149
transform 1 0 19780 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1644511149
transform -1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _341_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32476 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _342_
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _343_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32016 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _344_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _345_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _346_
timestamp 1644511149
transform -1 0 32752 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _347_
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1644511149
transform -1 0 34960 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _349_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26128 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1644511149
transform 1 0 5612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _351_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3128 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _352_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _353_
timestamp 1644511149
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _354_
timestamp 1644511149
transform 1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _355_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1644511149
transform 1 0 5336 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _357_
timestamp 1644511149
transform -1 0 7912 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1644511149
transform -1 0 6716 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _359_
timestamp 1644511149
transform -1 0 29992 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _360_
timestamp 1644511149
transform 1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _361_
timestamp 1644511149
transform -1 0 30820 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _363_
timestamp 1644511149
transform -1 0 31648 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1644511149
transform 1 0 10396 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _365_
timestamp 1644511149
transform -1 0 33672 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _366_
timestamp 1644511149
transform -1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _367_
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _369_
timestamp 1644511149
transform -1 0 15640 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1644511149
transform 1 0 14168 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _371_
timestamp 1644511149
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _373_
timestamp 1644511149
transform -1 0 18032 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp 1644511149
transform 1 0 17296 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _375_
timestamp 1644511149
transform -1 0 37720 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _376_
timestamp 1644511149
transform 1 0 37260 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _377_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1644511149
transform -1 0 20884 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _379_
timestamp 1644511149
transform 1 0 10120 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1644511149
transform -1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _381_
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _382_
timestamp 1644511149
transform -1 0 13616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _383_
timestamp 1644511149
transform -1 0 13064 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1644511149
transform -1 0 15364 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _385_
timestamp 1644511149
transform -1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1644511149
transform -1 0 16008 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1644511149
transform -1 0 26496 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _389_
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _390_
timestamp 1644511149
transform -1 0 26680 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _391_
timestamp 1644511149
transform 1 0 27968 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1644511149
transform -1 0 29440 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _393_
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _394_
timestamp 1644511149
transform 1 0 31372 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _395_
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _396_
timestamp 1644511149
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _397_
timestamp 1644511149
transform 1 0 20516 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _398_
timestamp 1644511149
transform 1 0 33028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _399_
timestamp 1644511149
transform 1 0 25208 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _400_
timestamp 1644511149
transform 1 0 33948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _401_
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _402_
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _403_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34960 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _404_
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _405_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33948 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _406_
timestamp 1644511149
transform -1 0 30452 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _407_
timestamp 1644511149
transform 1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _408_
timestamp 1644511149
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _409_
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _410_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23552 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _411_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _412_
timestamp 1644511149
transform -1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _413_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _414_
timestamp 1644511149
transform -1 0 27324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _415_
timestamp 1644511149
transform -1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _416_
timestamp 1644511149
transform 1 0 25024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _417_
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _418_
timestamp 1644511149
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _419_
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _420_
timestamp 1644511149
transform -1 0 21252 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _421_
timestamp 1644511149
transform 1 0 20976 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _422_
timestamp 1644511149
transform -1 0 18124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _423_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _424_
timestamp 1644511149
transform -1 0 20056 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _425_
timestamp 1644511149
transform -1 0 17940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _426_
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _427_
timestamp 1644511149
transform -1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _428_
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _429_
timestamp 1644511149
transform -1 0 13432 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _430_
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _431_
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _432_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _433_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1644511149
transform -1 0 9752 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1644511149
transform 1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1644511149
transform -1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _437_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13064 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _438_
timestamp 1644511149
transform 1 0 8096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _439_
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _440_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _441_
timestamp 1644511149
transform -1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1644511149
transform -1 0 4232 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _443_
timestamp 1644511149
transform -1 0 3312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _444_
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _445_
timestamp 1644511149
transform -1 0 7268 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _446_
timestamp 1644511149
transform -1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _447_
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _448_
timestamp 1644511149
transform 1 0 7360 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _449_
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _450_
timestamp 1644511149
transform 1 0 6808 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _451_
timestamp 1644511149
transform 1 0 6348 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _452_
timestamp 1644511149
transform 1 0 6716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _453_
timestamp 1644511149
transform 1 0 4416 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _454_
timestamp 1644511149
transform 1 0 5244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _455_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _456_
timestamp 1644511149
transform -1 0 5428 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _457_
timestamp 1644511149
transform 1 0 4784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _458_
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _459_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _460_
timestamp 1644511149
transform -1 0 6992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _461_
timestamp 1644511149
transform 1 0 5244 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _462_
timestamp 1644511149
transform -1 0 11868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _463_
timestamp 1644511149
transform 1 0 10120 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _464_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _465_
timestamp 1644511149
transform -1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _466_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _467_
timestamp 1644511149
transform -1 0 17572 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _468_
timestamp 1644511149
transform -1 0 15640 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _469_
timestamp 1644511149
transform 1 0 14352 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _470_
timestamp 1644511149
transform -1 0 19596 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _471_
timestamp 1644511149
transform 1 0 18400 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _472_
timestamp 1644511149
transform -1 0 19412 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _473_
timestamp 1644511149
transform -1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _474_
timestamp 1644511149
transform -1 0 18492 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _475_
timestamp 1644511149
transform -1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _476_
timestamp 1644511149
transform -1 0 22816 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _477_
timestamp 1644511149
transform -1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _478_
timestamp 1644511149
transform -1 0 27416 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _479_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _480_
timestamp 1644511149
transform -1 0 31648 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _481_
timestamp 1644511149
transform -1 0 23828 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1644511149
transform 1 0 25760 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1644511149
transform 1 0 25760 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1644511149
transform 1 0 17296 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1644511149
transform 1 0 6900 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1644511149
transform -1 0 15548 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1644511149
transform 1 0 2024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1644511149
transform 1 0 2668 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1644511149
transform 1 0 6900 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1644511149
transform 1 0 4600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1644511149
transform 1 0 2300 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1644511149
transform 1 0 1840 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1644511149
transform 1 0 4416 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1644511149
transform 1 0 9384 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1644511149
transform 1 0 8648 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1644511149
transform 1 0 14076 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1644511149
transform -1 0 23736 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1644511149
transform 1 0 27140 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1644511149
transform 1 0 36156 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1644511149
transform 1 0 35972 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1644511149
transform -1 0 35788 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1644511149
transform -1 0 36800 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _510__280 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _511__281
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _512__282
timestamp 1644511149
transform 1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _513__283
timestamp 1644511149
transform 1 0 37904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514__284
timestamp 1644511149
transform 1 0 37904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515__285
timestamp 1644511149
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _516_
timestamp 1644511149
transform 1 0 2576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1644511149
transform -1 0 30084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _518_
timestamp 1644511149
transform -1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1644511149
transform -1 0 36800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _520_
timestamp 1644511149
transform -1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1644511149
transform -1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _522_
timestamp 1644511149
transform -1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _523_
timestamp 1644511149
transform -1 0 30268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _524_
timestamp 1644511149
transform -1 0 36524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _525_
timestamp 1644511149
transform -1 0 37996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _526_
timestamp 1644511149
transform -1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _527_
timestamp 1644511149
transform -1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _528_
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _529_
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _530_
timestamp 1644511149
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _531_
timestamp 1644511149
transform 1 0 36984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _532_
timestamp 1644511149
transform 1 0 37628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _533_
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _534_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _535_
timestamp 1644511149
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _536_
timestamp 1644511149
transform 1 0 36432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform -1 0 10488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform -1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform -1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform -1 0 28612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform -1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 33028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 33856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform -1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1644511149
transform -1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform -1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 37444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform -1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform -1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform -1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1644511149
transform -1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 30544 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1644511149
transform 1 0 32200 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 33304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform -1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform -1 0 35420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform -1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 35880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform -1 0 38180 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform -1 0 35512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 27600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform -1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform -1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1644511149
transform -1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform -1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1644511149
transform 1 0 29992 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform -1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1644511149
transform 1 0 32476 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform -1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform -1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform -1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform -1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1644511149
transform 1 0 9476 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform -1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform -1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform -1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 24472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1644511149
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1644511149
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 11868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 12788 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1644511149
transform 1 0 12788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1644511149
transform -1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1644511149
transform 1 0 17020 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input85
timestamp 1644511149
transform 1 0 18032 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1644511149
transform 1 0 20148 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input88
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1644511149
transform -1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1644511149
transform -1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input93
timestamp 1644511149
transform 1 0 25392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1644511149
transform -1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1644511149
transform 1 0 31372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1644511149
transform -1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1644511149
transform 1 0 2668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1644511149
transform -1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1644511149
transform -1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1644511149
transform -1 0 35052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1644511149
transform -1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1644511149
transform -1 0 36524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1644511149
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1644511149
transform -1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1644511149
transform -1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1644511149
transform -1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input111
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 1644511149
transform 1 0 7636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input113
timestamp 1644511149
transform 1 0 9292 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1644511149
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input115
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1644511149
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input123
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input124
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1644511149
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input129
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1644511149
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1644511149
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1644511149
transform -1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1644511149
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1644511149
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input136
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input137
timestamp 1644511149
transform 1 0 8648 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1644511149
transform -1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1644511149
transform -1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1644511149
transform -1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1644511149
transform -1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1644511149
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1644511149
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1644511149
transform -1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input147
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1644511149
transform 1 0 37904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1644511149
transform 1 0 37904 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1644511149
transform 1 0 37904 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1644511149
transform -1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input153
timestamp 1644511149
transform -1 0 38180 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1644511149
transform 1 0 36340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1644511149
transform -1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input157
timestamp 1644511149
transform -1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input158
timestamp 1644511149
transform -1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1644511149
transform -1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1644511149
transform 1 0 35880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1644511149
transform 1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input162
timestamp 1644511149
transform 1 0 37260 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1644511149
transform 1 0 37904 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 32752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 35236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 36064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 36432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 37076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform -1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform -1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform 1 0 31004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform 1 0 32016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform -1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform -1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform -1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform -1 0 21068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform -1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform -1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform -1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform -1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1644511149
transform -1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1644511149
transform -1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1644511149
transform -1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1644511149
transform -1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1644511149
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1644511149
transform 1 0 10672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1644511149
transform -1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1644511149
transform -1 0 13892 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1644511149
transform 1 0 14260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1644511149
transform -1 0 16008 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1644511149
transform -1 0 16192 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1644511149
transform -1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1644511149
transform -1 0 18860 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1644511149
transform -1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1644511149
transform -1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1644511149
transform 1 0 24748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1644511149
transform 1 0 27876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1644511149
transform 1 0 3220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1644511149
transform 1 0 33120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1644511149
transform 1 0 34224 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1644511149
transform 1 0 35236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1644511149
transform 1 0 36340 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1644511149
transform 1 0 36432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1644511149
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1644511149
transform 1 0 37812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1644511149
transform -1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1644511149
transform -1 0 5060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1644511149
transform 1 0 7084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1644511149
transform -1 0 8188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1644511149
transform -1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1644511149
transform -1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1644511149
transform -1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1644511149
transform -1 0 11776 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1644511149
transform -1 0 12788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1644511149
transform 1 0 14996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1644511149
transform -1 0 15916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1644511149
transform -1 0 17020 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1644511149
transform -1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1644511149
transform -1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1644511149
transform -1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1644511149
transform -1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1644511149
transform -1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1644511149
transform 1 0 23000 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1644511149
transform -1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1644511149
transform 1 0 27692 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1644511149
transform -1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1644511149
transform -1 0 30728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1644511149
transform 1 0 31648 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1644511149
transform -1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1644511149
transform -1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1644511149
transform 1 0 34040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1644511149
transform 1 0 35604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1644511149
transform -1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1644511149
transform 1 0 37720 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1644511149
transform 1 0 37812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1644511149
transform 1 0 36984 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1644511149
transform -1 0 4324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1644511149
transform 1 0 5428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1644511149
transform -1 0 6440 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1644511149
transform -1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1644511149
transform -1 0 9292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1644511149
transform -1 0 10028 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1644511149
transform -1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1644511149
transform -1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1644511149
transform -1 0 35604 0 1 34816
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 9936 800 10056 6 clk
port 0 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 gpio0_input[0]
port 1 nsew signal tristate
rlabel metal2 s 32678 0 32734 800 6 gpio0_input[10]
port 2 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 gpio0_input[11]
port 3 nsew signal tristate
rlabel metal2 s 34334 0 34390 800 6 gpio0_input[12]
port 4 nsew signal tristate
rlabel metal2 s 35162 0 35218 800 6 gpio0_input[13]
port 5 nsew signal tristate
rlabel metal2 s 35990 0 36046 800 6 gpio0_input[14]
port 6 nsew signal tristate
rlabel metal2 s 36818 0 36874 800 6 gpio0_input[15]
port 7 nsew signal tristate
rlabel metal2 s 37646 0 37702 800 6 gpio0_input[16]
port 8 nsew signal tristate
rlabel metal2 s 38474 0 38530 800 6 gpio0_input[17]
port 9 nsew signal tristate
rlabel metal2 s 39302 0 39358 800 6 gpio0_input[18]
port 10 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 gpio0_input[1]
port 11 nsew signal tristate
rlabel metal2 s 26146 0 26202 800 6 gpio0_input[2]
port 12 nsew signal tristate
rlabel metal2 s 26882 0 26938 800 6 gpio0_input[3]
port 13 nsew signal tristate
rlabel metal2 s 27710 0 27766 800 6 gpio0_input[4]
port 14 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 gpio0_input[5]
port 15 nsew signal tristate
rlabel metal2 s 29366 0 29422 800 6 gpio0_input[6]
port 16 nsew signal tristate
rlabel metal2 s 30194 0 30250 800 6 gpio0_input[7]
port 17 nsew signal tristate
rlabel metal2 s 31022 0 31078 800 6 gpio0_input[8]
port 18 nsew signal tristate
rlabel metal2 s 31850 0 31906 800 6 gpio0_input[9]
port 19 nsew signal tristate
rlabel metal2 s 24766 0 24822 800 6 gpio0_oe[0]
port 20 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 gpio0_oe[10]
port 21 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 gpio0_oe[11]
port 22 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 gpio0_oe[12]
port 23 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 gpio0_oe[13]
port 24 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 gpio0_oe[14]
port 25 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 gpio0_oe[15]
port 26 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 gpio0_oe[16]
port 27 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 gpio0_oe[17]
port 28 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 gpio0_oe[18]
port 29 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 gpio0_oe[1]
port 30 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 gpio0_oe[2]
port 31 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 gpio0_oe[3]
port 32 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 gpio0_oe[4]
port 33 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 gpio0_oe[5]
port 34 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 gpio0_oe[6]
port 35 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 gpio0_oe[7]
port 36 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 gpio0_oe[8]
port 37 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 gpio0_oe[9]
port 38 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 gpio0_output[0]
port 39 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 gpio0_output[10]
port 40 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 gpio0_output[11]
port 41 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 gpio0_output[12]
port 42 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 gpio0_output[13]
port 43 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 gpio0_output[14]
port 44 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 gpio0_output[15]
port 45 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 gpio0_output[16]
port 46 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 gpio0_output[17]
port 47 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 gpio0_output[18]
port 48 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 gpio0_output[1]
port 49 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 gpio0_output[2]
port 50 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 gpio0_output[3]
port 51 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 gpio0_output[4]
port 52 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 gpio0_output[5]
port 53 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 gpio0_output[6]
port 54 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gpio0_output[7]
port 55 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 gpio0_output[8]
port 56 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 gpio0_output[9]
port 57 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 gpio1_input[0]
port 58 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 gpio1_input[10]
port 59 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 gpio1_input[11]
port 60 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 gpio1_input[12]
port 61 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 gpio1_input[13]
port 62 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 gpio1_input[14]
port 63 nsew signal tristate
rlabel metal2 s 21178 0 21234 800 6 gpio1_input[15]
port 64 nsew signal tristate
rlabel metal2 s 22006 0 22062 800 6 gpio1_input[16]
port 65 nsew signal tristate
rlabel metal2 s 22834 0 22890 800 6 gpio1_input[17]
port 66 nsew signal tristate
rlabel metal2 s 23662 0 23718 800 6 gpio1_input[18]
port 67 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 gpio1_input[1]
port 68 nsew signal tristate
rlabel metal2 s 10506 0 10562 800 6 gpio1_input[2]
port 69 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 gpio1_input[3]
port 70 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 gpio1_input[4]
port 71 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 gpio1_input[5]
port 72 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 gpio1_input[6]
port 73 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 gpio1_input[7]
port 74 nsew signal tristate
rlabel metal2 s 15382 0 15438 800 6 gpio1_input[8]
port 75 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 gpio1_input[9]
port 76 nsew signal tristate
rlabel metal2 s 9126 0 9182 800 6 gpio1_oe[0]
port 77 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 gpio1_oe[10]
port 78 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 gpio1_oe[11]
port 79 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 gpio1_oe[12]
port 80 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 gpio1_oe[13]
port 81 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 gpio1_oe[14]
port 82 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 gpio1_oe[15]
port 83 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 gpio1_oe[16]
port 84 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 gpio1_oe[17]
port 85 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 gpio1_oe[18]
port 86 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 gpio1_oe[1]
port 87 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 gpio1_oe[2]
port 88 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 gpio1_oe[3]
port 89 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 gpio1_oe[4]
port 90 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 gpio1_oe[5]
port 91 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 gpio1_oe[6]
port 92 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 gpio1_oe[7]
port 93 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 gpio1_oe[8]
port 94 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 gpio1_oe[9]
port 95 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 gpio1_output[0]
port 96 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 gpio1_output[10]
port 97 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 gpio1_output[11]
port 98 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 gpio1_output[12]
port 99 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 gpio1_output[13]
port 100 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 gpio1_output[14]
port 101 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 gpio1_output[15]
port 102 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 gpio1_output[16]
port 103 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 gpio1_output[17]
port 104 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 gpio1_output[18]
port 105 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 gpio1_output[1]
port 106 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 gpio1_output[2]
port 107 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 gpio1_output[3]
port 108 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 gpio1_output[4]
port 109 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 gpio1_output[5]
port 110 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 gpio1_output[6]
port 111 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 gpio1_output[7]
port 112 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 gpio1_output[8]
port 113 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 gpio1_output[9]
port 114 nsew signal input
rlabel metal2 s 110 39200 166 40000 6 io_in[0]
port 115 nsew signal input
rlabel metal2 s 10598 39200 10654 40000 6 io_in[10]
port 116 nsew signal input
rlabel metal2 s 11610 39200 11666 40000 6 io_in[11]
port 117 nsew signal input
rlabel metal2 s 12714 39200 12770 40000 6 io_in[12]
port 118 nsew signal input
rlabel metal2 s 13726 39200 13782 40000 6 io_in[13]
port 119 nsew signal input
rlabel metal2 s 14830 39200 14886 40000 6 io_in[14]
port 120 nsew signal input
rlabel metal2 s 15842 39200 15898 40000 6 io_in[15]
port 121 nsew signal input
rlabel metal2 s 16946 39200 17002 40000 6 io_in[16]
port 122 nsew signal input
rlabel metal2 s 17958 39200 18014 40000 6 io_in[17]
port 123 nsew signal input
rlabel metal2 s 19062 39200 19118 40000 6 io_in[18]
port 124 nsew signal input
rlabel metal2 s 20074 39200 20130 40000 6 io_in[19]
port 125 nsew signal input
rlabel metal2 s 1122 39200 1178 40000 6 io_in[1]
port 126 nsew signal input
rlabel metal2 s 21086 39200 21142 40000 6 io_in[20]
port 127 nsew signal input
rlabel metal2 s 22190 39200 22246 40000 6 io_in[21]
port 128 nsew signal input
rlabel metal2 s 23202 39200 23258 40000 6 io_in[22]
port 129 nsew signal input
rlabel metal2 s 24306 39200 24362 40000 6 io_in[23]
port 130 nsew signal input
rlabel metal2 s 25318 39200 25374 40000 6 io_in[24]
port 131 nsew signal input
rlabel metal2 s 26422 39200 26478 40000 6 io_in[25]
port 132 nsew signal input
rlabel metal2 s 27434 39200 27490 40000 6 io_in[26]
port 133 nsew signal input
rlabel metal2 s 28538 39200 28594 40000 6 io_in[27]
port 134 nsew signal input
rlabel metal2 s 29550 39200 29606 40000 6 io_in[28]
port 135 nsew signal input
rlabel metal2 s 30562 39200 30618 40000 6 io_in[29]
port 136 nsew signal input
rlabel metal2 s 2134 39200 2190 40000 6 io_in[2]
port 137 nsew signal input
rlabel metal2 s 31666 39200 31722 40000 6 io_in[30]
port 138 nsew signal input
rlabel metal2 s 32678 39200 32734 40000 6 io_in[31]
port 139 nsew signal input
rlabel metal2 s 33782 39200 33838 40000 6 io_in[32]
port 140 nsew signal input
rlabel metal2 s 34794 39200 34850 40000 6 io_in[33]
port 141 nsew signal input
rlabel metal2 s 35898 39200 35954 40000 6 io_in[34]
port 142 nsew signal input
rlabel metal2 s 36910 39200 36966 40000 6 io_in[35]
port 143 nsew signal input
rlabel metal2 s 38014 39200 38070 40000 6 io_in[36]
port 144 nsew signal input
rlabel metal2 s 39026 39200 39082 40000 6 io_in[37]
port 145 nsew signal input
rlabel metal2 s 3238 39200 3294 40000 6 io_in[3]
port 146 nsew signal input
rlabel metal2 s 4250 39200 4306 40000 6 io_in[4]
port 147 nsew signal input
rlabel metal2 s 5354 39200 5410 40000 6 io_in[5]
port 148 nsew signal input
rlabel metal2 s 6366 39200 6422 40000 6 io_in[6]
port 149 nsew signal input
rlabel metal2 s 7470 39200 7526 40000 6 io_in[7]
port 150 nsew signal input
rlabel metal2 s 8482 39200 8538 40000 6 io_in[8]
port 151 nsew signal input
rlabel metal2 s 9586 39200 9642 40000 6 io_in[9]
port 152 nsew signal input
rlabel metal2 s 386 39200 442 40000 6 io_oeb[0]
port 153 nsew signal tristate
rlabel metal2 s 10966 39200 11022 40000 6 io_oeb[10]
port 154 nsew signal tristate
rlabel metal2 s 11978 39200 12034 40000 6 io_oeb[11]
port 155 nsew signal tristate
rlabel metal2 s 13082 39200 13138 40000 6 io_oeb[12]
port 156 nsew signal tristate
rlabel metal2 s 14094 39200 14150 40000 6 io_oeb[13]
port 157 nsew signal tristate
rlabel metal2 s 15198 39200 15254 40000 6 io_oeb[14]
port 158 nsew signal tristate
rlabel metal2 s 16210 39200 16266 40000 6 io_oeb[15]
port 159 nsew signal tristate
rlabel metal2 s 17222 39200 17278 40000 6 io_oeb[16]
port 160 nsew signal tristate
rlabel metal2 s 18326 39200 18382 40000 6 io_oeb[17]
port 161 nsew signal tristate
rlabel metal2 s 19338 39200 19394 40000 6 io_oeb[18]
port 162 nsew signal tristate
rlabel metal2 s 20442 39200 20498 40000 6 io_oeb[19]
port 163 nsew signal tristate
rlabel metal2 s 1490 39200 1546 40000 6 io_oeb[1]
port 164 nsew signal tristate
rlabel metal2 s 21454 39200 21510 40000 6 io_oeb[20]
port 165 nsew signal tristate
rlabel metal2 s 22558 39200 22614 40000 6 io_oeb[21]
port 166 nsew signal tristate
rlabel metal2 s 23570 39200 23626 40000 6 io_oeb[22]
port 167 nsew signal tristate
rlabel metal2 s 24674 39200 24730 40000 6 io_oeb[23]
port 168 nsew signal tristate
rlabel metal2 s 25686 39200 25742 40000 6 io_oeb[24]
port 169 nsew signal tristate
rlabel metal2 s 26790 39200 26846 40000 6 io_oeb[25]
port 170 nsew signal tristate
rlabel metal2 s 27802 39200 27858 40000 6 io_oeb[26]
port 171 nsew signal tristate
rlabel metal2 s 28814 39200 28870 40000 6 io_oeb[27]
port 172 nsew signal tristate
rlabel metal2 s 29918 39200 29974 40000 6 io_oeb[28]
port 173 nsew signal tristate
rlabel metal2 s 30930 39200 30986 40000 6 io_oeb[29]
port 174 nsew signal tristate
rlabel metal2 s 2502 39200 2558 40000 6 io_oeb[2]
port 175 nsew signal tristate
rlabel metal2 s 32034 39200 32090 40000 6 io_oeb[30]
port 176 nsew signal tristate
rlabel metal2 s 33046 39200 33102 40000 6 io_oeb[31]
port 177 nsew signal tristate
rlabel metal2 s 34150 39200 34206 40000 6 io_oeb[32]
port 178 nsew signal tristate
rlabel metal2 s 35162 39200 35218 40000 6 io_oeb[33]
port 179 nsew signal tristate
rlabel metal2 s 36266 39200 36322 40000 6 io_oeb[34]
port 180 nsew signal tristate
rlabel metal2 s 37278 39200 37334 40000 6 io_oeb[35]
port 181 nsew signal tristate
rlabel metal2 s 38290 39200 38346 40000 6 io_oeb[36]
port 182 nsew signal tristate
rlabel metal2 s 39394 39200 39450 40000 6 io_oeb[37]
port 183 nsew signal tristate
rlabel metal2 s 3606 39200 3662 40000 6 io_oeb[3]
port 184 nsew signal tristate
rlabel metal2 s 4618 39200 4674 40000 6 io_oeb[4]
port 185 nsew signal tristate
rlabel metal2 s 5722 39200 5778 40000 6 io_oeb[5]
port 186 nsew signal tristate
rlabel metal2 s 6734 39200 6790 40000 6 io_oeb[6]
port 187 nsew signal tristate
rlabel metal2 s 7746 39200 7802 40000 6 io_oeb[7]
port 188 nsew signal tristate
rlabel metal2 s 8850 39200 8906 40000 6 io_oeb[8]
port 189 nsew signal tristate
rlabel metal2 s 9862 39200 9918 40000 6 io_oeb[9]
port 190 nsew signal tristate
rlabel metal2 s 754 39200 810 40000 6 io_out[0]
port 191 nsew signal tristate
rlabel metal2 s 11334 39200 11390 40000 6 io_out[10]
port 192 nsew signal tristate
rlabel metal2 s 12346 39200 12402 40000 6 io_out[11]
port 193 nsew signal tristate
rlabel metal2 s 13450 39200 13506 40000 6 io_out[12]
port 194 nsew signal tristate
rlabel metal2 s 14462 39200 14518 40000 6 io_out[13]
port 195 nsew signal tristate
rlabel metal2 s 15474 39200 15530 40000 6 io_out[14]
port 196 nsew signal tristate
rlabel metal2 s 16578 39200 16634 40000 6 io_out[15]
port 197 nsew signal tristate
rlabel metal2 s 17590 39200 17646 40000 6 io_out[16]
port 198 nsew signal tristate
rlabel metal2 s 18694 39200 18750 40000 6 io_out[17]
port 199 nsew signal tristate
rlabel metal2 s 19706 39200 19762 40000 6 io_out[18]
port 200 nsew signal tristate
rlabel metal2 s 20810 39200 20866 40000 6 io_out[19]
port 201 nsew signal tristate
rlabel metal2 s 1858 39200 1914 40000 6 io_out[1]
port 202 nsew signal tristate
rlabel metal2 s 21822 39200 21878 40000 6 io_out[20]
port 203 nsew signal tristate
rlabel metal2 s 22926 39200 22982 40000 6 io_out[21]
port 204 nsew signal tristate
rlabel metal2 s 23938 39200 23994 40000 6 io_out[22]
port 205 nsew signal tristate
rlabel metal2 s 24950 39200 25006 40000 6 io_out[23]
port 206 nsew signal tristate
rlabel metal2 s 26054 39200 26110 40000 6 io_out[24]
port 207 nsew signal tristate
rlabel metal2 s 27066 39200 27122 40000 6 io_out[25]
port 208 nsew signal tristate
rlabel metal2 s 28170 39200 28226 40000 6 io_out[26]
port 209 nsew signal tristate
rlabel metal2 s 29182 39200 29238 40000 6 io_out[27]
port 210 nsew signal tristate
rlabel metal2 s 30286 39200 30342 40000 6 io_out[28]
port 211 nsew signal tristate
rlabel metal2 s 31298 39200 31354 40000 6 io_out[29]
port 212 nsew signal tristate
rlabel metal2 s 2870 39200 2926 40000 6 io_out[2]
port 213 nsew signal tristate
rlabel metal2 s 32402 39200 32458 40000 6 io_out[30]
port 214 nsew signal tristate
rlabel metal2 s 33414 39200 33470 40000 6 io_out[31]
port 215 nsew signal tristate
rlabel metal2 s 34426 39200 34482 40000 6 io_out[32]
port 216 nsew signal tristate
rlabel metal2 s 35530 39200 35586 40000 6 io_out[33]
port 217 nsew signal tristate
rlabel metal2 s 36542 39200 36598 40000 6 io_out[34]
port 218 nsew signal tristate
rlabel metal2 s 37646 39200 37702 40000 6 io_out[35]
port 219 nsew signal tristate
rlabel metal2 s 38658 39200 38714 40000 6 io_out[36]
port 220 nsew signal tristate
rlabel metal2 s 39762 39200 39818 40000 6 io_out[37]
port 221 nsew signal tristate
rlabel metal2 s 3882 39200 3938 40000 6 io_out[3]
port 222 nsew signal tristate
rlabel metal2 s 4986 39200 5042 40000 6 io_out[4]
port 223 nsew signal tristate
rlabel metal2 s 5998 39200 6054 40000 6 io_out[5]
port 224 nsew signal tristate
rlabel metal2 s 7102 39200 7158 40000 6 io_out[6]
port 225 nsew signal tristate
rlabel metal2 s 8114 39200 8170 40000 6 io_out[7]
port 226 nsew signal tristate
rlabel metal2 s 9218 39200 9274 40000 6 io_out[8]
port 227 nsew signal tristate
rlabel metal2 s 10230 39200 10286 40000 6 io_out[9]
port 228 nsew signal tristate
rlabel metal3 s 39200 37408 40000 37528 6 la_blink[0]
port 229 nsew signal tristate
rlabel metal3 s 39200 39040 40000 39160 6 la_blink[1]
port 230 nsew signal tristate
rlabel metal2 s 110 0 166 800 6 pwm_en[0]
port 231 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 pwm_en[10]
port 232 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 pwm_en[11]
port 233 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 pwm_en[12]
port 234 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 pwm_en[13]
port 235 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 pwm_en[14]
port 236 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 pwm_en[15]
port 237 nsew signal input
rlabel metal2 s 570 0 626 800 6 pwm_en[1]
port 238 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 pwm_en[2]
port 239 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 pwm_en[3]
port 240 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 pwm_en[4]
port 241 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 pwm_en[5]
port 242 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 pwm_en[6]
port 243 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 pwm_en[7]
port 244 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 pwm_en[8]
port 245 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 pwm_en[9]
port 246 nsew signal input
rlabel metal2 s 294 0 350 800 6 pwm_out[0]
port 247 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 pwm_out[10]
port 248 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 pwm_out[11]
port 249 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 pwm_out[12]
port 250 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 pwm_out[13]
port 251 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 pwm_out[14]
port 252 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 pwm_out[15]
port 253 nsew signal input
rlabel metal2 s 846 0 902 800 6 pwm_out[1]
port 254 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 pwm_out[2]
port 255 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 pwm_out[3]
port 256 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 pwm_out[4]
port 257 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 pwm_out[5]
port 258 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 pwm_out[6]
port 259 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 pwm_out[7]
port 260 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 pwm_out[8]
port 261 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 pwm_out[9]
port 262 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 rst
port 263 nsew signal input
rlabel metal3 s 39200 20816 40000 20936 6 spi_clk[0]
port 264 nsew signal input
rlabel metal3 s 39200 29112 40000 29232 6 spi_clk[1]
port 265 nsew signal input
rlabel metal3 s 39200 22448 40000 22568 6 spi_cs[0]
port 266 nsew signal input
rlabel metal3 s 39200 30744 40000 30864 6 spi_cs[1]
port 267 nsew signal input
rlabel metal3 s 39200 24080 40000 24200 6 spi_en[0]
port 268 nsew signal input
rlabel metal3 s 39200 32376 40000 32496 6 spi_en[1]
port 269 nsew signal input
rlabel metal3 s 39200 25712 40000 25832 6 spi_miso[0]
port 270 nsew signal tristate
rlabel metal3 s 39200 34144 40000 34264 6 spi_miso[1]
port 271 nsew signal tristate
rlabel metal3 s 39200 27480 40000 27600 6 spi_mosi[0]
port 272 nsew signal input
rlabel metal3 s 39200 35776 40000 35896 6 spi_mosi[1]
port 273 nsew signal input
rlabel metal3 s 39200 824 40000 944 6 uart_en[0]
port 274 nsew signal input
rlabel metal3 s 39200 5720 40000 5840 6 uart_en[1]
port 275 nsew signal input
rlabel metal3 s 39200 10752 40000 10872 6 uart_en[2]
port 276 nsew signal input
rlabel metal3 s 39200 15784 40000 15904 6 uart_en[3]
port 277 nsew signal input
rlabel metal3 s 39200 2456 40000 2576 6 uart_rx[0]
port 278 nsew signal tristate
rlabel metal3 s 39200 7488 40000 7608 6 uart_rx[1]
port 279 nsew signal tristate
rlabel metal3 s 39200 12384 40000 12504 6 uart_rx[2]
port 280 nsew signal tristate
rlabel metal3 s 39200 17416 40000 17536 6 uart_rx[3]
port 281 nsew signal tristate
rlabel metal3 s 39200 4088 40000 4208 6 uart_tx[0]
port 282 nsew signal input
rlabel metal3 s 39200 9120 40000 9240 6 uart_tx[1]
port 283 nsew signal input
rlabel metal3 s 39200 14152 40000 14272 6 uart_tx[2]
port 284 nsew signal input
rlabel metal3 s 39200 19048 40000 19168 6 uart_tx[3]
port 285 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 286 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 286 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 287 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
